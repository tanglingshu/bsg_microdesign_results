

module top
(
  clk_i,
  data_i,
  sel_i,
  data_o
);

  input [63:0] data_i;
  input [1023:0] sel_i;
  output [63:0] data_o;
  input clk_i;

  bsg_fifo_shift_datapath
  wrapper
  (
    .data_i(data_i),
    .sel_i(sel_i),
    .data_o(data_o),
    .clk_i(clk_i)
  );


endmodule



module bsg_fifo_shift_datapath
(
  clk_i,
  data_i,
  sel_i,
  data_o
);

  input [63:0] data_i;
  input [1023:0] sel_i;
  output [63:0] data_o;
  input clk_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
  N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,
  N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,
  N1025,N1026,N1027,N1028,r_n_0__63_,r_n_0__62_,r_n_0__61_,r_n_0__60_,r_n_0__59_,
  r_n_0__58_,r_n_0__57_,r_n_0__56_,r_n_0__55_,r_n_0__54_,r_n_0__53_,r_n_0__52_,
  r_n_0__51_,r_n_0__50_,r_n_0__49_,r_n_0__48_,r_n_0__47_,r_n_0__46_,r_n_0__45_,
  r_n_0__44_,r_n_0__43_,r_n_0__42_,r_n_0__41_,r_n_0__40_,r_n_0__39_,r_n_0__38_,
  r_n_0__37_,r_n_0__36_,r_n_0__35_,r_n_0__34_,r_n_0__33_,r_n_0__32_,r_n_0__31_,r_n_0__30_,
  r_n_0__29_,r_n_0__28_,r_n_0__27_,r_n_0__26_,r_n_0__25_,r_n_0__24_,r_n_0__23_,
  r_n_0__22_,r_n_0__21_,r_n_0__20_,r_n_0__19_,r_n_0__18_,r_n_0__17_,r_n_0__16_,
  r_n_0__15_,r_n_0__14_,r_n_0__13_,r_n_0__12_,r_n_0__11_,r_n_0__10_,r_n_0__9_,r_n_0__8_,
  r_n_0__7_,r_n_0__6_,r_n_0__5_,r_n_0__4_,r_n_0__3_,r_n_0__2_,r_n_0__1_,r_n_0__0_,
  r_n_8__63_,r_n_8__62_,r_n_8__61_,r_n_8__60_,r_n_8__59_,r_n_8__58_,r_n_8__57_,
  r_n_8__56_,r_n_8__55_,r_n_8__54_,r_n_8__53_,r_n_8__52_,r_n_8__51_,r_n_8__50_,
  r_n_8__49_,r_n_8__48_,r_n_8__47_,r_n_8__46_,r_n_8__45_,r_n_8__44_,r_n_8__43_,r_n_8__42_,
  r_n_8__41_,r_n_8__40_,r_n_8__39_,r_n_8__38_,r_n_8__37_,r_n_8__36_,r_n_8__35_,
  r_n_8__34_,r_n_8__33_,r_n_8__32_,r_n_8__31_,r_n_8__30_,r_n_8__29_,r_n_8__28_,
  r_n_8__27_,r_n_8__26_,r_n_8__25_,r_n_8__24_,r_n_8__23_,r_n_8__22_,r_n_8__21_,
  r_n_8__20_,r_n_8__19_,r_n_8__18_,r_n_8__17_,r_n_8__16_,r_n_8__15_,r_n_8__14_,r_n_8__13_,
  r_n_8__12_,r_n_8__11_,r_n_8__10_,r_n_8__9_,r_n_8__8_,r_n_8__7_,r_n_8__6_,
  r_n_8__5_,r_n_8__4_,r_n_8__3_,r_n_8__2_,r_n_8__1_,r_n_8__0_,r_n_7__63_,r_n_7__62_,
  r_n_7__61_,r_n_7__60_,r_n_7__59_,r_n_7__58_,r_n_7__57_,r_n_7__56_,r_n_7__55_,
  r_n_7__54_,r_n_7__53_,r_n_7__52_,r_n_7__51_,r_n_7__50_,r_n_7__49_,r_n_7__48_,r_n_7__47_,
  r_n_7__46_,r_n_7__45_,r_n_7__44_,r_n_7__43_,r_n_7__42_,r_n_7__41_,r_n_7__40_,
  r_n_7__39_,r_n_7__38_,r_n_7__37_,r_n_7__36_,r_n_7__35_,r_n_7__34_,r_n_7__33_,
  r_n_7__32_,r_n_7__31_,r_n_7__30_,r_n_7__29_,r_n_7__28_,r_n_7__27_,r_n_7__26_,
  r_n_7__25_,r_n_7__24_,r_n_7__23_,r_n_7__22_,r_n_7__21_,r_n_7__20_,r_n_7__19_,r_n_7__18_,
  r_n_7__17_,r_n_7__16_,r_n_7__15_,r_n_7__14_,r_n_7__13_,r_n_7__12_,r_n_7__11_,
  r_n_7__10_,r_n_7__9_,r_n_7__8_,r_n_7__7_,r_n_7__6_,r_n_7__5_,r_n_7__4_,r_n_7__3_,
  r_n_7__2_,r_n_7__1_,r_n_7__0_,r_n_6__63_,r_n_6__62_,r_n_6__61_,r_n_6__60_,
  r_n_6__59_,r_n_6__58_,r_n_6__57_,r_n_6__56_,r_n_6__55_,r_n_6__54_,r_n_6__53_,r_n_6__52_,
  r_n_6__51_,r_n_6__50_,r_n_6__49_,r_n_6__48_,r_n_6__47_,r_n_6__46_,r_n_6__45_,
  r_n_6__44_,r_n_6__43_,r_n_6__42_,r_n_6__41_,r_n_6__40_,r_n_6__39_,r_n_6__38_,
  r_n_6__37_,r_n_6__36_,r_n_6__35_,r_n_6__34_,r_n_6__33_,r_n_6__32_,r_n_6__31_,r_n_6__30_,
  r_n_6__29_,r_n_6__28_,r_n_6__27_,r_n_6__26_,r_n_6__25_,r_n_6__24_,r_n_6__23_,
  r_n_6__22_,r_n_6__21_,r_n_6__20_,r_n_6__19_,r_n_6__18_,r_n_6__17_,r_n_6__16_,
  r_n_6__15_,r_n_6__14_,r_n_6__13_,r_n_6__12_,r_n_6__11_,r_n_6__10_,r_n_6__9_,r_n_6__8_,
  r_n_6__7_,r_n_6__6_,r_n_6__5_,r_n_6__4_,r_n_6__3_,r_n_6__2_,r_n_6__1_,r_n_6__0_,
  r_n_5__63_,r_n_5__62_,r_n_5__61_,r_n_5__60_,r_n_5__59_,r_n_5__58_,r_n_5__57_,
  r_n_5__56_,r_n_5__55_,r_n_5__54_,r_n_5__53_,r_n_5__52_,r_n_5__51_,r_n_5__50_,
  r_n_5__49_,r_n_5__48_,r_n_5__47_,r_n_5__46_,r_n_5__45_,r_n_5__44_,r_n_5__43_,
  r_n_5__42_,r_n_5__41_,r_n_5__40_,r_n_5__39_,r_n_5__38_,r_n_5__37_,r_n_5__36_,r_n_5__35_,
  r_n_5__34_,r_n_5__33_,r_n_5__32_,r_n_5__31_,r_n_5__30_,r_n_5__29_,r_n_5__28_,
  r_n_5__27_,r_n_5__26_,r_n_5__25_,r_n_5__24_,r_n_5__23_,r_n_5__22_,r_n_5__21_,
  r_n_5__20_,r_n_5__19_,r_n_5__18_,r_n_5__17_,r_n_5__16_,r_n_5__15_,r_n_5__14_,
  r_n_5__13_,r_n_5__12_,r_n_5__11_,r_n_5__10_,r_n_5__9_,r_n_5__8_,r_n_5__7_,r_n_5__6_,
  r_n_5__5_,r_n_5__4_,r_n_5__3_,r_n_5__2_,r_n_5__1_,r_n_5__0_,r_n_4__63_,r_n_4__62_,
  r_n_4__61_,r_n_4__60_,r_n_4__59_,r_n_4__58_,r_n_4__57_,r_n_4__56_,r_n_4__55_,
  r_n_4__54_,r_n_4__53_,r_n_4__52_,r_n_4__51_,r_n_4__50_,r_n_4__49_,r_n_4__48_,
  r_n_4__47_,r_n_4__46_,r_n_4__45_,r_n_4__44_,r_n_4__43_,r_n_4__42_,r_n_4__41_,r_n_4__40_,
  r_n_4__39_,r_n_4__38_,r_n_4__37_,r_n_4__36_,r_n_4__35_,r_n_4__34_,r_n_4__33_,
  r_n_4__32_,r_n_4__31_,r_n_4__30_,r_n_4__29_,r_n_4__28_,r_n_4__27_,r_n_4__26_,
  r_n_4__25_,r_n_4__24_,r_n_4__23_,r_n_4__22_,r_n_4__21_,r_n_4__20_,r_n_4__19_,r_n_4__18_,
  r_n_4__17_,r_n_4__16_,r_n_4__15_,r_n_4__14_,r_n_4__13_,r_n_4__12_,r_n_4__11_,
  r_n_4__10_,r_n_4__9_,r_n_4__8_,r_n_4__7_,r_n_4__6_,r_n_4__5_,r_n_4__4_,r_n_4__3_,
  r_n_4__2_,r_n_4__1_,r_n_4__0_,r_n_3__63_,r_n_3__62_,r_n_3__61_,r_n_3__60_,
  r_n_3__59_,r_n_3__58_,r_n_3__57_,r_n_3__56_,r_n_3__55_,r_n_3__54_,r_n_3__53_,r_n_3__52_,
  r_n_3__51_,r_n_3__50_,r_n_3__49_,r_n_3__48_,r_n_3__47_,r_n_3__46_,r_n_3__45_,
  r_n_3__44_,r_n_3__43_,r_n_3__42_,r_n_3__41_,r_n_3__40_,r_n_3__39_,r_n_3__38_,
  r_n_3__37_,r_n_3__36_,r_n_3__35_,r_n_3__34_,r_n_3__33_,r_n_3__32_,r_n_3__31_,
  r_n_3__30_,r_n_3__29_,r_n_3__28_,r_n_3__27_,r_n_3__26_,r_n_3__25_,r_n_3__24_,r_n_3__23_,
  r_n_3__22_,r_n_3__21_,r_n_3__20_,r_n_3__19_,r_n_3__18_,r_n_3__17_,r_n_3__16_,
  r_n_3__15_,r_n_3__14_,r_n_3__13_,r_n_3__12_,r_n_3__11_,r_n_3__10_,r_n_3__9_,
  r_n_3__8_,r_n_3__7_,r_n_3__6_,r_n_3__5_,r_n_3__4_,r_n_3__3_,r_n_3__2_,r_n_3__1_,
  r_n_3__0_,r_n_2__63_,r_n_2__62_,r_n_2__61_,r_n_2__60_,r_n_2__59_,r_n_2__58_,r_n_2__57_,
  r_n_2__56_,r_n_2__55_,r_n_2__54_,r_n_2__53_,r_n_2__52_,r_n_2__51_,r_n_2__50_,
  r_n_2__49_,r_n_2__48_,r_n_2__47_,r_n_2__46_,r_n_2__45_,r_n_2__44_,r_n_2__43_,
  r_n_2__42_,r_n_2__41_,r_n_2__40_,r_n_2__39_,r_n_2__38_,r_n_2__37_,r_n_2__36_,
  r_n_2__35_,r_n_2__34_,r_n_2__33_,r_n_2__32_,r_n_2__31_,r_n_2__30_,r_n_2__29_,r_n_2__28_,
  r_n_2__27_,r_n_2__26_,r_n_2__25_,r_n_2__24_,r_n_2__23_,r_n_2__22_,r_n_2__21_,
  r_n_2__20_,r_n_2__19_,r_n_2__18_,r_n_2__17_,r_n_2__16_,r_n_2__15_,r_n_2__14_,
  r_n_2__13_,r_n_2__12_,r_n_2__11_,r_n_2__10_,r_n_2__9_,r_n_2__8_,r_n_2__7_,r_n_2__6_,
  r_n_2__5_,r_n_2__4_,r_n_2__3_,r_n_2__2_,r_n_2__1_,r_n_2__0_,r_n_1__63_,r_n_1__62_,
  r_n_1__61_,r_n_1__60_,r_n_1__59_,r_n_1__58_,r_n_1__57_,r_n_1__56_,r_n_1__55_,
  r_n_1__54_,r_n_1__53_,r_n_1__52_,r_n_1__51_,r_n_1__50_,r_n_1__49_,r_n_1__48_,
  r_n_1__47_,r_n_1__46_,r_n_1__45_,r_n_1__44_,r_n_1__43_,r_n_1__42_,r_n_1__41_,r_n_1__40_,
  r_n_1__39_,r_n_1__38_,r_n_1__37_,r_n_1__36_,r_n_1__35_,r_n_1__34_,r_n_1__33_,
  r_n_1__32_,r_n_1__31_,r_n_1__30_,r_n_1__29_,r_n_1__28_,r_n_1__27_,r_n_1__26_,
  r_n_1__25_,r_n_1__24_,r_n_1__23_,r_n_1__22_,r_n_1__21_,r_n_1__20_,r_n_1__19_,
  r_n_1__18_,r_n_1__17_,r_n_1__16_,r_n_1__15_,r_n_1__14_,r_n_1__13_,r_n_1__12_,r_n_1__11_,
  r_n_1__10_,r_n_1__9_,r_n_1__8_,r_n_1__7_,r_n_1__6_,r_n_1__5_,r_n_1__4_,r_n_1__3_,
  r_n_1__2_,r_n_1__1_,r_n_1__0_,r_n_16__63_,r_n_16__62_,r_n_16__61_,r_n_16__60_,
  r_n_16__59_,r_n_16__58_,r_n_16__57_,r_n_16__56_,r_n_16__55_,r_n_16__54_,
  r_n_16__53_,r_n_16__52_,r_n_16__51_,r_n_16__50_,r_n_16__49_,r_n_16__48_,r_n_16__47_,
  r_n_16__46_,r_n_16__45_,r_n_16__44_,r_n_16__43_,r_n_16__42_,r_n_16__41_,r_n_16__40_,
  r_n_16__39_,r_n_16__38_,r_n_16__37_,r_n_16__36_,r_n_16__35_,r_n_16__34_,
  r_n_16__33_,r_n_16__32_,r_n_16__31_,r_n_16__30_,r_n_16__29_,r_n_16__28_,r_n_16__27_,
  r_n_16__26_,r_n_16__25_,r_n_16__24_,r_n_16__23_,r_n_16__22_,r_n_16__21_,r_n_16__20_,
  r_n_16__19_,r_n_16__18_,r_n_16__17_,r_n_16__16_,r_n_16__15_,r_n_16__14_,
  r_n_16__13_,r_n_16__12_,r_n_16__11_,r_n_16__10_,r_n_16__9_,r_n_16__8_,r_n_16__7_,
  r_n_16__6_,r_n_16__5_,r_n_16__4_,r_n_16__3_,r_n_16__2_,r_n_16__1_,r_n_16__0_,r_n_15__63_,
  r_n_15__62_,r_n_15__61_,r_n_15__60_,r_n_15__59_,r_n_15__58_,r_n_15__57_,
  r_n_15__56_,r_n_15__55_,r_n_15__54_,r_n_15__53_,r_n_15__52_,r_n_15__51_,r_n_15__50_,
  r_n_15__49_,r_n_15__48_,r_n_15__47_,r_n_15__46_,r_n_15__45_,r_n_15__44_,r_n_15__43_,
  r_n_15__42_,r_n_15__41_,r_n_15__40_,r_n_15__39_,r_n_15__38_,r_n_15__37_,
  r_n_15__36_,r_n_15__35_,r_n_15__34_,r_n_15__33_,r_n_15__32_,r_n_15__31_,r_n_15__30_,
  r_n_15__29_,r_n_15__28_,r_n_15__27_,r_n_15__26_,r_n_15__25_,r_n_15__24_,r_n_15__23_,
  r_n_15__22_,r_n_15__21_,r_n_15__20_,r_n_15__19_,r_n_15__18_,r_n_15__17_,
  r_n_15__16_,r_n_15__15_,r_n_15__14_,r_n_15__13_,r_n_15__12_,r_n_15__11_,r_n_15__10_,
  r_n_15__9_,r_n_15__8_,r_n_15__7_,r_n_15__6_,r_n_15__5_,r_n_15__4_,r_n_15__3_,
  r_n_15__2_,r_n_15__1_,r_n_15__0_,r_n_14__63_,r_n_14__62_,r_n_14__61_,r_n_14__60_,
  r_n_14__59_,r_n_14__58_,r_n_14__57_,r_n_14__56_,r_n_14__55_,r_n_14__54_,r_n_14__53_,
  r_n_14__52_,r_n_14__51_,r_n_14__50_,r_n_14__49_,r_n_14__48_,r_n_14__47_,
  r_n_14__46_,r_n_14__45_,r_n_14__44_,r_n_14__43_,r_n_14__42_,r_n_14__41_,r_n_14__40_,
  r_n_14__39_,r_n_14__38_,r_n_14__37_,r_n_14__36_,r_n_14__35_,r_n_14__34_,r_n_14__33_,
  r_n_14__32_,r_n_14__31_,r_n_14__30_,r_n_14__29_,r_n_14__28_,r_n_14__27_,
  r_n_14__26_,r_n_14__25_,r_n_14__24_,r_n_14__23_,r_n_14__22_,r_n_14__21_,r_n_14__20_,
  r_n_14__19_,r_n_14__18_,r_n_14__17_,r_n_14__16_,r_n_14__15_,r_n_14__14_,r_n_14__13_,
  r_n_14__12_,r_n_14__11_,r_n_14__10_,r_n_14__9_,r_n_14__8_,r_n_14__7_,r_n_14__6_,
  r_n_14__5_,r_n_14__4_,r_n_14__3_,r_n_14__2_,r_n_14__1_,r_n_14__0_,r_n_13__63_,
  r_n_13__62_,r_n_13__61_,r_n_13__60_,r_n_13__59_,r_n_13__58_,r_n_13__57_,r_n_13__56_,
  r_n_13__55_,r_n_13__54_,r_n_13__53_,r_n_13__52_,r_n_13__51_,r_n_13__50_,
  r_n_13__49_,r_n_13__48_,r_n_13__47_,r_n_13__46_,r_n_13__45_,r_n_13__44_,r_n_13__43_,
  r_n_13__42_,r_n_13__41_,r_n_13__40_,r_n_13__39_,r_n_13__38_,r_n_13__37_,r_n_13__36_,
  r_n_13__35_,r_n_13__34_,r_n_13__33_,r_n_13__32_,r_n_13__31_,r_n_13__30_,
  r_n_13__29_,r_n_13__28_,r_n_13__27_,r_n_13__26_,r_n_13__25_,r_n_13__24_,r_n_13__23_,
  r_n_13__22_,r_n_13__21_,r_n_13__20_,r_n_13__19_,r_n_13__18_,r_n_13__17_,r_n_13__16_,
  r_n_13__15_,r_n_13__14_,r_n_13__13_,r_n_13__12_,r_n_13__11_,r_n_13__10_,
  r_n_13__9_,r_n_13__8_,r_n_13__7_,r_n_13__6_,r_n_13__5_,r_n_13__4_,r_n_13__3_,r_n_13__2_,
  r_n_13__1_,r_n_13__0_,r_n_12__63_,r_n_12__62_,r_n_12__61_,r_n_12__60_,
  r_n_12__59_,r_n_12__58_,r_n_12__57_,r_n_12__56_,r_n_12__55_,r_n_12__54_,r_n_12__53_,
  r_n_12__52_,r_n_12__51_,r_n_12__50_,r_n_12__49_,r_n_12__48_,r_n_12__47_,r_n_12__46_,
  r_n_12__45_,r_n_12__44_,r_n_12__43_,r_n_12__42_,r_n_12__41_,r_n_12__40_,
  r_n_12__39_,r_n_12__38_,r_n_12__37_,r_n_12__36_,r_n_12__35_,r_n_12__34_,r_n_12__33_,
  r_n_12__32_,r_n_12__31_,r_n_12__30_,r_n_12__29_,r_n_12__28_,r_n_12__27_,r_n_12__26_,
  r_n_12__25_,r_n_12__24_,r_n_12__23_,r_n_12__22_,r_n_12__21_,r_n_12__20_,
  r_n_12__19_,r_n_12__18_,r_n_12__17_,r_n_12__16_,r_n_12__15_,r_n_12__14_,r_n_12__13_,
  r_n_12__12_,r_n_12__11_,r_n_12__10_,r_n_12__9_,r_n_12__8_,r_n_12__7_,r_n_12__6_,
  r_n_12__5_,r_n_12__4_,r_n_12__3_,r_n_12__2_,r_n_12__1_,r_n_12__0_,r_n_11__63_,
  r_n_11__62_,r_n_11__61_,r_n_11__60_,r_n_11__59_,r_n_11__58_,r_n_11__57_,r_n_11__56_,
  r_n_11__55_,r_n_11__54_,r_n_11__53_,r_n_11__52_,r_n_11__51_,r_n_11__50_,r_n_11__49_,
  r_n_11__48_,r_n_11__47_,r_n_11__46_,r_n_11__45_,r_n_11__44_,r_n_11__43_,
  r_n_11__42_,r_n_11__41_,r_n_11__40_,r_n_11__39_,r_n_11__38_,r_n_11__37_,r_n_11__36_,
  r_n_11__35_,r_n_11__34_,r_n_11__33_,r_n_11__32_,r_n_11__31_,r_n_11__30_,r_n_11__29_,
  r_n_11__28_,r_n_11__27_,r_n_11__26_,r_n_11__25_,r_n_11__24_,r_n_11__23_,
  r_n_11__22_,r_n_11__21_,r_n_11__20_,r_n_11__19_,r_n_11__18_,r_n_11__17_,r_n_11__16_,
  r_n_11__15_,r_n_11__14_,r_n_11__13_,r_n_11__12_,r_n_11__11_,r_n_11__10_,r_n_11__9_,
  r_n_11__8_,r_n_11__7_,r_n_11__6_,r_n_11__5_,r_n_11__4_,r_n_11__3_,r_n_11__2_,
  r_n_11__1_,r_n_11__0_,r_n_10__63_,r_n_10__62_,r_n_10__61_,r_n_10__60_,r_n_10__59_,
  r_n_10__58_,r_n_10__57_,r_n_10__56_,r_n_10__55_,r_n_10__54_,r_n_10__53_,
  r_n_10__52_,r_n_10__51_,r_n_10__50_,r_n_10__49_,r_n_10__48_,r_n_10__47_,r_n_10__46_,
  r_n_10__45_,r_n_10__44_,r_n_10__43_,r_n_10__42_,r_n_10__41_,r_n_10__40_,r_n_10__39_,
  r_n_10__38_,r_n_10__37_,r_n_10__36_,r_n_10__35_,r_n_10__34_,r_n_10__33_,
  r_n_10__32_,r_n_10__31_,r_n_10__30_,r_n_10__29_,r_n_10__28_,r_n_10__27_,r_n_10__26_,
  r_n_10__25_,r_n_10__24_,r_n_10__23_,r_n_10__22_,r_n_10__21_,r_n_10__20_,r_n_10__19_,
  r_n_10__18_,r_n_10__17_,r_n_10__16_,r_n_10__15_,r_n_10__14_,r_n_10__13_,
  r_n_10__12_,r_n_10__11_,r_n_10__10_,r_n_10__9_,r_n_10__8_,r_n_10__7_,r_n_10__6_,
  r_n_10__5_,r_n_10__4_,r_n_10__3_,r_n_10__2_,r_n_10__1_,r_n_10__0_,r_n_9__63_,r_n_9__62_,
  r_n_9__61_,r_n_9__60_,r_n_9__59_,r_n_9__58_,r_n_9__57_,r_n_9__56_,r_n_9__55_,
  r_n_9__54_,r_n_9__53_,r_n_9__52_,r_n_9__51_,r_n_9__50_,r_n_9__49_,r_n_9__48_,
  r_n_9__47_,r_n_9__46_,r_n_9__45_,r_n_9__44_,r_n_9__43_,r_n_9__42_,r_n_9__41_,r_n_9__40_,
  r_n_9__39_,r_n_9__38_,r_n_9__37_,r_n_9__36_,r_n_9__35_,r_n_9__34_,r_n_9__33_,
  r_n_9__32_,r_n_9__31_,r_n_9__30_,r_n_9__29_,r_n_9__28_,r_n_9__27_,r_n_9__26_,
  r_n_9__25_,r_n_9__24_,r_n_9__23_,r_n_9__22_,r_n_9__21_,r_n_9__20_,r_n_9__19_,
  r_n_9__18_,r_n_9__17_,r_n_9__16_,r_n_9__15_,r_n_9__14_,r_n_9__13_,r_n_9__12_,r_n_9__11_,
  r_n_9__10_,r_n_9__9_,r_n_9__8_,r_n_9__7_,r_n_9__6_,r_n_9__5_,r_n_9__4_,r_n_9__3_,
  r_n_9__2_,r_n_9__1_,r_n_9__0_,r_n_24__63_,r_n_24__62_,r_n_24__61_,r_n_24__60_,
  r_n_24__59_,r_n_24__58_,r_n_24__57_,r_n_24__56_,r_n_24__55_,r_n_24__54_,
  r_n_24__53_,r_n_24__52_,r_n_24__51_,r_n_24__50_,r_n_24__49_,r_n_24__48_,r_n_24__47_,
  r_n_24__46_,r_n_24__45_,r_n_24__44_,r_n_24__43_,r_n_24__42_,r_n_24__41_,r_n_24__40_,
  r_n_24__39_,r_n_24__38_,r_n_24__37_,r_n_24__36_,r_n_24__35_,r_n_24__34_,
  r_n_24__33_,r_n_24__32_,r_n_24__31_,r_n_24__30_,r_n_24__29_,r_n_24__28_,r_n_24__27_,
  r_n_24__26_,r_n_24__25_,r_n_24__24_,r_n_24__23_,r_n_24__22_,r_n_24__21_,r_n_24__20_,
  r_n_24__19_,r_n_24__18_,r_n_24__17_,r_n_24__16_,r_n_24__15_,r_n_24__14_,
  r_n_24__13_,r_n_24__12_,r_n_24__11_,r_n_24__10_,r_n_24__9_,r_n_24__8_,r_n_24__7_,
  r_n_24__6_,r_n_24__5_,r_n_24__4_,r_n_24__3_,r_n_24__2_,r_n_24__1_,r_n_24__0_,r_n_23__63_,
  r_n_23__62_,r_n_23__61_,r_n_23__60_,r_n_23__59_,r_n_23__58_,r_n_23__57_,
  r_n_23__56_,r_n_23__55_,r_n_23__54_,r_n_23__53_,r_n_23__52_,r_n_23__51_,r_n_23__50_,
  r_n_23__49_,r_n_23__48_,r_n_23__47_,r_n_23__46_,r_n_23__45_,r_n_23__44_,r_n_23__43_,
  r_n_23__42_,r_n_23__41_,r_n_23__40_,r_n_23__39_,r_n_23__38_,r_n_23__37_,
  r_n_23__36_,r_n_23__35_,r_n_23__34_,r_n_23__33_,r_n_23__32_,r_n_23__31_,r_n_23__30_,
  r_n_23__29_,r_n_23__28_,r_n_23__27_,r_n_23__26_,r_n_23__25_,r_n_23__24_,r_n_23__23_,
  r_n_23__22_,r_n_23__21_,r_n_23__20_,r_n_23__19_,r_n_23__18_,r_n_23__17_,
  r_n_23__16_,r_n_23__15_,r_n_23__14_,r_n_23__13_,r_n_23__12_,r_n_23__11_,r_n_23__10_,
  r_n_23__9_,r_n_23__8_,r_n_23__7_,r_n_23__6_,r_n_23__5_,r_n_23__4_,r_n_23__3_,
  r_n_23__2_,r_n_23__1_,r_n_23__0_,r_n_22__63_,r_n_22__62_,r_n_22__61_,r_n_22__60_,
  r_n_22__59_,r_n_22__58_,r_n_22__57_,r_n_22__56_,r_n_22__55_,r_n_22__54_,r_n_22__53_,
  r_n_22__52_,r_n_22__51_,r_n_22__50_,r_n_22__49_,r_n_22__48_,r_n_22__47_,
  r_n_22__46_,r_n_22__45_,r_n_22__44_,r_n_22__43_,r_n_22__42_,r_n_22__41_,r_n_22__40_,
  r_n_22__39_,r_n_22__38_,r_n_22__37_,r_n_22__36_,r_n_22__35_,r_n_22__34_,r_n_22__33_,
  r_n_22__32_,r_n_22__31_,r_n_22__30_,r_n_22__29_,r_n_22__28_,r_n_22__27_,
  r_n_22__26_,r_n_22__25_,r_n_22__24_,r_n_22__23_,r_n_22__22_,r_n_22__21_,r_n_22__20_,
  r_n_22__19_,r_n_22__18_,r_n_22__17_,r_n_22__16_,r_n_22__15_,r_n_22__14_,r_n_22__13_,
  r_n_22__12_,r_n_22__11_,r_n_22__10_,r_n_22__9_,r_n_22__8_,r_n_22__7_,r_n_22__6_,
  r_n_22__5_,r_n_22__4_,r_n_22__3_,r_n_22__2_,r_n_22__1_,r_n_22__0_,r_n_21__63_,
  r_n_21__62_,r_n_21__61_,r_n_21__60_,r_n_21__59_,r_n_21__58_,r_n_21__57_,r_n_21__56_,
  r_n_21__55_,r_n_21__54_,r_n_21__53_,r_n_21__52_,r_n_21__51_,r_n_21__50_,
  r_n_21__49_,r_n_21__48_,r_n_21__47_,r_n_21__46_,r_n_21__45_,r_n_21__44_,r_n_21__43_,
  r_n_21__42_,r_n_21__41_,r_n_21__40_,r_n_21__39_,r_n_21__38_,r_n_21__37_,r_n_21__36_,
  r_n_21__35_,r_n_21__34_,r_n_21__33_,r_n_21__32_,r_n_21__31_,r_n_21__30_,
  r_n_21__29_,r_n_21__28_,r_n_21__27_,r_n_21__26_,r_n_21__25_,r_n_21__24_,r_n_21__23_,
  r_n_21__22_,r_n_21__21_,r_n_21__20_,r_n_21__19_,r_n_21__18_,r_n_21__17_,r_n_21__16_,
  r_n_21__15_,r_n_21__14_,r_n_21__13_,r_n_21__12_,r_n_21__11_,r_n_21__10_,
  r_n_21__9_,r_n_21__8_,r_n_21__7_,r_n_21__6_,r_n_21__5_,r_n_21__4_,r_n_21__3_,r_n_21__2_,
  r_n_21__1_,r_n_21__0_,r_n_20__63_,r_n_20__62_,r_n_20__61_,r_n_20__60_,
  r_n_20__59_,r_n_20__58_,r_n_20__57_,r_n_20__56_,r_n_20__55_,r_n_20__54_,r_n_20__53_,
  r_n_20__52_,r_n_20__51_,r_n_20__50_,r_n_20__49_,r_n_20__48_,r_n_20__47_,r_n_20__46_,
  r_n_20__45_,r_n_20__44_,r_n_20__43_,r_n_20__42_,r_n_20__41_,r_n_20__40_,
  r_n_20__39_,r_n_20__38_,r_n_20__37_,r_n_20__36_,r_n_20__35_,r_n_20__34_,r_n_20__33_,
  r_n_20__32_,r_n_20__31_,r_n_20__30_,r_n_20__29_,r_n_20__28_,r_n_20__27_,r_n_20__26_,
  r_n_20__25_,r_n_20__24_,r_n_20__23_,r_n_20__22_,r_n_20__21_,r_n_20__20_,
  r_n_20__19_,r_n_20__18_,r_n_20__17_,r_n_20__16_,r_n_20__15_,r_n_20__14_,r_n_20__13_,
  r_n_20__12_,r_n_20__11_,r_n_20__10_,r_n_20__9_,r_n_20__8_,r_n_20__7_,r_n_20__6_,
  r_n_20__5_,r_n_20__4_,r_n_20__3_,r_n_20__2_,r_n_20__1_,r_n_20__0_,r_n_19__63_,
  r_n_19__62_,r_n_19__61_,r_n_19__60_,r_n_19__59_,r_n_19__58_,r_n_19__57_,r_n_19__56_,
  r_n_19__55_,r_n_19__54_,r_n_19__53_,r_n_19__52_,r_n_19__51_,r_n_19__50_,r_n_19__49_,
  r_n_19__48_,r_n_19__47_,r_n_19__46_,r_n_19__45_,r_n_19__44_,r_n_19__43_,
  r_n_19__42_,r_n_19__41_,r_n_19__40_,r_n_19__39_,r_n_19__38_,r_n_19__37_,r_n_19__36_,
  r_n_19__35_,r_n_19__34_,r_n_19__33_,r_n_19__32_,r_n_19__31_,r_n_19__30_,r_n_19__29_,
  r_n_19__28_,r_n_19__27_,r_n_19__26_,r_n_19__25_,r_n_19__24_,r_n_19__23_,
  r_n_19__22_,r_n_19__21_,r_n_19__20_,r_n_19__19_,r_n_19__18_,r_n_19__17_,r_n_19__16_,
  r_n_19__15_,r_n_19__14_,r_n_19__13_,r_n_19__12_,r_n_19__11_,r_n_19__10_,r_n_19__9_,
  r_n_19__8_,r_n_19__7_,r_n_19__6_,r_n_19__5_,r_n_19__4_,r_n_19__3_,r_n_19__2_,
  r_n_19__1_,r_n_19__0_,r_n_18__63_,r_n_18__62_,r_n_18__61_,r_n_18__60_,r_n_18__59_,
  r_n_18__58_,r_n_18__57_,r_n_18__56_,r_n_18__55_,r_n_18__54_,r_n_18__53_,
  r_n_18__52_,r_n_18__51_,r_n_18__50_,r_n_18__49_,r_n_18__48_,r_n_18__47_,r_n_18__46_,
  r_n_18__45_,r_n_18__44_,r_n_18__43_,r_n_18__42_,r_n_18__41_,r_n_18__40_,r_n_18__39_,
  r_n_18__38_,r_n_18__37_,r_n_18__36_,r_n_18__35_,r_n_18__34_,r_n_18__33_,
  r_n_18__32_,r_n_18__31_,r_n_18__30_,r_n_18__29_,r_n_18__28_,r_n_18__27_,r_n_18__26_,
  r_n_18__25_,r_n_18__24_,r_n_18__23_,r_n_18__22_,r_n_18__21_,r_n_18__20_,r_n_18__19_,
  r_n_18__18_,r_n_18__17_,r_n_18__16_,r_n_18__15_,r_n_18__14_,r_n_18__13_,
  r_n_18__12_,r_n_18__11_,r_n_18__10_,r_n_18__9_,r_n_18__8_,r_n_18__7_,r_n_18__6_,
  r_n_18__5_,r_n_18__4_,r_n_18__3_,r_n_18__2_,r_n_18__1_,r_n_18__0_,r_n_17__63_,r_n_17__62_,
  r_n_17__61_,r_n_17__60_,r_n_17__59_,r_n_17__58_,r_n_17__57_,r_n_17__56_,
  r_n_17__55_,r_n_17__54_,r_n_17__53_,r_n_17__52_,r_n_17__51_,r_n_17__50_,r_n_17__49_,
  r_n_17__48_,r_n_17__47_,r_n_17__46_,r_n_17__45_,r_n_17__44_,r_n_17__43_,r_n_17__42_,
  r_n_17__41_,r_n_17__40_,r_n_17__39_,r_n_17__38_,r_n_17__37_,r_n_17__36_,
  r_n_17__35_,r_n_17__34_,r_n_17__33_,r_n_17__32_,r_n_17__31_,r_n_17__30_,r_n_17__29_,
  r_n_17__28_,r_n_17__27_,r_n_17__26_,r_n_17__25_,r_n_17__24_,r_n_17__23_,r_n_17__22_,
  r_n_17__21_,r_n_17__20_,r_n_17__19_,r_n_17__18_,r_n_17__17_,r_n_17__16_,
  r_n_17__15_,r_n_17__14_,r_n_17__13_,r_n_17__12_,r_n_17__11_,r_n_17__10_,r_n_17__9_,
  r_n_17__8_,r_n_17__7_,r_n_17__6_,r_n_17__5_,r_n_17__4_,r_n_17__3_,r_n_17__2_,
  r_n_17__1_,r_n_17__0_,r_n_32__63_,r_n_32__62_,r_n_32__61_,r_n_32__60_,r_n_32__59_,
  r_n_32__58_,r_n_32__57_,r_n_32__56_,r_n_32__55_,r_n_32__54_,r_n_32__53_,r_n_32__52_,
  r_n_32__51_,r_n_32__50_,r_n_32__49_,r_n_32__48_,r_n_32__47_,r_n_32__46_,
  r_n_32__45_,r_n_32__44_,r_n_32__43_,r_n_32__42_,r_n_32__41_,r_n_32__40_,r_n_32__39_,
  r_n_32__38_,r_n_32__37_,r_n_32__36_,r_n_32__35_,r_n_32__34_,r_n_32__33_,r_n_32__32_,
  r_n_32__31_,r_n_32__30_,r_n_32__29_,r_n_32__28_,r_n_32__27_,r_n_32__26_,
  r_n_32__25_,r_n_32__24_,r_n_32__23_,r_n_32__22_,r_n_32__21_,r_n_32__20_,r_n_32__19_,
  r_n_32__18_,r_n_32__17_,r_n_32__16_,r_n_32__15_,r_n_32__14_,r_n_32__13_,r_n_32__12_,
  r_n_32__11_,r_n_32__10_,r_n_32__9_,r_n_32__8_,r_n_32__7_,r_n_32__6_,r_n_32__5_,
  r_n_32__4_,r_n_32__3_,r_n_32__2_,r_n_32__1_,r_n_32__0_,r_n_31__63_,r_n_31__62_,
  r_n_31__61_,r_n_31__60_,r_n_31__59_,r_n_31__58_,r_n_31__57_,r_n_31__56_,r_n_31__55_,
  r_n_31__54_,r_n_31__53_,r_n_31__52_,r_n_31__51_,r_n_31__50_,r_n_31__49_,
  r_n_31__48_,r_n_31__47_,r_n_31__46_,r_n_31__45_,r_n_31__44_,r_n_31__43_,r_n_31__42_,
  r_n_31__41_,r_n_31__40_,r_n_31__39_,r_n_31__38_,r_n_31__37_,r_n_31__36_,r_n_31__35_,
  r_n_31__34_,r_n_31__33_,r_n_31__32_,r_n_31__31_,r_n_31__30_,r_n_31__29_,
  r_n_31__28_,r_n_31__27_,r_n_31__26_,r_n_31__25_,r_n_31__24_,r_n_31__23_,r_n_31__22_,
  r_n_31__21_,r_n_31__20_,r_n_31__19_,r_n_31__18_,r_n_31__17_,r_n_31__16_,r_n_31__15_,
  r_n_31__14_,r_n_31__13_,r_n_31__12_,r_n_31__11_,r_n_31__10_,r_n_31__9_,
  r_n_31__8_,r_n_31__7_,r_n_31__6_,r_n_31__5_,r_n_31__4_,r_n_31__3_,r_n_31__2_,r_n_31__1_,
  r_n_31__0_,r_n_30__63_,r_n_30__62_,r_n_30__61_,r_n_30__60_,r_n_30__59_,
  r_n_30__58_,r_n_30__57_,r_n_30__56_,r_n_30__55_,r_n_30__54_,r_n_30__53_,r_n_30__52_,
  r_n_30__51_,r_n_30__50_,r_n_30__49_,r_n_30__48_,r_n_30__47_,r_n_30__46_,r_n_30__45_,
  r_n_30__44_,r_n_30__43_,r_n_30__42_,r_n_30__41_,r_n_30__40_,r_n_30__39_,
  r_n_30__38_,r_n_30__37_,r_n_30__36_,r_n_30__35_,r_n_30__34_,r_n_30__33_,r_n_30__32_,
  r_n_30__31_,r_n_30__30_,r_n_30__29_,r_n_30__28_,r_n_30__27_,r_n_30__26_,r_n_30__25_,
  r_n_30__24_,r_n_30__23_,r_n_30__22_,r_n_30__21_,r_n_30__20_,r_n_30__19_,
  r_n_30__18_,r_n_30__17_,r_n_30__16_,r_n_30__15_,r_n_30__14_,r_n_30__13_,r_n_30__12_,
  r_n_30__11_,r_n_30__10_,r_n_30__9_,r_n_30__8_,r_n_30__7_,r_n_30__6_,r_n_30__5_,
  r_n_30__4_,r_n_30__3_,r_n_30__2_,r_n_30__1_,r_n_30__0_,r_n_29__63_,r_n_29__62_,
  r_n_29__61_,r_n_29__60_,r_n_29__59_,r_n_29__58_,r_n_29__57_,r_n_29__56_,r_n_29__55_,
  r_n_29__54_,r_n_29__53_,r_n_29__52_,r_n_29__51_,r_n_29__50_,r_n_29__49_,r_n_29__48_,
  r_n_29__47_,r_n_29__46_,r_n_29__45_,r_n_29__44_,r_n_29__43_,r_n_29__42_,
  r_n_29__41_,r_n_29__40_,r_n_29__39_,r_n_29__38_,r_n_29__37_,r_n_29__36_,r_n_29__35_,
  r_n_29__34_,r_n_29__33_,r_n_29__32_,r_n_29__31_,r_n_29__30_,r_n_29__29_,r_n_29__28_,
  r_n_29__27_,r_n_29__26_,r_n_29__25_,r_n_29__24_,r_n_29__23_,r_n_29__22_,
  r_n_29__21_,r_n_29__20_,r_n_29__19_,r_n_29__18_,r_n_29__17_,r_n_29__16_,r_n_29__15_,
  r_n_29__14_,r_n_29__13_,r_n_29__12_,r_n_29__11_,r_n_29__10_,r_n_29__9_,r_n_29__8_,
  r_n_29__7_,r_n_29__6_,r_n_29__5_,r_n_29__4_,r_n_29__3_,r_n_29__2_,r_n_29__1_,
  r_n_29__0_,r_n_28__63_,r_n_28__62_,r_n_28__61_,r_n_28__60_,r_n_28__59_,r_n_28__58_,
  r_n_28__57_,r_n_28__56_,r_n_28__55_,r_n_28__54_,r_n_28__53_,r_n_28__52_,
  r_n_28__51_,r_n_28__50_,r_n_28__49_,r_n_28__48_,r_n_28__47_,r_n_28__46_,r_n_28__45_,
  r_n_28__44_,r_n_28__43_,r_n_28__42_,r_n_28__41_,r_n_28__40_,r_n_28__39_,r_n_28__38_,
  r_n_28__37_,r_n_28__36_,r_n_28__35_,r_n_28__34_,r_n_28__33_,r_n_28__32_,
  r_n_28__31_,r_n_28__30_,r_n_28__29_,r_n_28__28_,r_n_28__27_,r_n_28__26_,r_n_28__25_,
  r_n_28__24_,r_n_28__23_,r_n_28__22_,r_n_28__21_,r_n_28__20_,r_n_28__19_,r_n_28__18_,
  r_n_28__17_,r_n_28__16_,r_n_28__15_,r_n_28__14_,r_n_28__13_,r_n_28__12_,
  r_n_28__11_,r_n_28__10_,r_n_28__9_,r_n_28__8_,r_n_28__7_,r_n_28__6_,r_n_28__5_,r_n_28__4_,
  r_n_28__3_,r_n_28__2_,r_n_28__1_,r_n_28__0_,r_n_27__63_,r_n_27__62_,r_n_27__61_,
  r_n_27__60_,r_n_27__59_,r_n_27__58_,r_n_27__57_,r_n_27__56_,r_n_27__55_,
  r_n_27__54_,r_n_27__53_,r_n_27__52_,r_n_27__51_,r_n_27__50_,r_n_27__49_,r_n_27__48_,
  r_n_27__47_,r_n_27__46_,r_n_27__45_,r_n_27__44_,r_n_27__43_,r_n_27__42_,r_n_27__41_,
  r_n_27__40_,r_n_27__39_,r_n_27__38_,r_n_27__37_,r_n_27__36_,r_n_27__35_,
  r_n_27__34_,r_n_27__33_,r_n_27__32_,r_n_27__31_,r_n_27__30_,r_n_27__29_,r_n_27__28_,
  r_n_27__27_,r_n_27__26_,r_n_27__25_,r_n_27__24_,r_n_27__23_,r_n_27__22_,r_n_27__21_,
  r_n_27__20_,r_n_27__19_,r_n_27__18_,r_n_27__17_,r_n_27__16_,r_n_27__15_,
  r_n_27__14_,r_n_27__13_,r_n_27__12_,r_n_27__11_,r_n_27__10_,r_n_27__9_,r_n_27__8_,
  r_n_27__7_,r_n_27__6_,r_n_27__5_,r_n_27__4_,r_n_27__3_,r_n_27__2_,r_n_27__1_,
  r_n_27__0_,r_n_26__63_,r_n_26__62_,r_n_26__61_,r_n_26__60_,r_n_26__59_,r_n_26__58_,
  r_n_26__57_,r_n_26__56_,r_n_26__55_,r_n_26__54_,r_n_26__53_,r_n_26__52_,r_n_26__51_,
  r_n_26__50_,r_n_26__49_,r_n_26__48_,r_n_26__47_,r_n_26__46_,r_n_26__45_,
  r_n_26__44_,r_n_26__43_,r_n_26__42_,r_n_26__41_,r_n_26__40_,r_n_26__39_,r_n_26__38_,
  r_n_26__37_,r_n_26__36_,r_n_26__35_,r_n_26__34_,r_n_26__33_,r_n_26__32_,r_n_26__31_,
  r_n_26__30_,r_n_26__29_,r_n_26__28_,r_n_26__27_,r_n_26__26_,r_n_26__25_,
  r_n_26__24_,r_n_26__23_,r_n_26__22_,r_n_26__21_,r_n_26__20_,r_n_26__19_,r_n_26__18_,
  r_n_26__17_,r_n_26__16_,r_n_26__15_,r_n_26__14_,r_n_26__13_,r_n_26__12_,r_n_26__11_,
  r_n_26__10_,r_n_26__9_,r_n_26__8_,r_n_26__7_,r_n_26__6_,r_n_26__5_,r_n_26__4_,
  r_n_26__3_,r_n_26__2_,r_n_26__1_,r_n_26__0_,r_n_25__63_,r_n_25__62_,r_n_25__61_,
  r_n_25__60_,r_n_25__59_,r_n_25__58_,r_n_25__57_,r_n_25__56_,r_n_25__55_,r_n_25__54_,
  r_n_25__53_,r_n_25__52_,r_n_25__51_,r_n_25__50_,r_n_25__49_,r_n_25__48_,
  r_n_25__47_,r_n_25__46_,r_n_25__45_,r_n_25__44_,r_n_25__43_,r_n_25__42_,r_n_25__41_,
  r_n_25__40_,r_n_25__39_,r_n_25__38_,r_n_25__37_,r_n_25__36_,r_n_25__35_,r_n_25__34_,
  r_n_25__33_,r_n_25__32_,r_n_25__31_,r_n_25__30_,r_n_25__29_,r_n_25__28_,
  r_n_25__27_,r_n_25__26_,r_n_25__25_,r_n_25__24_,r_n_25__23_,r_n_25__22_,r_n_25__21_,
  r_n_25__20_,r_n_25__19_,r_n_25__18_,r_n_25__17_,r_n_25__16_,r_n_25__15_,r_n_25__14_,
  r_n_25__13_,r_n_25__12_,r_n_25__11_,r_n_25__10_,r_n_25__9_,r_n_25__8_,
  r_n_25__7_,r_n_25__6_,r_n_25__5_,r_n_25__4_,r_n_25__3_,r_n_25__2_,r_n_25__1_,r_n_25__0_,
  r_n_40__63_,r_n_40__62_,r_n_40__61_,r_n_40__60_,r_n_40__59_,r_n_40__58_,
  r_n_40__57_,r_n_40__56_,r_n_40__55_,r_n_40__54_,r_n_40__53_,r_n_40__52_,r_n_40__51_,
  r_n_40__50_,r_n_40__49_,r_n_40__48_,r_n_40__47_,r_n_40__46_,r_n_40__45_,r_n_40__44_,
  r_n_40__43_,r_n_40__42_,r_n_40__41_,r_n_40__40_,r_n_40__39_,r_n_40__38_,
  r_n_40__37_,r_n_40__36_,r_n_40__35_,r_n_40__34_,r_n_40__33_,r_n_40__32_,r_n_40__31_,
  r_n_40__30_,r_n_40__29_,r_n_40__28_,r_n_40__27_,r_n_40__26_,r_n_40__25_,r_n_40__24_,
  r_n_40__23_,r_n_40__22_,r_n_40__21_,r_n_40__20_,r_n_40__19_,r_n_40__18_,
  r_n_40__17_,r_n_40__16_,r_n_40__15_,r_n_40__14_,r_n_40__13_,r_n_40__12_,r_n_40__11_,
  r_n_40__10_,r_n_40__9_,r_n_40__8_,r_n_40__7_,r_n_40__6_,r_n_40__5_,r_n_40__4_,
  r_n_40__3_,r_n_40__2_,r_n_40__1_,r_n_40__0_,r_n_39__63_,r_n_39__62_,r_n_39__61_,
  r_n_39__60_,r_n_39__59_,r_n_39__58_,r_n_39__57_,r_n_39__56_,r_n_39__55_,r_n_39__54_,
  r_n_39__53_,r_n_39__52_,r_n_39__51_,r_n_39__50_,r_n_39__49_,r_n_39__48_,r_n_39__47_,
  r_n_39__46_,r_n_39__45_,r_n_39__44_,r_n_39__43_,r_n_39__42_,r_n_39__41_,
  r_n_39__40_,r_n_39__39_,r_n_39__38_,r_n_39__37_,r_n_39__36_,r_n_39__35_,r_n_39__34_,
  r_n_39__33_,r_n_39__32_,r_n_39__31_,r_n_39__30_,r_n_39__29_,r_n_39__28_,r_n_39__27_,
  r_n_39__26_,r_n_39__25_,r_n_39__24_,r_n_39__23_,r_n_39__22_,r_n_39__21_,
  r_n_39__20_,r_n_39__19_,r_n_39__18_,r_n_39__17_,r_n_39__16_,r_n_39__15_,r_n_39__14_,
  r_n_39__13_,r_n_39__12_,r_n_39__11_,r_n_39__10_,r_n_39__9_,r_n_39__8_,r_n_39__7_,
  r_n_39__6_,r_n_39__5_,r_n_39__4_,r_n_39__3_,r_n_39__2_,r_n_39__1_,r_n_39__0_,
  r_n_38__63_,r_n_38__62_,r_n_38__61_,r_n_38__60_,r_n_38__59_,r_n_38__58_,r_n_38__57_,
  r_n_38__56_,r_n_38__55_,r_n_38__54_,r_n_38__53_,r_n_38__52_,r_n_38__51_,
  r_n_38__50_,r_n_38__49_,r_n_38__48_,r_n_38__47_,r_n_38__46_,r_n_38__45_,r_n_38__44_,
  r_n_38__43_,r_n_38__42_,r_n_38__41_,r_n_38__40_,r_n_38__39_,r_n_38__38_,r_n_38__37_,
  r_n_38__36_,r_n_38__35_,r_n_38__34_,r_n_38__33_,r_n_38__32_,r_n_38__31_,
  r_n_38__30_,r_n_38__29_,r_n_38__28_,r_n_38__27_,r_n_38__26_,r_n_38__25_,r_n_38__24_,
  r_n_38__23_,r_n_38__22_,r_n_38__21_,r_n_38__20_,r_n_38__19_,r_n_38__18_,r_n_38__17_,
  r_n_38__16_,r_n_38__15_,r_n_38__14_,r_n_38__13_,r_n_38__12_,r_n_38__11_,
  r_n_38__10_,r_n_38__9_,r_n_38__8_,r_n_38__7_,r_n_38__6_,r_n_38__5_,r_n_38__4_,r_n_38__3_,
  r_n_38__2_,r_n_38__1_,r_n_38__0_,r_n_37__63_,r_n_37__62_,r_n_37__61_,r_n_37__60_,
  r_n_37__59_,r_n_37__58_,r_n_37__57_,r_n_37__56_,r_n_37__55_,r_n_37__54_,
  r_n_37__53_,r_n_37__52_,r_n_37__51_,r_n_37__50_,r_n_37__49_,r_n_37__48_,r_n_37__47_,
  r_n_37__46_,r_n_37__45_,r_n_37__44_,r_n_37__43_,r_n_37__42_,r_n_37__41_,r_n_37__40_,
  r_n_37__39_,r_n_37__38_,r_n_37__37_,r_n_37__36_,r_n_37__35_,r_n_37__34_,
  r_n_37__33_,r_n_37__32_,r_n_37__31_,r_n_37__30_,r_n_37__29_,r_n_37__28_,r_n_37__27_,
  r_n_37__26_,r_n_37__25_,r_n_37__24_,r_n_37__23_,r_n_37__22_,r_n_37__21_,r_n_37__20_,
  r_n_37__19_,r_n_37__18_,r_n_37__17_,r_n_37__16_,r_n_37__15_,r_n_37__14_,
  r_n_37__13_,r_n_37__12_,r_n_37__11_,r_n_37__10_,r_n_37__9_,r_n_37__8_,r_n_37__7_,
  r_n_37__6_,r_n_37__5_,r_n_37__4_,r_n_37__3_,r_n_37__2_,r_n_37__1_,r_n_37__0_,
  r_n_36__63_,r_n_36__62_,r_n_36__61_,r_n_36__60_,r_n_36__59_,r_n_36__58_,r_n_36__57_,
  r_n_36__56_,r_n_36__55_,r_n_36__54_,r_n_36__53_,r_n_36__52_,r_n_36__51_,r_n_36__50_,
  r_n_36__49_,r_n_36__48_,r_n_36__47_,r_n_36__46_,r_n_36__45_,r_n_36__44_,
  r_n_36__43_,r_n_36__42_,r_n_36__41_,r_n_36__40_,r_n_36__39_,r_n_36__38_,r_n_36__37_,
  r_n_36__36_,r_n_36__35_,r_n_36__34_,r_n_36__33_,r_n_36__32_,r_n_36__31_,r_n_36__30_,
  r_n_36__29_,r_n_36__28_,r_n_36__27_,r_n_36__26_,r_n_36__25_,r_n_36__24_,
  r_n_36__23_,r_n_36__22_,r_n_36__21_,r_n_36__20_,r_n_36__19_,r_n_36__18_,r_n_36__17_,
  r_n_36__16_,r_n_36__15_,r_n_36__14_,r_n_36__13_,r_n_36__12_,r_n_36__11_,r_n_36__10_,
  r_n_36__9_,r_n_36__8_,r_n_36__7_,r_n_36__6_,r_n_36__5_,r_n_36__4_,r_n_36__3_,
  r_n_36__2_,r_n_36__1_,r_n_36__0_,r_n_35__63_,r_n_35__62_,r_n_35__61_,r_n_35__60_,
  r_n_35__59_,r_n_35__58_,r_n_35__57_,r_n_35__56_,r_n_35__55_,r_n_35__54_,r_n_35__53_,
  r_n_35__52_,r_n_35__51_,r_n_35__50_,r_n_35__49_,r_n_35__48_,r_n_35__47_,
  r_n_35__46_,r_n_35__45_,r_n_35__44_,r_n_35__43_,r_n_35__42_,r_n_35__41_,r_n_35__40_,
  r_n_35__39_,r_n_35__38_,r_n_35__37_,r_n_35__36_,r_n_35__35_,r_n_35__34_,r_n_35__33_,
  r_n_35__32_,r_n_35__31_,r_n_35__30_,r_n_35__29_,r_n_35__28_,r_n_35__27_,
  r_n_35__26_,r_n_35__25_,r_n_35__24_,r_n_35__23_,r_n_35__22_,r_n_35__21_,r_n_35__20_,
  r_n_35__19_,r_n_35__18_,r_n_35__17_,r_n_35__16_,r_n_35__15_,r_n_35__14_,r_n_35__13_,
  r_n_35__12_,r_n_35__11_,r_n_35__10_,r_n_35__9_,r_n_35__8_,r_n_35__7_,r_n_35__6_,
  r_n_35__5_,r_n_35__4_,r_n_35__3_,r_n_35__2_,r_n_35__1_,r_n_35__0_,r_n_34__63_,
  r_n_34__62_,r_n_34__61_,r_n_34__60_,r_n_34__59_,r_n_34__58_,r_n_34__57_,
  r_n_34__56_,r_n_34__55_,r_n_34__54_,r_n_34__53_,r_n_34__52_,r_n_34__51_,r_n_34__50_,
  r_n_34__49_,r_n_34__48_,r_n_34__47_,r_n_34__46_,r_n_34__45_,r_n_34__44_,r_n_34__43_,
  r_n_34__42_,r_n_34__41_,r_n_34__40_,r_n_34__39_,r_n_34__38_,r_n_34__37_,
  r_n_34__36_,r_n_34__35_,r_n_34__34_,r_n_34__33_,r_n_34__32_,r_n_34__31_,r_n_34__30_,
  r_n_34__29_,r_n_34__28_,r_n_34__27_,r_n_34__26_,r_n_34__25_,r_n_34__24_,r_n_34__23_,
  r_n_34__22_,r_n_34__21_,r_n_34__20_,r_n_34__19_,r_n_34__18_,r_n_34__17_,
  r_n_34__16_,r_n_34__15_,r_n_34__14_,r_n_34__13_,r_n_34__12_,r_n_34__11_,r_n_34__10_,
  r_n_34__9_,r_n_34__8_,r_n_34__7_,r_n_34__6_,r_n_34__5_,r_n_34__4_,r_n_34__3_,
  r_n_34__2_,r_n_34__1_,r_n_34__0_,r_n_33__63_,r_n_33__62_,r_n_33__61_,r_n_33__60_,
  r_n_33__59_,r_n_33__58_,r_n_33__57_,r_n_33__56_,r_n_33__55_,r_n_33__54_,r_n_33__53_,
  r_n_33__52_,r_n_33__51_,r_n_33__50_,r_n_33__49_,r_n_33__48_,r_n_33__47_,r_n_33__46_,
  r_n_33__45_,r_n_33__44_,r_n_33__43_,r_n_33__42_,r_n_33__41_,r_n_33__40_,
  r_n_33__39_,r_n_33__38_,r_n_33__37_,r_n_33__36_,r_n_33__35_,r_n_33__34_,r_n_33__33_,
  r_n_33__32_,r_n_33__31_,r_n_33__30_,r_n_33__29_,r_n_33__28_,r_n_33__27_,r_n_33__26_,
  r_n_33__25_,r_n_33__24_,r_n_33__23_,r_n_33__22_,r_n_33__21_,r_n_33__20_,
  r_n_33__19_,r_n_33__18_,r_n_33__17_,r_n_33__16_,r_n_33__15_,r_n_33__14_,r_n_33__13_,
  r_n_33__12_,r_n_33__11_,r_n_33__10_,r_n_33__9_,r_n_33__8_,r_n_33__7_,r_n_33__6_,
  r_n_33__5_,r_n_33__4_,r_n_33__3_,r_n_33__2_,r_n_33__1_,r_n_33__0_,r_n_48__63_,
  r_n_48__62_,r_n_48__61_,r_n_48__60_,r_n_48__59_,r_n_48__58_,r_n_48__57_,r_n_48__56_,
  r_n_48__55_,r_n_48__54_,r_n_48__53_,r_n_48__52_,r_n_48__51_,r_n_48__50_,
  r_n_48__49_,r_n_48__48_,r_n_48__47_,r_n_48__46_,r_n_48__45_,r_n_48__44_,r_n_48__43_,
  r_n_48__42_,r_n_48__41_,r_n_48__40_,r_n_48__39_,r_n_48__38_,r_n_48__37_,r_n_48__36_,
  r_n_48__35_,r_n_48__34_,r_n_48__33_,r_n_48__32_,r_n_48__31_,r_n_48__30_,
  r_n_48__29_,r_n_48__28_,r_n_48__27_,r_n_48__26_,r_n_48__25_,r_n_48__24_,r_n_48__23_,
  r_n_48__22_,r_n_48__21_,r_n_48__20_,r_n_48__19_,r_n_48__18_,r_n_48__17_,r_n_48__16_,
  r_n_48__15_,r_n_48__14_,r_n_48__13_,r_n_48__12_,r_n_48__11_,r_n_48__10_,
  r_n_48__9_,r_n_48__8_,r_n_48__7_,r_n_48__6_,r_n_48__5_,r_n_48__4_,r_n_48__3_,r_n_48__2_,
  r_n_48__1_,r_n_48__0_,r_n_47__63_,r_n_47__62_,r_n_47__61_,r_n_47__60_,r_n_47__59_,
  r_n_47__58_,r_n_47__57_,r_n_47__56_,r_n_47__55_,r_n_47__54_,r_n_47__53_,
  r_n_47__52_,r_n_47__51_,r_n_47__50_,r_n_47__49_,r_n_47__48_,r_n_47__47_,r_n_47__46_,
  r_n_47__45_,r_n_47__44_,r_n_47__43_,r_n_47__42_,r_n_47__41_,r_n_47__40_,r_n_47__39_,
  r_n_47__38_,r_n_47__37_,r_n_47__36_,r_n_47__35_,r_n_47__34_,r_n_47__33_,
  r_n_47__32_,r_n_47__31_,r_n_47__30_,r_n_47__29_,r_n_47__28_,r_n_47__27_,r_n_47__26_,
  r_n_47__25_,r_n_47__24_,r_n_47__23_,r_n_47__22_,r_n_47__21_,r_n_47__20_,r_n_47__19_,
  r_n_47__18_,r_n_47__17_,r_n_47__16_,r_n_47__15_,r_n_47__14_,r_n_47__13_,
  r_n_47__12_,r_n_47__11_,r_n_47__10_,r_n_47__9_,r_n_47__8_,r_n_47__7_,r_n_47__6_,
  r_n_47__5_,r_n_47__4_,r_n_47__3_,r_n_47__2_,r_n_47__1_,r_n_47__0_,r_n_46__63_,
  r_n_46__62_,r_n_46__61_,r_n_46__60_,r_n_46__59_,r_n_46__58_,r_n_46__57_,r_n_46__56_,
  r_n_46__55_,r_n_46__54_,r_n_46__53_,r_n_46__52_,r_n_46__51_,r_n_46__50_,r_n_46__49_,
  r_n_46__48_,r_n_46__47_,r_n_46__46_,r_n_46__45_,r_n_46__44_,r_n_46__43_,
  r_n_46__42_,r_n_46__41_,r_n_46__40_,r_n_46__39_,r_n_46__38_,r_n_46__37_,r_n_46__36_,
  r_n_46__35_,r_n_46__34_,r_n_46__33_,r_n_46__32_,r_n_46__31_,r_n_46__30_,r_n_46__29_,
  r_n_46__28_,r_n_46__27_,r_n_46__26_,r_n_46__25_,r_n_46__24_,r_n_46__23_,
  r_n_46__22_,r_n_46__21_,r_n_46__20_,r_n_46__19_,r_n_46__18_,r_n_46__17_,r_n_46__16_,
  r_n_46__15_,r_n_46__14_,r_n_46__13_,r_n_46__12_,r_n_46__11_,r_n_46__10_,r_n_46__9_,
  r_n_46__8_,r_n_46__7_,r_n_46__6_,r_n_46__5_,r_n_46__4_,r_n_46__3_,r_n_46__2_,
  r_n_46__1_,r_n_46__0_,r_n_45__63_,r_n_45__62_,r_n_45__61_,r_n_45__60_,r_n_45__59_,
  r_n_45__58_,r_n_45__57_,r_n_45__56_,r_n_45__55_,r_n_45__54_,r_n_45__53_,r_n_45__52_,
  r_n_45__51_,r_n_45__50_,r_n_45__49_,r_n_45__48_,r_n_45__47_,r_n_45__46_,
  r_n_45__45_,r_n_45__44_,r_n_45__43_,r_n_45__42_,r_n_45__41_,r_n_45__40_,r_n_45__39_,
  r_n_45__38_,r_n_45__37_,r_n_45__36_,r_n_45__35_,r_n_45__34_,r_n_45__33_,r_n_45__32_,
  r_n_45__31_,r_n_45__30_,r_n_45__29_,r_n_45__28_,r_n_45__27_,r_n_45__26_,
  r_n_45__25_,r_n_45__24_,r_n_45__23_,r_n_45__22_,r_n_45__21_,r_n_45__20_,r_n_45__19_,
  r_n_45__18_,r_n_45__17_,r_n_45__16_,r_n_45__15_,r_n_45__14_,r_n_45__13_,r_n_45__12_,
  r_n_45__11_,r_n_45__10_,r_n_45__9_,r_n_45__8_,r_n_45__7_,r_n_45__6_,r_n_45__5_,
  r_n_45__4_,r_n_45__3_,r_n_45__2_,r_n_45__1_,r_n_45__0_,r_n_44__63_,r_n_44__62_,
  r_n_44__61_,r_n_44__60_,r_n_44__59_,r_n_44__58_,r_n_44__57_,r_n_44__56_,
  r_n_44__55_,r_n_44__54_,r_n_44__53_,r_n_44__52_,r_n_44__51_,r_n_44__50_,r_n_44__49_,
  r_n_44__48_,r_n_44__47_,r_n_44__46_,r_n_44__45_,r_n_44__44_,r_n_44__43_,r_n_44__42_,
  r_n_44__41_,r_n_44__40_,r_n_44__39_,r_n_44__38_,r_n_44__37_,r_n_44__36_,
  r_n_44__35_,r_n_44__34_,r_n_44__33_,r_n_44__32_,r_n_44__31_,r_n_44__30_,r_n_44__29_,
  r_n_44__28_,r_n_44__27_,r_n_44__26_,r_n_44__25_,r_n_44__24_,r_n_44__23_,r_n_44__22_,
  r_n_44__21_,r_n_44__20_,r_n_44__19_,r_n_44__18_,r_n_44__17_,r_n_44__16_,
  r_n_44__15_,r_n_44__14_,r_n_44__13_,r_n_44__12_,r_n_44__11_,r_n_44__10_,r_n_44__9_,
  r_n_44__8_,r_n_44__7_,r_n_44__6_,r_n_44__5_,r_n_44__4_,r_n_44__3_,r_n_44__2_,
  r_n_44__1_,r_n_44__0_,r_n_43__63_,r_n_43__62_,r_n_43__61_,r_n_43__60_,r_n_43__59_,
  r_n_43__58_,r_n_43__57_,r_n_43__56_,r_n_43__55_,r_n_43__54_,r_n_43__53_,r_n_43__52_,
  r_n_43__51_,r_n_43__50_,r_n_43__49_,r_n_43__48_,r_n_43__47_,r_n_43__46_,r_n_43__45_,
  r_n_43__44_,r_n_43__43_,r_n_43__42_,r_n_43__41_,r_n_43__40_,r_n_43__39_,
  r_n_43__38_,r_n_43__37_,r_n_43__36_,r_n_43__35_,r_n_43__34_,r_n_43__33_,r_n_43__32_,
  r_n_43__31_,r_n_43__30_,r_n_43__29_,r_n_43__28_,r_n_43__27_,r_n_43__26_,r_n_43__25_,
  r_n_43__24_,r_n_43__23_,r_n_43__22_,r_n_43__21_,r_n_43__20_,r_n_43__19_,
  r_n_43__18_,r_n_43__17_,r_n_43__16_,r_n_43__15_,r_n_43__14_,r_n_43__13_,r_n_43__12_,
  r_n_43__11_,r_n_43__10_,r_n_43__9_,r_n_43__8_,r_n_43__7_,r_n_43__6_,r_n_43__5_,
  r_n_43__4_,r_n_43__3_,r_n_43__2_,r_n_43__1_,r_n_43__0_,r_n_42__63_,r_n_42__62_,
  r_n_42__61_,r_n_42__60_,r_n_42__59_,r_n_42__58_,r_n_42__57_,r_n_42__56_,r_n_42__55_,
  r_n_42__54_,r_n_42__53_,r_n_42__52_,r_n_42__51_,r_n_42__50_,r_n_42__49_,
  r_n_42__48_,r_n_42__47_,r_n_42__46_,r_n_42__45_,r_n_42__44_,r_n_42__43_,r_n_42__42_,
  r_n_42__41_,r_n_42__40_,r_n_42__39_,r_n_42__38_,r_n_42__37_,r_n_42__36_,r_n_42__35_,
  r_n_42__34_,r_n_42__33_,r_n_42__32_,r_n_42__31_,r_n_42__30_,r_n_42__29_,
  r_n_42__28_,r_n_42__27_,r_n_42__26_,r_n_42__25_,r_n_42__24_,r_n_42__23_,r_n_42__22_,
  r_n_42__21_,r_n_42__20_,r_n_42__19_,r_n_42__18_,r_n_42__17_,r_n_42__16_,r_n_42__15_,
  r_n_42__14_,r_n_42__13_,r_n_42__12_,r_n_42__11_,r_n_42__10_,r_n_42__9_,r_n_42__8_,
  r_n_42__7_,r_n_42__6_,r_n_42__5_,r_n_42__4_,r_n_42__3_,r_n_42__2_,r_n_42__1_,
  r_n_42__0_,r_n_41__63_,r_n_41__62_,r_n_41__61_,r_n_41__60_,r_n_41__59_,r_n_41__58_,
  r_n_41__57_,r_n_41__56_,r_n_41__55_,r_n_41__54_,r_n_41__53_,r_n_41__52_,
  r_n_41__51_,r_n_41__50_,r_n_41__49_,r_n_41__48_,r_n_41__47_,r_n_41__46_,r_n_41__45_,
  r_n_41__44_,r_n_41__43_,r_n_41__42_,r_n_41__41_,r_n_41__40_,r_n_41__39_,r_n_41__38_,
  r_n_41__37_,r_n_41__36_,r_n_41__35_,r_n_41__34_,r_n_41__33_,r_n_41__32_,
  r_n_41__31_,r_n_41__30_,r_n_41__29_,r_n_41__28_,r_n_41__27_,r_n_41__26_,r_n_41__25_,
  r_n_41__24_,r_n_41__23_,r_n_41__22_,r_n_41__21_,r_n_41__20_,r_n_41__19_,r_n_41__18_,
  r_n_41__17_,r_n_41__16_,r_n_41__15_,r_n_41__14_,r_n_41__13_,r_n_41__12_,
  r_n_41__11_,r_n_41__10_,r_n_41__9_,r_n_41__8_,r_n_41__7_,r_n_41__6_,r_n_41__5_,
  r_n_41__4_,r_n_41__3_,r_n_41__2_,r_n_41__1_,r_n_41__0_,r_n_56__63_,r_n_56__62_,
  r_n_56__61_,r_n_56__60_,r_n_56__59_,r_n_56__58_,r_n_56__57_,r_n_56__56_,r_n_56__55_,
  r_n_56__54_,r_n_56__53_,r_n_56__52_,r_n_56__51_,r_n_56__50_,r_n_56__49_,r_n_56__48_,
  r_n_56__47_,r_n_56__46_,r_n_56__45_,r_n_56__44_,r_n_56__43_,r_n_56__42_,
  r_n_56__41_,r_n_56__40_,r_n_56__39_,r_n_56__38_,r_n_56__37_,r_n_56__36_,r_n_56__35_,
  r_n_56__34_,r_n_56__33_,r_n_56__32_,r_n_56__31_,r_n_56__30_,r_n_56__29_,r_n_56__28_,
  r_n_56__27_,r_n_56__26_,r_n_56__25_,r_n_56__24_,r_n_56__23_,r_n_56__22_,
  r_n_56__21_,r_n_56__20_,r_n_56__19_,r_n_56__18_,r_n_56__17_,r_n_56__16_,r_n_56__15_,
  r_n_56__14_,r_n_56__13_,r_n_56__12_,r_n_56__11_,r_n_56__10_,r_n_56__9_,r_n_56__8_,
  r_n_56__7_,r_n_56__6_,r_n_56__5_,r_n_56__4_,r_n_56__3_,r_n_56__2_,r_n_56__1_,
  r_n_56__0_,r_n_55__63_,r_n_55__62_,r_n_55__61_,r_n_55__60_,r_n_55__59_,r_n_55__58_,
  r_n_55__57_,r_n_55__56_,r_n_55__55_,r_n_55__54_,r_n_55__53_,r_n_55__52_,r_n_55__51_,
  r_n_55__50_,r_n_55__49_,r_n_55__48_,r_n_55__47_,r_n_55__46_,r_n_55__45_,
  r_n_55__44_,r_n_55__43_,r_n_55__42_,r_n_55__41_,r_n_55__40_,r_n_55__39_,r_n_55__38_,
  r_n_55__37_,r_n_55__36_,r_n_55__35_,r_n_55__34_,r_n_55__33_,r_n_55__32_,r_n_55__31_,
  r_n_55__30_,r_n_55__29_,r_n_55__28_,r_n_55__27_,r_n_55__26_,r_n_55__25_,
  r_n_55__24_,r_n_55__23_,r_n_55__22_,r_n_55__21_,r_n_55__20_,r_n_55__19_,r_n_55__18_,
  r_n_55__17_,r_n_55__16_,r_n_55__15_,r_n_55__14_,r_n_55__13_,r_n_55__12_,r_n_55__11_,
  r_n_55__10_,r_n_55__9_,r_n_55__8_,r_n_55__7_,r_n_55__6_,r_n_55__5_,r_n_55__4_,
  r_n_55__3_,r_n_55__2_,r_n_55__1_,r_n_55__0_,r_n_54__63_,r_n_54__62_,r_n_54__61_,
  r_n_54__60_,r_n_54__59_,r_n_54__58_,r_n_54__57_,r_n_54__56_,r_n_54__55_,
  r_n_54__54_,r_n_54__53_,r_n_54__52_,r_n_54__51_,r_n_54__50_,r_n_54__49_,r_n_54__48_,
  r_n_54__47_,r_n_54__46_,r_n_54__45_,r_n_54__44_,r_n_54__43_,r_n_54__42_,r_n_54__41_,
  r_n_54__40_,r_n_54__39_,r_n_54__38_,r_n_54__37_,r_n_54__36_,r_n_54__35_,
  r_n_54__34_,r_n_54__33_,r_n_54__32_,r_n_54__31_,r_n_54__30_,r_n_54__29_,r_n_54__28_,
  r_n_54__27_,r_n_54__26_,r_n_54__25_,r_n_54__24_,r_n_54__23_,r_n_54__22_,r_n_54__21_,
  r_n_54__20_,r_n_54__19_,r_n_54__18_,r_n_54__17_,r_n_54__16_,r_n_54__15_,
  r_n_54__14_,r_n_54__13_,r_n_54__12_,r_n_54__11_,r_n_54__10_,r_n_54__9_,r_n_54__8_,
  r_n_54__7_,r_n_54__6_,r_n_54__5_,r_n_54__4_,r_n_54__3_,r_n_54__2_,r_n_54__1_,r_n_54__0_,
  r_n_53__63_,r_n_53__62_,r_n_53__61_,r_n_53__60_,r_n_53__59_,r_n_53__58_,
  r_n_53__57_,r_n_53__56_,r_n_53__55_,r_n_53__54_,r_n_53__53_,r_n_53__52_,r_n_53__51_,
  r_n_53__50_,r_n_53__49_,r_n_53__48_,r_n_53__47_,r_n_53__46_,r_n_53__45_,r_n_53__44_,
  r_n_53__43_,r_n_53__42_,r_n_53__41_,r_n_53__40_,r_n_53__39_,r_n_53__38_,
  r_n_53__37_,r_n_53__36_,r_n_53__35_,r_n_53__34_,r_n_53__33_,r_n_53__32_,r_n_53__31_,
  r_n_53__30_,r_n_53__29_,r_n_53__28_,r_n_53__27_,r_n_53__26_,r_n_53__25_,r_n_53__24_,
  r_n_53__23_,r_n_53__22_,r_n_53__21_,r_n_53__20_,r_n_53__19_,r_n_53__18_,
  r_n_53__17_,r_n_53__16_,r_n_53__15_,r_n_53__14_,r_n_53__13_,r_n_53__12_,r_n_53__11_,
  r_n_53__10_,r_n_53__9_,r_n_53__8_,r_n_53__7_,r_n_53__6_,r_n_53__5_,r_n_53__4_,
  r_n_53__3_,r_n_53__2_,r_n_53__1_,r_n_53__0_,r_n_52__63_,r_n_52__62_,r_n_52__61_,
  r_n_52__60_,r_n_52__59_,r_n_52__58_,r_n_52__57_,r_n_52__56_,r_n_52__55_,r_n_52__54_,
  r_n_52__53_,r_n_52__52_,r_n_52__51_,r_n_52__50_,r_n_52__49_,r_n_52__48_,
  r_n_52__47_,r_n_52__46_,r_n_52__45_,r_n_52__44_,r_n_52__43_,r_n_52__42_,r_n_52__41_,
  r_n_52__40_,r_n_52__39_,r_n_52__38_,r_n_52__37_,r_n_52__36_,r_n_52__35_,r_n_52__34_,
  r_n_52__33_,r_n_52__32_,r_n_52__31_,r_n_52__30_,r_n_52__29_,r_n_52__28_,
  r_n_52__27_,r_n_52__26_,r_n_52__25_,r_n_52__24_,r_n_52__23_,r_n_52__22_,r_n_52__21_,
  r_n_52__20_,r_n_52__19_,r_n_52__18_,r_n_52__17_,r_n_52__16_,r_n_52__15_,r_n_52__14_,
  r_n_52__13_,r_n_52__12_,r_n_52__11_,r_n_52__10_,r_n_52__9_,r_n_52__8_,r_n_52__7_,
  r_n_52__6_,r_n_52__5_,r_n_52__4_,r_n_52__3_,r_n_52__2_,r_n_52__1_,r_n_52__0_,
  r_n_51__63_,r_n_51__62_,r_n_51__61_,r_n_51__60_,r_n_51__59_,r_n_51__58_,r_n_51__57_,
  r_n_51__56_,r_n_51__55_,r_n_51__54_,r_n_51__53_,r_n_51__52_,r_n_51__51_,
  r_n_51__50_,r_n_51__49_,r_n_51__48_,r_n_51__47_,r_n_51__46_,r_n_51__45_,r_n_51__44_,
  r_n_51__43_,r_n_51__42_,r_n_51__41_,r_n_51__40_,r_n_51__39_,r_n_51__38_,r_n_51__37_,
  r_n_51__36_,r_n_51__35_,r_n_51__34_,r_n_51__33_,r_n_51__32_,r_n_51__31_,
  r_n_51__30_,r_n_51__29_,r_n_51__28_,r_n_51__27_,r_n_51__26_,r_n_51__25_,r_n_51__24_,
  r_n_51__23_,r_n_51__22_,r_n_51__21_,r_n_51__20_,r_n_51__19_,r_n_51__18_,r_n_51__17_,
  r_n_51__16_,r_n_51__15_,r_n_51__14_,r_n_51__13_,r_n_51__12_,r_n_51__11_,
  r_n_51__10_,r_n_51__9_,r_n_51__8_,r_n_51__7_,r_n_51__6_,r_n_51__5_,r_n_51__4_,
  r_n_51__3_,r_n_51__2_,r_n_51__1_,r_n_51__0_,r_n_50__63_,r_n_50__62_,r_n_50__61_,
  r_n_50__60_,r_n_50__59_,r_n_50__58_,r_n_50__57_,r_n_50__56_,r_n_50__55_,r_n_50__54_,
  r_n_50__53_,r_n_50__52_,r_n_50__51_,r_n_50__50_,r_n_50__49_,r_n_50__48_,r_n_50__47_,
  r_n_50__46_,r_n_50__45_,r_n_50__44_,r_n_50__43_,r_n_50__42_,r_n_50__41_,
  r_n_50__40_,r_n_50__39_,r_n_50__38_,r_n_50__37_,r_n_50__36_,r_n_50__35_,r_n_50__34_,
  r_n_50__33_,r_n_50__32_,r_n_50__31_,r_n_50__30_,r_n_50__29_,r_n_50__28_,r_n_50__27_,
  r_n_50__26_,r_n_50__25_,r_n_50__24_,r_n_50__23_,r_n_50__22_,r_n_50__21_,
  r_n_50__20_,r_n_50__19_,r_n_50__18_,r_n_50__17_,r_n_50__16_,r_n_50__15_,r_n_50__14_,
  r_n_50__13_,r_n_50__12_,r_n_50__11_,r_n_50__10_,r_n_50__9_,r_n_50__8_,r_n_50__7_,
  r_n_50__6_,r_n_50__5_,r_n_50__4_,r_n_50__3_,r_n_50__2_,r_n_50__1_,r_n_50__0_,
  r_n_49__63_,r_n_49__62_,r_n_49__61_,r_n_49__60_,r_n_49__59_,r_n_49__58_,r_n_49__57_,
  r_n_49__56_,r_n_49__55_,r_n_49__54_,r_n_49__53_,r_n_49__52_,r_n_49__51_,r_n_49__50_,
  r_n_49__49_,r_n_49__48_,r_n_49__47_,r_n_49__46_,r_n_49__45_,r_n_49__44_,
  r_n_49__43_,r_n_49__42_,r_n_49__41_,r_n_49__40_,r_n_49__39_,r_n_49__38_,r_n_49__37_,
  r_n_49__36_,r_n_49__35_,r_n_49__34_,r_n_49__33_,r_n_49__32_,r_n_49__31_,r_n_49__30_,
  r_n_49__29_,r_n_49__28_,r_n_49__27_,r_n_49__26_,r_n_49__25_,r_n_49__24_,
  r_n_49__23_,r_n_49__22_,r_n_49__21_,r_n_49__20_,r_n_49__19_,r_n_49__18_,r_n_49__17_,
  r_n_49__16_,r_n_49__15_,r_n_49__14_,r_n_49__13_,r_n_49__12_,r_n_49__11_,r_n_49__10_,
  r_n_49__9_,r_n_49__8_,r_n_49__7_,r_n_49__6_,r_n_49__5_,r_n_49__4_,r_n_49__3_,
  r_n_49__2_,r_n_49__1_,r_n_49__0_,r_n_64__63_,r_n_64__62_,r_n_64__61_,r_n_64__60_,
  r_n_64__59_,r_n_64__58_,r_n_64__57_,r_n_64__56_,r_n_64__55_,r_n_64__54_,
  r_n_64__53_,r_n_64__52_,r_n_64__51_,r_n_64__50_,r_n_64__49_,r_n_64__48_,r_n_64__47_,
  r_n_64__46_,r_n_64__45_,r_n_64__44_,r_n_64__43_,r_n_64__42_,r_n_64__41_,r_n_64__40_,
  r_n_64__39_,r_n_64__38_,r_n_64__37_,r_n_64__36_,r_n_64__35_,r_n_64__34_,
  r_n_64__33_,r_n_64__32_,r_n_64__31_,r_n_64__30_,r_n_64__29_,r_n_64__28_,r_n_64__27_,
  r_n_64__26_,r_n_64__25_,r_n_64__24_,r_n_64__23_,r_n_64__22_,r_n_64__21_,r_n_64__20_,
  r_n_64__19_,r_n_64__18_,r_n_64__17_,r_n_64__16_,r_n_64__15_,r_n_64__14_,
  r_n_64__13_,r_n_64__12_,r_n_64__11_,r_n_64__10_,r_n_64__9_,r_n_64__8_,r_n_64__7_,
  r_n_64__6_,r_n_64__5_,r_n_64__4_,r_n_64__3_,r_n_64__2_,r_n_64__1_,r_n_64__0_,r_n_63__63_,
  r_n_63__62_,r_n_63__61_,r_n_63__60_,r_n_63__59_,r_n_63__58_,r_n_63__57_,
  r_n_63__56_,r_n_63__55_,r_n_63__54_,r_n_63__53_,r_n_63__52_,r_n_63__51_,r_n_63__50_,
  r_n_63__49_,r_n_63__48_,r_n_63__47_,r_n_63__46_,r_n_63__45_,r_n_63__44_,r_n_63__43_,
  r_n_63__42_,r_n_63__41_,r_n_63__40_,r_n_63__39_,r_n_63__38_,r_n_63__37_,
  r_n_63__36_,r_n_63__35_,r_n_63__34_,r_n_63__33_,r_n_63__32_,r_n_63__31_,r_n_63__30_,
  r_n_63__29_,r_n_63__28_,r_n_63__27_,r_n_63__26_,r_n_63__25_,r_n_63__24_,r_n_63__23_,
  r_n_63__22_,r_n_63__21_,r_n_63__20_,r_n_63__19_,r_n_63__18_,r_n_63__17_,
  r_n_63__16_,r_n_63__15_,r_n_63__14_,r_n_63__13_,r_n_63__12_,r_n_63__11_,r_n_63__10_,
  r_n_63__9_,r_n_63__8_,r_n_63__7_,r_n_63__6_,r_n_63__5_,r_n_63__4_,r_n_63__3_,
  r_n_63__2_,r_n_63__1_,r_n_63__0_,r_n_62__63_,r_n_62__62_,r_n_62__61_,r_n_62__60_,
  r_n_62__59_,r_n_62__58_,r_n_62__57_,r_n_62__56_,r_n_62__55_,r_n_62__54_,r_n_62__53_,
  r_n_62__52_,r_n_62__51_,r_n_62__50_,r_n_62__49_,r_n_62__48_,r_n_62__47_,
  r_n_62__46_,r_n_62__45_,r_n_62__44_,r_n_62__43_,r_n_62__42_,r_n_62__41_,r_n_62__40_,
  r_n_62__39_,r_n_62__38_,r_n_62__37_,r_n_62__36_,r_n_62__35_,r_n_62__34_,r_n_62__33_,
  r_n_62__32_,r_n_62__31_,r_n_62__30_,r_n_62__29_,r_n_62__28_,r_n_62__27_,
  r_n_62__26_,r_n_62__25_,r_n_62__24_,r_n_62__23_,r_n_62__22_,r_n_62__21_,r_n_62__20_,
  r_n_62__19_,r_n_62__18_,r_n_62__17_,r_n_62__16_,r_n_62__15_,r_n_62__14_,r_n_62__13_,
  r_n_62__12_,r_n_62__11_,r_n_62__10_,r_n_62__9_,r_n_62__8_,r_n_62__7_,r_n_62__6_,
  r_n_62__5_,r_n_62__4_,r_n_62__3_,r_n_62__2_,r_n_62__1_,r_n_62__0_,r_n_61__63_,
  r_n_61__62_,r_n_61__61_,r_n_61__60_,r_n_61__59_,r_n_61__58_,r_n_61__57_,r_n_61__56_,
  r_n_61__55_,r_n_61__54_,r_n_61__53_,r_n_61__52_,r_n_61__51_,r_n_61__50_,
  r_n_61__49_,r_n_61__48_,r_n_61__47_,r_n_61__46_,r_n_61__45_,r_n_61__44_,r_n_61__43_,
  r_n_61__42_,r_n_61__41_,r_n_61__40_,r_n_61__39_,r_n_61__38_,r_n_61__37_,r_n_61__36_,
  r_n_61__35_,r_n_61__34_,r_n_61__33_,r_n_61__32_,r_n_61__31_,r_n_61__30_,
  r_n_61__29_,r_n_61__28_,r_n_61__27_,r_n_61__26_,r_n_61__25_,r_n_61__24_,r_n_61__23_,
  r_n_61__22_,r_n_61__21_,r_n_61__20_,r_n_61__19_,r_n_61__18_,r_n_61__17_,r_n_61__16_,
  r_n_61__15_,r_n_61__14_,r_n_61__13_,r_n_61__12_,r_n_61__11_,r_n_61__10_,
  r_n_61__9_,r_n_61__8_,r_n_61__7_,r_n_61__6_,r_n_61__5_,r_n_61__4_,r_n_61__3_,r_n_61__2_,
  r_n_61__1_,r_n_61__0_,r_n_60__63_,r_n_60__62_,r_n_60__61_,r_n_60__60_,
  r_n_60__59_,r_n_60__58_,r_n_60__57_,r_n_60__56_,r_n_60__55_,r_n_60__54_,r_n_60__53_,
  r_n_60__52_,r_n_60__51_,r_n_60__50_,r_n_60__49_,r_n_60__48_,r_n_60__47_,r_n_60__46_,
  r_n_60__45_,r_n_60__44_,r_n_60__43_,r_n_60__42_,r_n_60__41_,r_n_60__40_,
  r_n_60__39_,r_n_60__38_,r_n_60__37_,r_n_60__36_,r_n_60__35_,r_n_60__34_,r_n_60__33_,
  r_n_60__32_,r_n_60__31_,r_n_60__30_,r_n_60__29_,r_n_60__28_,r_n_60__27_,r_n_60__26_,
  r_n_60__25_,r_n_60__24_,r_n_60__23_,r_n_60__22_,r_n_60__21_,r_n_60__20_,
  r_n_60__19_,r_n_60__18_,r_n_60__17_,r_n_60__16_,r_n_60__15_,r_n_60__14_,r_n_60__13_,
  r_n_60__12_,r_n_60__11_,r_n_60__10_,r_n_60__9_,r_n_60__8_,r_n_60__7_,r_n_60__6_,
  r_n_60__5_,r_n_60__4_,r_n_60__3_,r_n_60__2_,r_n_60__1_,r_n_60__0_,r_n_59__63_,
  r_n_59__62_,r_n_59__61_,r_n_59__60_,r_n_59__59_,r_n_59__58_,r_n_59__57_,r_n_59__56_,
  r_n_59__55_,r_n_59__54_,r_n_59__53_,r_n_59__52_,r_n_59__51_,r_n_59__50_,r_n_59__49_,
  r_n_59__48_,r_n_59__47_,r_n_59__46_,r_n_59__45_,r_n_59__44_,r_n_59__43_,
  r_n_59__42_,r_n_59__41_,r_n_59__40_,r_n_59__39_,r_n_59__38_,r_n_59__37_,r_n_59__36_,
  r_n_59__35_,r_n_59__34_,r_n_59__33_,r_n_59__32_,r_n_59__31_,r_n_59__30_,r_n_59__29_,
  r_n_59__28_,r_n_59__27_,r_n_59__26_,r_n_59__25_,r_n_59__24_,r_n_59__23_,
  r_n_59__22_,r_n_59__21_,r_n_59__20_,r_n_59__19_,r_n_59__18_,r_n_59__17_,r_n_59__16_,
  r_n_59__15_,r_n_59__14_,r_n_59__13_,r_n_59__12_,r_n_59__11_,r_n_59__10_,r_n_59__9_,
  r_n_59__8_,r_n_59__7_,r_n_59__6_,r_n_59__5_,r_n_59__4_,r_n_59__3_,r_n_59__2_,
  r_n_59__1_,r_n_59__0_,r_n_58__63_,r_n_58__62_,r_n_58__61_,r_n_58__60_,r_n_58__59_,
  r_n_58__58_,r_n_58__57_,r_n_58__56_,r_n_58__55_,r_n_58__54_,r_n_58__53_,
  r_n_58__52_,r_n_58__51_,r_n_58__50_,r_n_58__49_,r_n_58__48_,r_n_58__47_,r_n_58__46_,
  r_n_58__45_,r_n_58__44_,r_n_58__43_,r_n_58__42_,r_n_58__41_,r_n_58__40_,r_n_58__39_,
  r_n_58__38_,r_n_58__37_,r_n_58__36_,r_n_58__35_,r_n_58__34_,r_n_58__33_,
  r_n_58__32_,r_n_58__31_,r_n_58__30_,r_n_58__29_,r_n_58__28_,r_n_58__27_,r_n_58__26_,
  r_n_58__25_,r_n_58__24_,r_n_58__23_,r_n_58__22_,r_n_58__21_,r_n_58__20_,r_n_58__19_,
  r_n_58__18_,r_n_58__17_,r_n_58__16_,r_n_58__15_,r_n_58__14_,r_n_58__13_,
  r_n_58__12_,r_n_58__11_,r_n_58__10_,r_n_58__9_,r_n_58__8_,r_n_58__7_,r_n_58__6_,
  r_n_58__5_,r_n_58__4_,r_n_58__3_,r_n_58__2_,r_n_58__1_,r_n_58__0_,r_n_57__63_,r_n_57__62_,
  r_n_57__61_,r_n_57__60_,r_n_57__59_,r_n_57__58_,r_n_57__57_,r_n_57__56_,
  r_n_57__55_,r_n_57__54_,r_n_57__53_,r_n_57__52_,r_n_57__51_,r_n_57__50_,r_n_57__49_,
  r_n_57__48_,r_n_57__47_,r_n_57__46_,r_n_57__45_,r_n_57__44_,r_n_57__43_,r_n_57__42_,
  r_n_57__41_,r_n_57__40_,r_n_57__39_,r_n_57__38_,r_n_57__37_,r_n_57__36_,
  r_n_57__35_,r_n_57__34_,r_n_57__33_,r_n_57__32_,r_n_57__31_,r_n_57__30_,r_n_57__29_,
  r_n_57__28_,r_n_57__27_,r_n_57__26_,r_n_57__25_,r_n_57__24_,r_n_57__23_,r_n_57__22_,
  r_n_57__21_,r_n_57__20_,r_n_57__19_,r_n_57__18_,r_n_57__17_,r_n_57__16_,
  r_n_57__15_,r_n_57__14_,r_n_57__13_,r_n_57__12_,r_n_57__11_,r_n_57__10_,r_n_57__9_,
  r_n_57__8_,r_n_57__7_,r_n_57__6_,r_n_57__5_,r_n_57__4_,r_n_57__3_,r_n_57__2_,
  r_n_57__1_,r_n_57__0_,r_n_72__63_,r_n_72__62_,r_n_72__61_,r_n_72__60_,r_n_72__59_,
  r_n_72__58_,r_n_72__57_,r_n_72__56_,r_n_72__55_,r_n_72__54_,r_n_72__53_,r_n_72__52_,
  r_n_72__51_,r_n_72__50_,r_n_72__49_,r_n_72__48_,r_n_72__47_,r_n_72__46_,
  r_n_72__45_,r_n_72__44_,r_n_72__43_,r_n_72__42_,r_n_72__41_,r_n_72__40_,r_n_72__39_,
  r_n_72__38_,r_n_72__37_,r_n_72__36_,r_n_72__35_,r_n_72__34_,r_n_72__33_,r_n_72__32_,
  r_n_72__31_,r_n_72__30_,r_n_72__29_,r_n_72__28_,r_n_72__27_,r_n_72__26_,
  r_n_72__25_,r_n_72__24_,r_n_72__23_,r_n_72__22_,r_n_72__21_,r_n_72__20_,r_n_72__19_,
  r_n_72__18_,r_n_72__17_,r_n_72__16_,r_n_72__15_,r_n_72__14_,r_n_72__13_,r_n_72__12_,
  r_n_72__11_,r_n_72__10_,r_n_72__9_,r_n_72__8_,r_n_72__7_,r_n_72__6_,r_n_72__5_,
  r_n_72__4_,r_n_72__3_,r_n_72__2_,r_n_72__1_,r_n_72__0_,r_n_71__63_,r_n_71__62_,
  r_n_71__61_,r_n_71__60_,r_n_71__59_,r_n_71__58_,r_n_71__57_,r_n_71__56_,r_n_71__55_,
  r_n_71__54_,r_n_71__53_,r_n_71__52_,r_n_71__51_,r_n_71__50_,r_n_71__49_,
  r_n_71__48_,r_n_71__47_,r_n_71__46_,r_n_71__45_,r_n_71__44_,r_n_71__43_,r_n_71__42_,
  r_n_71__41_,r_n_71__40_,r_n_71__39_,r_n_71__38_,r_n_71__37_,r_n_71__36_,r_n_71__35_,
  r_n_71__34_,r_n_71__33_,r_n_71__32_,r_n_71__31_,r_n_71__30_,r_n_71__29_,
  r_n_71__28_,r_n_71__27_,r_n_71__26_,r_n_71__25_,r_n_71__24_,r_n_71__23_,r_n_71__22_,
  r_n_71__21_,r_n_71__20_,r_n_71__19_,r_n_71__18_,r_n_71__17_,r_n_71__16_,r_n_71__15_,
  r_n_71__14_,r_n_71__13_,r_n_71__12_,r_n_71__11_,r_n_71__10_,r_n_71__9_,
  r_n_71__8_,r_n_71__7_,r_n_71__6_,r_n_71__5_,r_n_71__4_,r_n_71__3_,r_n_71__2_,r_n_71__1_,
  r_n_71__0_,r_n_70__63_,r_n_70__62_,r_n_70__61_,r_n_70__60_,r_n_70__59_,
  r_n_70__58_,r_n_70__57_,r_n_70__56_,r_n_70__55_,r_n_70__54_,r_n_70__53_,r_n_70__52_,
  r_n_70__51_,r_n_70__50_,r_n_70__49_,r_n_70__48_,r_n_70__47_,r_n_70__46_,r_n_70__45_,
  r_n_70__44_,r_n_70__43_,r_n_70__42_,r_n_70__41_,r_n_70__40_,r_n_70__39_,
  r_n_70__38_,r_n_70__37_,r_n_70__36_,r_n_70__35_,r_n_70__34_,r_n_70__33_,r_n_70__32_,
  r_n_70__31_,r_n_70__30_,r_n_70__29_,r_n_70__28_,r_n_70__27_,r_n_70__26_,r_n_70__25_,
  r_n_70__24_,r_n_70__23_,r_n_70__22_,r_n_70__21_,r_n_70__20_,r_n_70__19_,
  r_n_70__18_,r_n_70__17_,r_n_70__16_,r_n_70__15_,r_n_70__14_,r_n_70__13_,r_n_70__12_,
  r_n_70__11_,r_n_70__10_,r_n_70__9_,r_n_70__8_,r_n_70__7_,r_n_70__6_,r_n_70__5_,
  r_n_70__4_,r_n_70__3_,r_n_70__2_,r_n_70__1_,r_n_70__0_,r_n_69__63_,r_n_69__62_,
  r_n_69__61_,r_n_69__60_,r_n_69__59_,r_n_69__58_,r_n_69__57_,r_n_69__56_,r_n_69__55_,
  r_n_69__54_,r_n_69__53_,r_n_69__52_,r_n_69__51_,r_n_69__50_,r_n_69__49_,r_n_69__48_,
  r_n_69__47_,r_n_69__46_,r_n_69__45_,r_n_69__44_,r_n_69__43_,r_n_69__42_,
  r_n_69__41_,r_n_69__40_,r_n_69__39_,r_n_69__38_,r_n_69__37_,r_n_69__36_,r_n_69__35_,
  r_n_69__34_,r_n_69__33_,r_n_69__32_,r_n_69__31_,r_n_69__30_,r_n_69__29_,r_n_69__28_,
  r_n_69__27_,r_n_69__26_,r_n_69__25_,r_n_69__24_,r_n_69__23_,r_n_69__22_,
  r_n_69__21_,r_n_69__20_,r_n_69__19_,r_n_69__18_,r_n_69__17_,r_n_69__16_,r_n_69__15_,
  r_n_69__14_,r_n_69__13_,r_n_69__12_,r_n_69__11_,r_n_69__10_,r_n_69__9_,r_n_69__8_,
  r_n_69__7_,r_n_69__6_,r_n_69__5_,r_n_69__4_,r_n_69__3_,r_n_69__2_,r_n_69__1_,
  r_n_69__0_,r_n_68__63_,r_n_68__62_,r_n_68__61_,r_n_68__60_,r_n_68__59_,r_n_68__58_,
  r_n_68__57_,r_n_68__56_,r_n_68__55_,r_n_68__54_,r_n_68__53_,r_n_68__52_,
  r_n_68__51_,r_n_68__50_,r_n_68__49_,r_n_68__48_,r_n_68__47_,r_n_68__46_,r_n_68__45_,
  r_n_68__44_,r_n_68__43_,r_n_68__42_,r_n_68__41_,r_n_68__40_,r_n_68__39_,r_n_68__38_,
  r_n_68__37_,r_n_68__36_,r_n_68__35_,r_n_68__34_,r_n_68__33_,r_n_68__32_,
  r_n_68__31_,r_n_68__30_,r_n_68__29_,r_n_68__28_,r_n_68__27_,r_n_68__26_,r_n_68__25_,
  r_n_68__24_,r_n_68__23_,r_n_68__22_,r_n_68__21_,r_n_68__20_,r_n_68__19_,r_n_68__18_,
  r_n_68__17_,r_n_68__16_,r_n_68__15_,r_n_68__14_,r_n_68__13_,r_n_68__12_,
  r_n_68__11_,r_n_68__10_,r_n_68__9_,r_n_68__8_,r_n_68__7_,r_n_68__6_,r_n_68__5_,r_n_68__4_,
  r_n_68__3_,r_n_68__2_,r_n_68__1_,r_n_68__0_,r_n_67__63_,r_n_67__62_,r_n_67__61_,
  r_n_67__60_,r_n_67__59_,r_n_67__58_,r_n_67__57_,r_n_67__56_,r_n_67__55_,
  r_n_67__54_,r_n_67__53_,r_n_67__52_,r_n_67__51_,r_n_67__50_,r_n_67__49_,r_n_67__48_,
  r_n_67__47_,r_n_67__46_,r_n_67__45_,r_n_67__44_,r_n_67__43_,r_n_67__42_,r_n_67__41_,
  r_n_67__40_,r_n_67__39_,r_n_67__38_,r_n_67__37_,r_n_67__36_,r_n_67__35_,
  r_n_67__34_,r_n_67__33_,r_n_67__32_,r_n_67__31_,r_n_67__30_,r_n_67__29_,r_n_67__28_,
  r_n_67__27_,r_n_67__26_,r_n_67__25_,r_n_67__24_,r_n_67__23_,r_n_67__22_,r_n_67__21_,
  r_n_67__20_,r_n_67__19_,r_n_67__18_,r_n_67__17_,r_n_67__16_,r_n_67__15_,
  r_n_67__14_,r_n_67__13_,r_n_67__12_,r_n_67__11_,r_n_67__10_,r_n_67__9_,r_n_67__8_,
  r_n_67__7_,r_n_67__6_,r_n_67__5_,r_n_67__4_,r_n_67__3_,r_n_67__2_,r_n_67__1_,
  r_n_67__0_,r_n_66__63_,r_n_66__62_,r_n_66__61_,r_n_66__60_,r_n_66__59_,r_n_66__58_,
  r_n_66__57_,r_n_66__56_,r_n_66__55_,r_n_66__54_,r_n_66__53_,r_n_66__52_,r_n_66__51_,
  r_n_66__50_,r_n_66__49_,r_n_66__48_,r_n_66__47_,r_n_66__46_,r_n_66__45_,
  r_n_66__44_,r_n_66__43_,r_n_66__42_,r_n_66__41_,r_n_66__40_,r_n_66__39_,r_n_66__38_,
  r_n_66__37_,r_n_66__36_,r_n_66__35_,r_n_66__34_,r_n_66__33_,r_n_66__32_,r_n_66__31_,
  r_n_66__30_,r_n_66__29_,r_n_66__28_,r_n_66__27_,r_n_66__26_,r_n_66__25_,
  r_n_66__24_,r_n_66__23_,r_n_66__22_,r_n_66__21_,r_n_66__20_,r_n_66__19_,r_n_66__18_,
  r_n_66__17_,r_n_66__16_,r_n_66__15_,r_n_66__14_,r_n_66__13_,r_n_66__12_,r_n_66__11_,
  r_n_66__10_,r_n_66__9_,r_n_66__8_,r_n_66__7_,r_n_66__6_,r_n_66__5_,r_n_66__4_,
  r_n_66__3_,r_n_66__2_,r_n_66__1_,r_n_66__0_,r_n_65__63_,r_n_65__62_,r_n_65__61_,
  r_n_65__60_,r_n_65__59_,r_n_65__58_,r_n_65__57_,r_n_65__56_,r_n_65__55_,r_n_65__54_,
  r_n_65__53_,r_n_65__52_,r_n_65__51_,r_n_65__50_,r_n_65__49_,r_n_65__48_,
  r_n_65__47_,r_n_65__46_,r_n_65__45_,r_n_65__44_,r_n_65__43_,r_n_65__42_,r_n_65__41_,
  r_n_65__40_,r_n_65__39_,r_n_65__38_,r_n_65__37_,r_n_65__36_,r_n_65__35_,r_n_65__34_,
  r_n_65__33_,r_n_65__32_,r_n_65__31_,r_n_65__30_,r_n_65__29_,r_n_65__28_,
  r_n_65__27_,r_n_65__26_,r_n_65__25_,r_n_65__24_,r_n_65__23_,r_n_65__22_,r_n_65__21_,
  r_n_65__20_,r_n_65__19_,r_n_65__18_,r_n_65__17_,r_n_65__16_,r_n_65__15_,r_n_65__14_,
  r_n_65__13_,r_n_65__12_,r_n_65__11_,r_n_65__10_,r_n_65__9_,r_n_65__8_,
  r_n_65__7_,r_n_65__6_,r_n_65__5_,r_n_65__4_,r_n_65__3_,r_n_65__2_,r_n_65__1_,r_n_65__0_,
  r_n_80__63_,r_n_80__62_,r_n_80__61_,r_n_80__60_,r_n_80__59_,r_n_80__58_,
  r_n_80__57_,r_n_80__56_,r_n_80__55_,r_n_80__54_,r_n_80__53_,r_n_80__52_,r_n_80__51_,
  r_n_80__50_,r_n_80__49_,r_n_80__48_,r_n_80__47_,r_n_80__46_,r_n_80__45_,r_n_80__44_,
  r_n_80__43_,r_n_80__42_,r_n_80__41_,r_n_80__40_,r_n_80__39_,r_n_80__38_,
  r_n_80__37_,r_n_80__36_,r_n_80__35_,r_n_80__34_,r_n_80__33_,r_n_80__32_,r_n_80__31_,
  r_n_80__30_,r_n_80__29_,r_n_80__28_,r_n_80__27_,r_n_80__26_,r_n_80__25_,r_n_80__24_,
  r_n_80__23_,r_n_80__22_,r_n_80__21_,r_n_80__20_,r_n_80__19_,r_n_80__18_,
  r_n_80__17_,r_n_80__16_,r_n_80__15_,r_n_80__14_,r_n_80__13_,r_n_80__12_,r_n_80__11_,
  r_n_80__10_,r_n_80__9_,r_n_80__8_,r_n_80__7_,r_n_80__6_,r_n_80__5_,r_n_80__4_,
  r_n_80__3_,r_n_80__2_,r_n_80__1_,r_n_80__0_,r_n_79__63_,r_n_79__62_,r_n_79__61_,
  r_n_79__60_,r_n_79__59_,r_n_79__58_,r_n_79__57_,r_n_79__56_,r_n_79__55_,r_n_79__54_,
  r_n_79__53_,r_n_79__52_,r_n_79__51_,r_n_79__50_,r_n_79__49_,r_n_79__48_,r_n_79__47_,
  r_n_79__46_,r_n_79__45_,r_n_79__44_,r_n_79__43_,r_n_79__42_,r_n_79__41_,
  r_n_79__40_,r_n_79__39_,r_n_79__38_,r_n_79__37_,r_n_79__36_,r_n_79__35_,r_n_79__34_,
  r_n_79__33_,r_n_79__32_,r_n_79__31_,r_n_79__30_,r_n_79__29_,r_n_79__28_,r_n_79__27_,
  r_n_79__26_,r_n_79__25_,r_n_79__24_,r_n_79__23_,r_n_79__22_,r_n_79__21_,
  r_n_79__20_,r_n_79__19_,r_n_79__18_,r_n_79__17_,r_n_79__16_,r_n_79__15_,r_n_79__14_,
  r_n_79__13_,r_n_79__12_,r_n_79__11_,r_n_79__10_,r_n_79__9_,r_n_79__8_,r_n_79__7_,
  r_n_79__6_,r_n_79__5_,r_n_79__4_,r_n_79__3_,r_n_79__2_,r_n_79__1_,r_n_79__0_,
  r_n_78__63_,r_n_78__62_,r_n_78__61_,r_n_78__60_,r_n_78__59_,r_n_78__58_,r_n_78__57_,
  r_n_78__56_,r_n_78__55_,r_n_78__54_,r_n_78__53_,r_n_78__52_,r_n_78__51_,
  r_n_78__50_,r_n_78__49_,r_n_78__48_,r_n_78__47_,r_n_78__46_,r_n_78__45_,r_n_78__44_,
  r_n_78__43_,r_n_78__42_,r_n_78__41_,r_n_78__40_,r_n_78__39_,r_n_78__38_,r_n_78__37_,
  r_n_78__36_,r_n_78__35_,r_n_78__34_,r_n_78__33_,r_n_78__32_,r_n_78__31_,
  r_n_78__30_,r_n_78__29_,r_n_78__28_,r_n_78__27_,r_n_78__26_,r_n_78__25_,r_n_78__24_,
  r_n_78__23_,r_n_78__22_,r_n_78__21_,r_n_78__20_,r_n_78__19_,r_n_78__18_,r_n_78__17_,
  r_n_78__16_,r_n_78__15_,r_n_78__14_,r_n_78__13_,r_n_78__12_,r_n_78__11_,
  r_n_78__10_,r_n_78__9_,r_n_78__8_,r_n_78__7_,r_n_78__6_,r_n_78__5_,r_n_78__4_,r_n_78__3_,
  r_n_78__2_,r_n_78__1_,r_n_78__0_,r_n_77__63_,r_n_77__62_,r_n_77__61_,r_n_77__60_,
  r_n_77__59_,r_n_77__58_,r_n_77__57_,r_n_77__56_,r_n_77__55_,r_n_77__54_,
  r_n_77__53_,r_n_77__52_,r_n_77__51_,r_n_77__50_,r_n_77__49_,r_n_77__48_,r_n_77__47_,
  r_n_77__46_,r_n_77__45_,r_n_77__44_,r_n_77__43_,r_n_77__42_,r_n_77__41_,r_n_77__40_,
  r_n_77__39_,r_n_77__38_,r_n_77__37_,r_n_77__36_,r_n_77__35_,r_n_77__34_,
  r_n_77__33_,r_n_77__32_,r_n_77__31_,r_n_77__30_,r_n_77__29_,r_n_77__28_,r_n_77__27_,
  r_n_77__26_,r_n_77__25_,r_n_77__24_,r_n_77__23_,r_n_77__22_,r_n_77__21_,r_n_77__20_,
  r_n_77__19_,r_n_77__18_,r_n_77__17_,r_n_77__16_,r_n_77__15_,r_n_77__14_,
  r_n_77__13_,r_n_77__12_,r_n_77__11_,r_n_77__10_,r_n_77__9_,r_n_77__8_,r_n_77__7_,
  r_n_77__6_,r_n_77__5_,r_n_77__4_,r_n_77__3_,r_n_77__2_,r_n_77__1_,r_n_77__0_,
  r_n_76__63_,r_n_76__62_,r_n_76__61_,r_n_76__60_,r_n_76__59_,r_n_76__58_,r_n_76__57_,
  r_n_76__56_,r_n_76__55_,r_n_76__54_,r_n_76__53_,r_n_76__52_,r_n_76__51_,r_n_76__50_,
  r_n_76__49_,r_n_76__48_,r_n_76__47_,r_n_76__46_,r_n_76__45_,r_n_76__44_,
  r_n_76__43_,r_n_76__42_,r_n_76__41_,r_n_76__40_,r_n_76__39_,r_n_76__38_,r_n_76__37_,
  r_n_76__36_,r_n_76__35_,r_n_76__34_,r_n_76__33_,r_n_76__32_,r_n_76__31_,r_n_76__30_,
  r_n_76__29_,r_n_76__28_,r_n_76__27_,r_n_76__26_,r_n_76__25_,r_n_76__24_,
  r_n_76__23_,r_n_76__22_,r_n_76__21_,r_n_76__20_,r_n_76__19_,r_n_76__18_,r_n_76__17_,
  r_n_76__16_,r_n_76__15_,r_n_76__14_,r_n_76__13_,r_n_76__12_,r_n_76__11_,r_n_76__10_,
  r_n_76__9_,r_n_76__8_,r_n_76__7_,r_n_76__6_,r_n_76__5_,r_n_76__4_,r_n_76__3_,
  r_n_76__2_,r_n_76__1_,r_n_76__0_,r_n_75__63_,r_n_75__62_,r_n_75__61_,r_n_75__60_,
  r_n_75__59_,r_n_75__58_,r_n_75__57_,r_n_75__56_,r_n_75__55_,r_n_75__54_,r_n_75__53_,
  r_n_75__52_,r_n_75__51_,r_n_75__50_,r_n_75__49_,r_n_75__48_,r_n_75__47_,
  r_n_75__46_,r_n_75__45_,r_n_75__44_,r_n_75__43_,r_n_75__42_,r_n_75__41_,r_n_75__40_,
  r_n_75__39_,r_n_75__38_,r_n_75__37_,r_n_75__36_,r_n_75__35_,r_n_75__34_,r_n_75__33_,
  r_n_75__32_,r_n_75__31_,r_n_75__30_,r_n_75__29_,r_n_75__28_,r_n_75__27_,
  r_n_75__26_,r_n_75__25_,r_n_75__24_,r_n_75__23_,r_n_75__22_,r_n_75__21_,r_n_75__20_,
  r_n_75__19_,r_n_75__18_,r_n_75__17_,r_n_75__16_,r_n_75__15_,r_n_75__14_,r_n_75__13_,
  r_n_75__12_,r_n_75__11_,r_n_75__10_,r_n_75__9_,r_n_75__8_,r_n_75__7_,r_n_75__6_,
  r_n_75__5_,r_n_75__4_,r_n_75__3_,r_n_75__2_,r_n_75__1_,r_n_75__0_,r_n_74__63_,
  r_n_74__62_,r_n_74__61_,r_n_74__60_,r_n_74__59_,r_n_74__58_,r_n_74__57_,
  r_n_74__56_,r_n_74__55_,r_n_74__54_,r_n_74__53_,r_n_74__52_,r_n_74__51_,r_n_74__50_,
  r_n_74__49_,r_n_74__48_,r_n_74__47_,r_n_74__46_,r_n_74__45_,r_n_74__44_,r_n_74__43_,
  r_n_74__42_,r_n_74__41_,r_n_74__40_,r_n_74__39_,r_n_74__38_,r_n_74__37_,
  r_n_74__36_,r_n_74__35_,r_n_74__34_,r_n_74__33_,r_n_74__32_,r_n_74__31_,r_n_74__30_,
  r_n_74__29_,r_n_74__28_,r_n_74__27_,r_n_74__26_,r_n_74__25_,r_n_74__24_,r_n_74__23_,
  r_n_74__22_,r_n_74__21_,r_n_74__20_,r_n_74__19_,r_n_74__18_,r_n_74__17_,
  r_n_74__16_,r_n_74__15_,r_n_74__14_,r_n_74__13_,r_n_74__12_,r_n_74__11_,r_n_74__10_,
  r_n_74__9_,r_n_74__8_,r_n_74__7_,r_n_74__6_,r_n_74__5_,r_n_74__4_,r_n_74__3_,
  r_n_74__2_,r_n_74__1_,r_n_74__0_,r_n_73__63_,r_n_73__62_,r_n_73__61_,r_n_73__60_,
  r_n_73__59_,r_n_73__58_,r_n_73__57_,r_n_73__56_,r_n_73__55_,r_n_73__54_,r_n_73__53_,
  r_n_73__52_,r_n_73__51_,r_n_73__50_,r_n_73__49_,r_n_73__48_,r_n_73__47_,r_n_73__46_,
  r_n_73__45_,r_n_73__44_,r_n_73__43_,r_n_73__42_,r_n_73__41_,r_n_73__40_,
  r_n_73__39_,r_n_73__38_,r_n_73__37_,r_n_73__36_,r_n_73__35_,r_n_73__34_,r_n_73__33_,
  r_n_73__32_,r_n_73__31_,r_n_73__30_,r_n_73__29_,r_n_73__28_,r_n_73__27_,r_n_73__26_,
  r_n_73__25_,r_n_73__24_,r_n_73__23_,r_n_73__22_,r_n_73__21_,r_n_73__20_,
  r_n_73__19_,r_n_73__18_,r_n_73__17_,r_n_73__16_,r_n_73__15_,r_n_73__14_,r_n_73__13_,
  r_n_73__12_,r_n_73__11_,r_n_73__10_,r_n_73__9_,r_n_73__8_,r_n_73__7_,r_n_73__6_,
  r_n_73__5_,r_n_73__4_,r_n_73__3_,r_n_73__2_,r_n_73__1_,r_n_73__0_,r_n_88__63_,
  r_n_88__62_,r_n_88__61_,r_n_88__60_,r_n_88__59_,r_n_88__58_,r_n_88__57_,r_n_88__56_,
  r_n_88__55_,r_n_88__54_,r_n_88__53_,r_n_88__52_,r_n_88__51_,r_n_88__50_,
  r_n_88__49_,r_n_88__48_,r_n_88__47_,r_n_88__46_,r_n_88__45_,r_n_88__44_,r_n_88__43_,
  r_n_88__42_,r_n_88__41_,r_n_88__40_,r_n_88__39_,r_n_88__38_,r_n_88__37_,r_n_88__36_,
  r_n_88__35_,r_n_88__34_,r_n_88__33_,r_n_88__32_,r_n_88__31_,r_n_88__30_,
  r_n_88__29_,r_n_88__28_,r_n_88__27_,r_n_88__26_,r_n_88__25_,r_n_88__24_,r_n_88__23_,
  r_n_88__22_,r_n_88__21_,r_n_88__20_,r_n_88__19_,r_n_88__18_,r_n_88__17_,r_n_88__16_,
  r_n_88__15_,r_n_88__14_,r_n_88__13_,r_n_88__12_,r_n_88__11_,r_n_88__10_,
  r_n_88__9_,r_n_88__8_,r_n_88__7_,r_n_88__6_,r_n_88__5_,r_n_88__4_,r_n_88__3_,r_n_88__2_,
  r_n_88__1_,r_n_88__0_,r_n_87__63_,r_n_87__62_,r_n_87__61_,r_n_87__60_,r_n_87__59_,
  r_n_87__58_,r_n_87__57_,r_n_87__56_,r_n_87__55_,r_n_87__54_,r_n_87__53_,
  r_n_87__52_,r_n_87__51_,r_n_87__50_,r_n_87__49_,r_n_87__48_,r_n_87__47_,r_n_87__46_,
  r_n_87__45_,r_n_87__44_,r_n_87__43_,r_n_87__42_,r_n_87__41_,r_n_87__40_,r_n_87__39_,
  r_n_87__38_,r_n_87__37_,r_n_87__36_,r_n_87__35_,r_n_87__34_,r_n_87__33_,
  r_n_87__32_,r_n_87__31_,r_n_87__30_,r_n_87__29_,r_n_87__28_,r_n_87__27_,r_n_87__26_,
  r_n_87__25_,r_n_87__24_,r_n_87__23_,r_n_87__22_,r_n_87__21_,r_n_87__20_,r_n_87__19_,
  r_n_87__18_,r_n_87__17_,r_n_87__16_,r_n_87__15_,r_n_87__14_,r_n_87__13_,
  r_n_87__12_,r_n_87__11_,r_n_87__10_,r_n_87__9_,r_n_87__8_,r_n_87__7_,r_n_87__6_,
  r_n_87__5_,r_n_87__4_,r_n_87__3_,r_n_87__2_,r_n_87__1_,r_n_87__0_,r_n_86__63_,
  r_n_86__62_,r_n_86__61_,r_n_86__60_,r_n_86__59_,r_n_86__58_,r_n_86__57_,r_n_86__56_,
  r_n_86__55_,r_n_86__54_,r_n_86__53_,r_n_86__52_,r_n_86__51_,r_n_86__50_,r_n_86__49_,
  r_n_86__48_,r_n_86__47_,r_n_86__46_,r_n_86__45_,r_n_86__44_,r_n_86__43_,
  r_n_86__42_,r_n_86__41_,r_n_86__40_,r_n_86__39_,r_n_86__38_,r_n_86__37_,r_n_86__36_,
  r_n_86__35_,r_n_86__34_,r_n_86__33_,r_n_86__32_,r_n_86__31_,r_n_86__30_,r_n_86__29_,
  r_n_86__28_,r_n_86__27_,r_n_86__26_,r_n_86__25_,r_n_86__24_,r_n_86__23_,
  r_n_86__22_,r_n_86__21_,r_n_86__20_,r_n_86__19_,r_n_86__18_,r_n_86__17_,r_n_86__16_,
  r_n_86__15_,r_n_86__14_,r_n_86__13_,r_n_86__12_,r_n_86__11_,r_n_86__10_,r_n_86__9_,
  r_n_86__8_,r_n_86__7_,r_n_86__6_,r_n_86__5_,r_n_86__4_,r_n_86__3_,r_n_86__2_,
  r_n_86__1_,r_n_86__0_,r_n_85__63_,r_n_85__62_,r_n_85__61_,r_n_85__60_,r_n_85__59_,
  r_n_85__58_,r_n_85__57_,r_n_85__56_,r_n_85__55_,r_n_85__54_,r_n_85__53_,r_n_85__52_,
  r_n_85__51_,r_n_85__50_,r_n_85__49_,r_n_85__48_,r_n_85__47_,r_n_85__46_,
  r_n_85__45_,r_n_85__44_,r_n_85__43_,r_n_85__42_,r_n_85__41_,r_n_85__40_,r_n_85__39_,
  r_n_85__38_,r_n_85__37_,r_n_85__36_,r_n_85__35_,r_n_85__34_,r_n_85__33_,r_n_85__32_,
  r_n_85__31_,r_n_85__30_,r_n_85__29_,r_n_85__28_,r_n_85__27_,r_n_85__26_,
  r_n_85__25_,r_n_85__24_,r_n_85__23_,r_n_85__22_,r_n_85__21_,r_n_85__20_,r_n_85__19_,
  r_n_85__18_,r_n_85__17_,r_n_85__16_,r_n_85__15_,r_n_85__14_,r_n_85__13_,r_n_85__12_,
  r_n_85__11_,r_n_85__10_,r_n_85__9_,r_n_85__8_,r_n_85__7_,r_n_85__6_,r_n_85__5_,
  r_n_85__4_,r_n_85__3_,r_n_85__2_,r_n_85__1_,r_n_85__0_,r_n_84__63_,r_n_84__62_,
  r_n_84__61_,r_n_84__60_,r_n_84__59_,r_n_84__58_,r_n_84__57_,r_n_84__56_,
  r_n_84__55_,r_n_84__54_,r_n_84__53_,r_n_84__52_,r_n_84__51_,r_n_84__50_,r_n_84__49_,
  r_n_84__48_,r_n_84__47_,r_n_84__46_,r_n_84__45_,r_n_84__44_,r_n_84__43_,r_n_84__42_,
  r_n_84__41_,r_n_84__40_,r_n_84__39_,r_n_84__38_,r_n_84__37_,r_n_84__36_,
  r_n_84__35_,r_n_84__34_,r_n_84__33_,r_n_84__32_,r_n_84__31_,r_n_84__30_,r_n_84__29_,
  r_n_84__28_,r_n_84__27_,r_n_84__26_,r_n_84__25_,r_n_84__24_,r_n_84__23_,r_n_84__22_,
  r_n_84__21_,r_n_84__20_,r_n_84__19_,r_n_84__18_,r_n_84__17_,r_n_84__16_,
  r_n_84__15_,r_n_84__14_,r_n_84__13_,r_n_84__12_,r_n_84__11_,r_n_84__10_,r_n_84__9_,
  r_n_84__8_,r_n_84__7_,r_n_84__6_,r_n_84__5_,r_n_84__4_,r_n_84__3_,r_n_84__2_,
  r_n_84__1_,r_n_84__0_,r_n_83__63_,r_n_83__62_,r_n_83__61_,r_n_83__60_,r_n_83__59_,
  r_n_83__58_,r_n_83__57_,r_n_83__56_,r_n_83__55_,r_n_83__54_,r_n_83__53_,r_n_83__52_,
  r_n_83__51_,r_n_83__50_,r_n_83__49_,r_n_83__48_,r_n_83__47_,r_n_83__46_,r_n_83__45_,
  r_n_83__44_,r_n_83__43_,r_n_83__42_,r_n_83__41_,r_n_83__40_,r_n_83__39_,
  r_n_83__38_,r_n_83__37_,r_n_83__36_,r_n_83__35_,r_n_83__34_,r_n_83__33_,r_n_83__32_,
  r_n_83__31_,r_n_83__30_,r_n_83__29_,r_n_83__28_,r_n_83__27_,r_n_83__26_,r_n_83__25_,
  r_n_83__24_,r_n_83__23_,r_n_83__22_,r_n_83__21_,r_n_83__20_,r_n_83__19_,
  r_n_83__18_,r_n_83__17_,r_n_83__16_,r_n_83__15_,r_n_83__14_,r_n_83__13_,r_n_83__12_,
  r_n_83__11_,r_n_83__10_,r_n_83__9_,r_n_83__8_,r_n_83__7_,r_n_83__6_,r_n_83__5_,
  r_n_83__4_,r_n_83__3_,r_n_83__2_,r_n_83__1_,r_n_83__0_,r_n_82__63_,r_n_82__62_,
  r_n_82__61_,r_n_82__60_,r_n_82__59_,r_n_82__58_,r_n_82__57_,r_n_82__56_,r_n_82__55_,
  r_n_82__54_,r_n_82__53_,r_n_82__52_,r_n_82__51_,r_n_82__50_,r_n_82__49_,
  r_n_82__48_,r_n_82__47_,r_n_82__46_,r_n_82__45_,r_n_82__44_,r_n_82__43_,r_n_82__42_,
  r_n_82__41_,r_n_82__40_,r_n_82__39_,r_n_82__38_,r_n_82__37_,r_n_82__36_,r_n_82__35_,
  r_n_82__34_,r_n_82__33_,r_n_82__32_,r_n_82__31_,r_n_82__30_,r_n_82__29_,
  r_n_82__28_,r_n_82__27_,r_n_82__26_,r_n_82__25_,r_n_82__24_,r_n_82__23_,r_n_82__22_,
  r_n_82__21_,r_n_82__20_,r_n_82__19_,r_n_82__18_,r_n_82__17_,r_n_82__16_,r_n_82__15_,
  r_n_82__14_,r_n_82__13_,r_n_82__12_,r_n_82__11_,r_n_82__10_,r_n_82__9_,r_n_82__8_,
  r_n_82__7_,r_n_82__6_,r_n_82__5_,r_n_82__4_,r_n_82__3_,r_n_82__2_,r_n_82__1_,
  r_n_82__0_,r_n_81__63_,r_n_81__62_,r_n_81__61_,r_n_81__60_,r_n_81__59_,r_n_81__58_,
  r_n_81__57_,r_n_81__56_,r_n_81__55_,r_n_81__54_,r_n_81__53_,r_n_81__52_,
  r_n_81__51_,r_n_81__50_,r_n_81__49_,r_n_81__48_,r_n_81__47_,r_n_81__46_,r_n_81__45_,
  r_n_81__44_,r_n_81__43_,r_n_81__42_,r_n_81__41_,r_n_81__40_,r_n_81__39_,r_n_81__38_,
  r_n_81__37_,r_n_81__36_,r_n_81__35_,r_n_81__34_,r_n_81__33_,r_n_81__32_,
  r_n_81__31_,r_n_81__30_,r_n_81__29_,r_n_81__28_,r_n_81__27_,r_n_81__26_,r_n_81__25_,
  r_n_81__24_,r_n_81__23_,r_n_81__22_,r_n_81__21_,r_n_81__20_,r_n_81__19_,r_n_81__18_,
  r_n_81__17_,r_n_81__16_,r_n_81__15_,r_n_81__14_,r_n_81__13_,r_n_81__12_,
  r_n_81__11_,r_n_81__10_,r_n_81__9_,r_n_81__8_,r_n_81__7_,r_n_81__6_,r_n_81__5_,
  r_n_81__4_,r_n_81__3_,r_n_81__2_,r_n_81__1_,r_n_81__0_,r_n_96__63_,r_n_96__62_,
  r_n_96__61_,r_n_96__60_,r_n_96__59_,r_n_96__58_,r_n_96__57_,r_n_96__56_,r_n_96__55_,
  r_n_96__54_,r_n_96__53_,r_n_96__52_,r_n_96__51_,r_n_96__50_,r_n_96__49_,r_n_96__48_,
  r_n_96__47_,r_n_96__46_,r_n_96__45_,r_n_96__44_,r_n_96__43_,r_n_96__42_,
  r_n_96__41_,r_n_96__40_,r_n_96__39_,r_n_96__38_,r_n_96__37_,r_n_96__36_,r_n_96__35_,
  r_n_96__34_,r_n_96__33_,r_n_96__32_,r_n_96__31_,r_n_96__30_,r_n_96__29_,r_n_96__28_,
  r_n_96__27_,r_n_96__26_,r_n_96__25_,r_n_96__24_,r_n_96__23_,r_n_96__22_,
  r_n_96__21_,r_n_96__20_,r_n_96__19_,r_n_96__18_,r_n_96__17_,r_n_96__16_,r_n_96__15_,
  r_n_96__14_,r_n_96__13_,r_n_96__12_,r_n_96__11_,r_n_96__10_,r_n_96__9_,r_n_96__8_,
  r_n_96__7_,r_n_96__6_,r_n_96__5_,r_n_96__4_,r_n_96__3_,r_n_96__2_,r_n_96__1_,
  r_n_96__0_,r_n_95__63_,r_n_95__62_,r_n_95__61_,r_n_95__60_,r_n_95__59_,r_n_95__58_,
  r_n_95__57_,r_n_95__56_,r_n_95__55_,r_n_95__54_,r_n_95__53_,r_n_95__52_,r_n_95__51_,
  r_n_95__50_,r_n_95__49_,r_n_95__48_,r_n_95__47_,r_n_95__46_,r_n_95__45_,
  r_n_95__44_,r_n_95__43_,r_n_95__42_,r_n_95__41_,r_n_95__40_,r_n_95__39_,r_n_95__38_,
  r_n_95__37_,r_n_95__36_,r_n_95__35_,r_n_95__34_,r_n_95__33_,r_n_95__32_,r_n_95__31_,
  r_n_95__30_,r_n_95__29_,r_n_95__28_,r_n_95__27_,r_n_95__26_,r_n_95__25_,
  r_n_95__24_,r_n_95__23_,r_n_95__22_,r_n_95__21_,r_n_95__20_,r_n_95__19_,r_n_95__18_,
  r_n_95__17_,r_n_95__16_,r_n_95__15_,r_n_95__14_,r_n_95__13_,r_n_95__12_,r_n_95__11_,
  r_n_95__10_,r_n_95__9_,r_n_95__8_,r_n_95__7_,r_n_95__6_,r_n_95__5_,r_n_95__4_,
  r_n_95__3_,r_n_95__2_,r_n_95__1_,r_n_95__0_,r_n_94__63_,r_n_94__62_,r_n_94__61_,
  r_n_94__60_,r_n_94__59_,r_n_94__58_,r_n_94__57_,r_n_94__56_,r_n_94__55_,
  r_n_94__54_,r_n_94__53_,r_n_94__52_,r_n_94__51_,r_n_94__50_,r_n_94__49_,r_n_94__48_,
  r_n_94__47_,r_n_94__46_,r_n_94__45_,r_n_94__44_,r_n_94__43_,r_n_94__42_,r_n_94__41_,
  r_n_94__40_,r_n_94__39_,r_n_94__38_,r_n_94__37_,r_n_94__36_,r_n_94__35_,
  r_n_94__34_,r_n_94__33_,r_n_94__32_,r_n_94__31_,r_n_94__30_,r_n_94__29_,r_n_94__28_,
  r_n_94__27_,r_n_94__26_,r_n_94__25_,r_n_94__24_,r_n_94__23_,r_n_94__22_,r_n_94__21_,
  r_n_94__20_,r_n_94__19_,r_n_94__18_,r_n_94__17_,r_n_94__16_,r_n_94__15_,
  r_n_94__14_,r_n_94__13_,r_n_94__12_,r_n_94__11_,r_n_94__10_,r_n_94__9_,r_n_94__8_,
  r_n_94__7_,r_n_94__6_,r_n_94__5_,r_n_94__4_,r_n_94__3_,r_n_94__2_,r_n_94__1_,r_n_94__0_,
  r_n_93__63_,r_n_93__62_,r_n_93__61_,r_n_93__60_,r_n_93__59_,r_n_93__58_,
  r_n_93__57_,r_n_93__56_,r_n_93__55_,r_n_93__54_,r_n_93__53_,r_n_93__52_,r_n_93__51_,
  r_n_93__50_,r_n_93__49_,r_n_93__48_,r_n_93__47_,r_n_93__46_,r_n_93__45_,r_n_93__44_,
  r_n_93__43_,r_n_93__42_,r_n_93__41_,r_n_93__40_,r_n_93__39_,r_n_93__38_,
  r_n_93__37_,r_n_93__36_,r_n_93__35_,r_n_93__34_,r_n_93__33_,r_n_93__32_,r_n_93__31_,
  r_n_93__30_,r_n_93__29_,r_n_93__28_,r_n_93__27_,r_n_93__26_,r_n_93__25_,r_n_93__24_,
  r_n_93__23_,r_n_93__22_,r_n_93__21_,r_n_93__20_,r_n_93__19_,r_n_93__18_,
  r_n_93__17_,r_n_93__16_,r_n_93__15_,r_n_93__14_,r_n_93__13_,r_n_93__12_,r_n_93__11_,
  r_n_93__10_,r_n_93__9_,r_n_93__8_,r_n_93__7_,r_n_93__6_,r_n_93__5_,r_n_93__4_,
  r_n_93__3_,r_n_93__2_,r_n_93__1_,r_n_93__0_,r_n_92__63_,r_n_92__62_,r_n_92__61_,
  r_n_92__60_,r_n_92__59_,r_n_92__58_,r_n_92__57_,r_n_92__56_,r_n_92__55_,r_n_92__54_,
  r_n_92__53_,r_n_92__52_,r_n_92__51_,r_n_92__50_,r_n_92__49_,r_n_92__48_,
  r_n_92__47_,r_n_92__46_,r_n_92__45_,r_n_92__44_,r_n_92__43_,r_n_92__42_,r_n_92__41_,
  r_n_92__40_,r_n_92__39_,r_n_92__38_,r_n_92__37_,r_n_92__36_,r_n_92__35_,r_n_92__34_,
  r_n_92__33_,r_n_92__32_,r_n_92__31_,r_n_92__30_,r_n_92__29_,r_n_92__28_,
  r_n_92__27_,r_n_92__26_,r_n_92__25_,r_n_92__24_,r_n_92__23_,r_n_92__22_,r_n_92__21_,
  r_n_92__20_,r_n_92__19_,r_n_92__18_,r_n_92__17_,r_n_92__16_,r_n_92__15_,r_n_92__14_,
  r_n_92__13_,r_n_92__12_,r_n_92__11_,r_n_92__10_,r_n_92__9_,r_n_92__8_,r_n_92__7_,
  r_n_92__6_,r_n_92__5_,r_n_92__4_,r_n_92__3_,r_n_92__2_,r_n_92__1_,r_n_92__0_,
  r_n_91__63_,r_n_91__62_,r_n_91__61_,r_n_91__60_,r_n_91__59_,r_n_91__58_,r_n_91__57_,
  r_n_91__56_,r_n_91__55_,r_n_91__54_,r_n_91__53_,r_n_91__52_,r_n_91__51_,
  r_n_91__50_,r_n_91__49_,r_n_91__48_,r_n_91__47_,r_n_91__46_,r_n_91__45_,r_n_91__44_,
  r_n_91__43_,r_n_91__42_,r_n_91__41_,r_n_91__40_,r_n_91__39_,r_n_91__38_,r_n_91__37_,
  r_n_91__36_,r_n_91__35_,r_n_91__34_,r_n_91__33_,r_n_91__32_,r_n_91__31_,
  r_n_91__30_,r_n_91__29_,r_n_91__28_,r_n_91__27_,r_n_91__26_,r_n_91__25_,r_n_91__24_,
  r_n_91__23_,r_n_91__22_,r_n_91__21_,r_n_91__20_,r_n_91__19_,r_n_91__18_,r_n_91__17_,
  r_n_91__16_,r_n_91__15_,r_n_91__14_,r_n_91__13_,r_n_91__12_,r_n_91__11_,
  r_n_91__10_,r_n_91__9_,r_n_91__8_,r_n_91__7_,r_n_91__6_,r_n_91__5_,r_n_91__4_,
  r_n_91__3_,r_n_91__2_,r_n_91__1_,r_n_91__0_,r_n_90__63_,r_n_90__62_,r_n_90__61_,
  r_n_90__60_,r_n_90__59_,r_n_90__58_,r_n_90__57_,r_n_90__56_,r_n_90__55_,r_n_90__54_,
  r_n_90__53_,r_n_90__52_,r_n_90__51_,r_n_90__50_,r_n_90__49_,r_n_90__48_,r_n_90__47_,
  r_n_90__46_,r_n_90__45_,r_n_90__44_,r_n_90__43_,r_n_90__42_,r_n_90__41_,
  r_n_90__40_,r_n_90__39_,r_n_90__38_,r_n_90__37_,r_n_90__36_,r_n_90__35_,r_n_90__34_,
  r_n_90__33_,r_n_90__32_,r_n_90__31_,r_n_90__30_,r_n_90__29_,r_n_90__28_,r_n_90__27_,
  r_n_90__26_,r_n_90__25_,r_n_90__24_,r_n_90__23_,r_n_90__22_,r_n_90__21_,
  r_n_90__20_,r_n_90__19_,r_n_90__18_,r_n_90__17_,r_n_90__16_,r_n_90__15_,r_n_90__14_,
  r_n_90__13_,r_n_90__12_,r_n_90__11_,r_n_90__10_,r_n_90__9_,r_n_90__8_,r_n_90__7_,
  r_n_90__6_,r_n_90__5_,r_n_90__4_,r_n_90__3_,r_n_90__2_,r_n_90__1_,r_n_90__0_,
  r_n_89__63_,r_n_89__62_,r_n_89__61_,r_n_89__60_,r_n_89__59_,r_n_89__58_,r_n_89__57_,
  r_n_89__56_,r_n_89__55_,r_n_89__54_,r_n_89__53_,r_n_89__52_,r_n_89__51_,r_n_89__50_,
  r_n_89__49_,r_n_89__48_,r_n_89__47_,r_n_89__46_,r_n_89__45_,r_n_89__44_,
  r_n_89__43_,r_n_89__42_,r_n_89__41_,r_n_89__40_,r_n_89__39_,r_n_89__38_,r_n_89__37_,
  r_n_89__36_,r_n_89__35_,r_n_89__34_,r_n_89__33_,r_n_89__32_,r_n_89__31_,r_n_89__30_,
  r_n_89__29_,r_n_89__28_,r_n_89__27_,r_n_89__26_,r_n_89__25_,r_n_89__24_,
  r_n_89__23_,r_n_89__22_,r_n_89__21_,r_n_89__20_,r_n_89__19_,r_n_89__18_,r_n_89__17_,
  r_n_89__16_,r_n_89__15_,r_n_89__14_,r_n_89__13_,r_n_89__12_,r_n_89__11_,r_n_89__10_,
  r_n_89__9_,r_n_89__8_,r_n_89__7_,r_n_89__6_,r_n_89__5_,r_n_89__4_,r_n_89__3_,
  r_n_89__2_,r_n_89__1_,r_n_89__0_,r_n_104__63_,r_n_104__62_,r_n_104__61_,
  r_n_104__60_,r_n_104__59_,r_n_104__58_,r_n_104__57_,r_n_104__56_,r_n_104__55_,r_n_104__54_,
  r_n_104__53_,r_n_104__52_,r_n_104__51_,r_n_104__50_,r_n_104__49_,r_n_104__48_,
  r_n_104__47_,r_n_104__46_,r_n_104__45_,r_n_104__44_,r_n_104__43_,r_n_104__42_,
  r_n_104__41_,r_n_104__40_,r_n_104__39_,r_n_104__38_,r_n_104__37_,r_n_104__36_,
  r_n_104__35_,r_n_104__34_,r_n_104__33_,r_n_104__32_,r_n_104__31_,r_n_104__30_,
  r_n_104__29_,r_n_104__28_,r_n_104__27_,r_n_104__26_,r_n_104__25_,r_n_104__24_,
  r_n_104__23_,r_n_104__22_,r_n_104__21_,r_n_104__20_,r_n_104__19_,r_n_104__18_,
  r_n_104__17_,r_n_104__16_,r_n_104__15_,r_n_104__14_,r_n_104__13_,r_n_104__12_,r_n_104__11_,
  r_n_104__10_,r_n_104__9_,r_n_104__8_,r_n_104__7_,r_n_104__6_,r_n_104__5_,
  r_n_104__4_,r_n_104__3_,r_n_104__2_,r_n_104__1_,r_n_104__0_,r_n_103__63_,r_n_103__62_,
  r_n_103__61_,r_n_103__60_,r_n_103__59_,r_n_103__58_,r_n_103__57_,r_n_103__56_,
  r_n_103__55_,r_n_103__54_,r_n_103__53_,r_n_103__52_,r_n_103__51_,r_n_103__50_,
  r_n_103__49_,r_n_103__48_,r_n_103__47_,r_n_103__46_,r_n_103__45_,r_n_103__44_,
  r_n_103__43_,r_n_103__42_,r_n_103__41_,r_n_103__40_,r_n_103__39_,r_n_103__38_,
  r_n_103__37_,r_n_103__36_,r_n_103__35_,r_n_103__34_,r_n_103__33_,r_n_103__32_,
  r_n_103__31_,r_n_103__30_,r_n_103__29_,r_n_103__28_,r_n_103__27_,r_n_103__26_,r_n_103__25_,
  r_n_103__24_,r_n_103__23_,r_n_103__22_,r_n_103__21_,r_n_103__20_,r_n_103__19_,
  r_n_103__18_,r_n_103__17_,r_n_103__16_,r_n_103__15_,r_n_103__14_,r_n_103__13_,
  r_n_103__12_,r_n_103__11_,r_n_103__10_,r_n_103__9_,r_n_103__8_,r_n_103__7_,
  r_n_103__6_,r_n_103__5_,r_n_103__4_,r_n_103__3_,r_n_103__2_,r_n_103__1_,r_n_103__0_,
  r_n_102__63_,r_n_102__62_,r_n_102__61_,r_n_102__60_,r_n_102__59_,r_n_102__58_,
  r_n_102__57_,r_n_102__56_,r_n_102__55_,r_n_102__54_,r_n_102__53_,r_n_102__52_,
  r_n_102__51_,r_n_102__50_,r_n_102__49_,r_n_102__48_,r_n_102__47_,r_n_102__46_,
  r_n_102__45_,r_n_102__44_,r_n_102__43_,r_n_102__42_,r_n_102__41_,r_n_102__40_,r_n_102__39_,
  r_n_102__38_,r_n_102__37_,r_n_102__36_,r_n_102__35_,r_n_102__34_,r_n_102__33_,
  r_n_102__32_,r_n_102__31_,r_n_102__30_,r_n_102__29_,r_n_102__28_,r_n_102__27_,
  r_n_102__26_,r_n_102__25_,r_n_102__24_,r_n_102__23_,r_n_102__22_,r_n_102__21_,
  r_n_102__20_,r_n_102__19_,r_n_102__18_,r_n_102__17_,r_n_102__16_,r_n_102__15_,
  r_n_102__14_,r_n_102__13_,r_n_102__12_,r_n_102__11_,r_n_102__10_,r_n_102__9_,r_n_102__8_,
  r_n_102__7_,r_n_102__6_,r_n_102__5_,r_n_102__4_,r_n_102__3_,r_n_102__2_,
  r_n_102__1_,r_n_102__0_,r_n_101__63_,r_n_101__62_,r_n_101__61_,r_n_101__60_,
  r_n_101__59_,r_n_101__58_,r_n_101__57_,r_n_101__56_,r_n_101__55_,r_n_101__54_,r_n_101__53_,
  r_n_101__52_,r_n_101__51_,r_n_101__50_,r_n_101__49_,r_n_101__48_,r_n_101__47_,
  r_n_101__46_,r_n_101__45_,r_n_101__44_,r_n_101__43_,r_n_101__42_,r_n_101__41_,
  r_n_101__40_,r_n_101__39_,r_n_101__38_,r_n_101__37_,r_n_101__36_,r_n_101__35_,
  r_n_101__34_,r_n_101__33_,r_n_101__32_,r_n_101__31_,r_n_101__30_,r_n_101__29_,
  r_n_101__28_,r_n_101__27_,r_n_101__26_,r_n_101__25_,r_n_101__24_,r_n_101__23_,
  r_n_101__22_,r_n_101__21_,r_n_101__20_,r_n_101__19_,r_n_101__18_,r_n_101__17_,r_n_101__16_,
  r_n_101__15_,r_n_101__14_,r_n_101__13_,r_n_101__12_,r_n_101__11_,r_n_101__10_,
  r_n_101__9_,r_n_101__8_,r_n_101__7_,r_n_101__6_,r_n_101__5_,r_n_101__4_,
  r_n_101__3_,r_n_101__2_,r_n_101__1_,r_n_101__0_,r_n_100__63_,r_n_100__62_,r_n_100__61_,
  r_n_100__60_,r_n_100__59_,r_n_100__58_,r_n_100__57_,r_n_100__56_,r_n_100__55_,
  r_n_100__54_,r_n_100__53_,r_n_100__52_,r_n_100__51_,r_n_100__50_,r_n_100__49_,
  r_n_100__48_,r_n_100__47_,r_n_100__46_,r_n_100__45_,r_n_100__44_,r_n_100__43_,
  r_n_100__42_,r_n_100__41_,r_n_100__40_,r_n_100__39_,r_n_100__38_,r_n_100__37_,
  r_n_100__36_,r_n_100__35_,r_n_100__34_,r_n_100__33_,r_n_100__32_,r_n_100__31_,r_n_100__30_,
  r_n_100__29_,r_n_100__28_,r_n_100__27_,r_n_100__26_,r_n_100__25_,r_n_100__24_,
  r_n_100__23_,r_n_100__22_,r_n_100__21_,r_n_100__20_,r_n_100__19_,r_n_100__18_,
  r_n_100__17_,r_n_100__16_,r_n_100__15_,r_n_100__14_,r_n_100__13_,r_n_100__12_,
  r_n_100__11_,r_n_100__10_,r_n_100__9_,r_n_100__8_,r_n_100__7_,r_n_100__6_,r_n_100__5_,
  r_n_100__4_,r_n_100__3_,r_n_100__2_,r_n_100__1_,r_n_100__0_,r_n_99__63_,
  r_n_99__62_,r_n_99__61_,r_n_99__60_,r_n_99__59_,r_n_99__58_,r_n_99__57_,r_n_99__56_,
  r_n_99__55_,r_n_99__54_,r_n_99__53_,r_n_99__52_,r_n_99__51_,r_n_99__50_,r_n_99__49_,
  r_n_99__48_,r_n_99__47_,r_n_99__46_,r_n_99__45_,r_n_99__44_,r_n_99__43_,
  r_n_99__42_,r_n_99__41_,r_n_99__40_,r_n_99__39_,r_n_99__38_,r_n_99__37_,r_n_99__36_,
  r_n_99__35_,r_n_99__34_,r_n_99__33_,r_n_99__32_,r_n_99__31_,r_n_99__30_,r_n_99__29_,
  r_n_99__28_,r_n_99__27_,r_n_99__26_,r_n_99__25_,r_n_99__24_,r_n_99__23_,
  r_n_99__22_,r_n_99__21_,r_n_99__20_,r_n_99__19_,r_n_99__18_,r_n_99__17_,r_n_99__16_,
  r_n_99__15_,r_n_99__14_,r_n_99__13_,r_n_99__12_,r_n_99__11_,r_n_99__10_,r_n_99__9_,
  r_n_99__8_,r_n_99__7_,r_n_99__6_,r_n_99__5_,r_n_99__4_,r_n_99__3_,r_n_99__2_,
  r_n_99__1_,r_n_99__0_,r_n_98__63_,r_n_98__62_,r_n_98__61_,r_n_98__60_,r_n_98__59_,
  r_n_98__58_,r_n_98__57_,r_n_98__56_,r_n_98__55_,r_n_98__54_,r_n_98__53_,
  r_n_98__52_,r_n_98__51_,r_n_98__50_,r_n_98__49_,r_n_98__48_,r_n_98__47_,r_n_98__46_,
  r_n_98__45_,r_n_98__44_,r_n_98__43_,r_n_98__42_,r_n_98__41_,r_n_98__40_,r_n_98__39_,
  r_n_98__38_,r_n_98__37_,r_n_98__36_,r_n_98__35_,r_n_98__34_,r_n_98__33_,
  r_n_98__32_,r_n_98__31_,r_n_98__30_,r_n_98__29_,r_n_98__28_,r_n_98__27_,r_n_98__26_,
  r_n_98__25_,r_n_98__24_,r_n_98__23_,r_n_98__22_,r_n_98__21_,r_n_98__20_,r_n_98__19_,
  r_n_98__18_,r_n_98__17_,r_n_98__16_,r_n_98__15_,r_n_98__14_,r_n_98__13_,
  r_n_98__12_,r_n_98__11_,r_n_98__10_,r_n_98__9_,r_n_98__8_,r_n_98__7_,r_n_98__6_,
  r_n_98__5_,r_n_98__4_,r_n_98__3_,r_n_98__2_,r_n_98__1_,r_n_98__0_,r_n_97__63_,r_n_97__62_,
  r_n_97__61_,r_n_97__60_,r_n_97__59_,r_n_97__58_,r_n_97__57_,r_n_97__56_,
  r_n_97__55_,r_n_97__54_,r_n_97__53_,r_n_97__52_,r_n_97__51_,r_n_97__50_,r_n_97__49_,
  r_n_97__48_,r_n_97__47_,r_n_97__46_,r_n_97__45_,r_n_97__44_,r_n_97__43_,r_n_97__42_,
  r_n_97__41_,r_n_97__40_,r_n_97__39_,r_n_97__38_,r_n_97__37_,r_n_97__36_,
  r_n_97__35_,r_n_97__34_,r_n_97__33_,r_n_97__32_,r_n_97__31_,r_n_97__30_,r_n_97__29_,
  r_n_97__28_,r_n_97__27_,r_n_97__26_,r_n_97__25_,r_n_97__24_,r_n_97__23_,r_n_97__22_,
  r_n_97__21_,r_n_97__20_,r_n_97__19_,r_n_97__18_,r_n_97__17_,r_n_97__16_,
  r_n_97__15_,r_n_97__14_,r_n_97__13_,r_n_97__12_,r_n_97__11_,r_n_97__10_,r_n_97__9_,
  r_n_97__8_,r_n_97__7_,r_n_97__6_,r_n_97__5_,r_n_97__4_,r_n_97__3_,r_n_97__2_,
  r_n_97__1_,r_n_97__0_,r_n_112__63_,r_n_112__62_,r_n_112__61_,r_n_112__60_,r_n_112__59_,
  r_n_112__58_,r_n_112__57_,r_n_112__56_,r_n_112__55_,r_n_112__54_,r_n_112__53_,
  r_n_112__52_,r_n_112__51_,r_n_112__50_,r_n_112__49_,r_n_112__48_,r_n_112__47_,
  r_n_112__46_,r_n_112__45_,r_n_112__44_,r_n_112__43_,r_n_112__42_,r_n_112__41_,
  r_n_112__40_,r_n_112__39_,r_n_112__38_,r_n_112__37_,r_n_112__36_,r_n_112__35_,
  r_n_112__34_,r_n_112__33_,r_n_112__32_,r_n_112__31_,r_n_112__30_,r_n_112__29_,
  r_n_112__28_,r_n_112__27_,r_n_112__26_,r_n_112__25_,r_n_112__24_,r_n_112__23_,r_n_112__22_,
  r_n_112__21_,r_n_112__20_,r_n_112__19_,r_n_112__18_,r_n_112__17_,r_n_112__16_,
  r_n_112__15_,r_n_112__14_,r_n_112__13_,r_n_112__12_,r_n_112__11_,r_n_112__10_,
  r_n_112__9_,r_n_112__8_,r_n_112__7_,r_n_112__6_,r_n_112__5_,r_n_112__4_,r_n_112__3_,
  r_n_112__2_,r_n_112__1_,r_n_112__0_,r_n_111__63_,r_n_111__62_,r_n_111__61_,
  r_n_111__60_,r_n_111__59_,r_n_111__58_,r_n_111__57_,r_n_111__56_,r_n_111__55_,
  r_n_111__54_,r_n_111__53_,r_n_111__52_,r_n_111__51_,r_n_111__50_,r_n_111__49_,
  r_n_111__48_,r_n_111__47_,r_n_111__46_,r_n_111__45_,r_n_111__44_,r_n_111__43_,
  r_n_111__42_,r_n_111__41_,r_n_111__40_,r_n_111__39_,r_n_111__38_,r_n_111__37_,r_n_111__36_,
  r_n_111__35_,r_n_111__34_,r_n_111__33_,r_n_111__32_,r_n_111__31_,r_n_111__30_,
  r_n_111__29_,r_n_111__28_,r_n_111__27_,r_n_111__26_,r_n_111__25_,r_n_111__24_,
  r_n_111__23_,r_n_111__22_,r_n_111__21_,r_n_111__20_,r_n_111__19_,r_n_111__18_,
  r_n_111__17_,r_n_111__16_,r_n_111__15_,r_n_111__14_,r_n_111__13_,r_n_111__12_,
  r_n_111__11_,r_n_111__10_,r_n_111__9_,r_n_111__8_,r_n_111__7_,r_n_111__6_,r_n_111__5_,
  r_n_111__4_,r_n_111__3_,r_n_111__2_,r_n_111__1_,r_n_111__0_,r_n_110__63_,
  r_n_110__62_,r_n_110__61_,r_n_110__60_,r_n_110__59_,r_n_110__58_,r_n_110__57_,
  r_n_110__56_,r_n_110__55_,r_n_110__54_,r_n_110__53_,r_n_110__52_,r_n_110__51_,r_n_110__50_,
  r_n_110__49_,r_n_110__48_,r_n_110__47_,r_n_110__46_,r_n_110__45_,r_n_110__44_,
  r_n_110__43_,r_n_110__42_,r_n_110__41_,r_n_110__40_,r_n_110__39_,r_n_110__38_,
  r_n_110__37_,r_n_110__36_,r_n_110__35_,r_n_110__34_,r_n_110__33_,r_n_110__32_,
  r_n_110__31_,r_n_110__30_,r_n_110__29_,r_n_110__28_,r_n_110__27_,r_n_110__26_,
  r_n_110__25_,r_n_110__24_,r_n_110__23_,r_n_110__22_,r_n_110__21_,r_n_110__20_,
  r_n_110__19_,r_n_110__18_,r_n_110__17_,r_n_110__16_,r_n_110__15_,r_n_110__14_,
  r_n_110__13_,r_n_110__12_,r_n_110__11_,r_n_110__10_,r_n_110__9_,r_n_110__8_,r_n_110__7_,
  r_n_110__6_,r_n_110__5_,r_n_110__4_,r_n_110__3_,r_n_110__2_,r_n_110__1_,r_n_110__0_,
  r_n_109__63_,r_n_109__62_,r_n_109__61_,r_n_109__60_,r_n_109__59_,r_n_109__58_,
  r_n_109__57_,r_n_109__56_,r_n_109__55_,r_n_109__54_,r_n_109__53_,r_n_109__52_,
  r_n_109__51_,r_n_109__50_,r_n_109__49_,r_n_109__48_,r_n_109__47_,r_n_109__46_,
  r_n_109__45_,r_n_109__44_,r_n_109__43_,r_n_109__42_,r_n_109__41_,r_n_109__40_,
  r_n_109__39_,r_n_109__38_,r_n_109__37_,r_n_109__36_,r_n_109__35_,r_n_109__34_,
  r_n_109__33_,r_n_109__32_,r_n_109__31_,r_n_109__30_,r_n_109__29_,r_n_109__28_,
  r_n_109__27_,r_n_109__26_,r_n_109__25_,r_n_109__24_,r_n_109__23_,r_n_109__22_,r_n_109__21_,
  r_n_109__20_,r_n_109__19_,r_n_109__18_,r_n_109__17_,r_n_109__16_,r_n_109__15_,
  r_n_109__14_,r_n_109__13_,r_n_109__12_,r_n_109__11_,r_n_109__10_,r_n_109__9_,
  r_n_109__8_,r_n_109__7_,r_n_109__6_,r_n_109__5_,r_n_109__4_,r_n_109__3_,r_n_109__2_,
  r_n_109__1_,r_n_109__0_,r_n_108__63_,r_n_108__62_,r_n_108__61_,r_n_108__60_,
  r_n_108__59_,r_n_108__58_,r_n_108__57_,r_n_108__56_,r_n_108__55_,r_n_108__54_,
  r_n_108__53_,r_n_108__52_,r_n_108__51_,r_n_108__50_,r_n_108__49_,r_n_108__48_,
  r_n_108__47_,r_n_108__46_,r_n_108__45_,r_n_108__44_,r_n_108__43_,r_n_108__42_,
  r_n_108__41_,r_n_108__40_,r_n_108__39_,r_n_108__38_,r_n_108__37_,r_n_108__36_,r_n_108__35_,
  r_n_108__34_,r_n_108__33_,r_n_108__32_,r_n_108__31_,r_n_108__30_,r_n_108__29_,
  r_n_108__28_,r_n_108__27_,r_n_108__26_,r_n_108__25_,r_n_108__24_,r_n_108__23_,
  r_n_108__22_,r_n_108__21_,r_n_108__20_,r_n_108__19_,r_n_108__18_,r_n_108__17_,
  r_n_108__16_,r_n_108__15_,r_n_108__14_,r_n_108__13_,r_n_108__12_,r_n_108__11_,
  r_n_108__10_,r_n_108__9_,r_n_108__8_,r_n_108__7_,r_n_108__6_,r_n_108__5_,r_n_108__4_,
  r_n_108__3_,r_n_108__2_,r_n_108__1_,r_n_108__0_,r_n_107__63_,r_n_107__62_,
  r_n_107__61_,r_n_107__60_,r_n_107__59_,r_n_107__58_,r_n_107__57_,r_n_107__56_,
  r_n_107__55_,r_n_107__54_,r_n_107__53_,r_n_107__52_,r_n_107__51_,r_n_107__50_,r_n_107__49_,
  r_n_107__48_,r_n_107__47_,r_n_107__46_,r_n_107__45_,r_n_107__44_,r_n_107__43_,
  r_n_107__42_,r_n_107__41_,r_n_107__40_,r_n_107__39_,r_n_107__38_,r_n_107__37_,
  r_n_107__36_,r_n_107__35_,r_n_107__34_,r_n_107__33_,r_n_107__32_,r_n_107__31_,
  r_n_107__30_,r_n_107__29_,r_n_107__28_,r_n_107__27_,r_n_107__26_,r_n_107__25_,
  r_n_107__24_,r_n_107__23_,r_n_107__22_,r_n_107__21_,r_n_107__20_,r_n_107__19_,
  r_n_107__18_,r_n_107__17_,r_n_107__16_,r_n_107__15_,r_n_107__14_,r_n_107__13_,r_n_107__12_,
  r_n_107__11_,r_n_107__10_,r_n_107__9_,r_n_107__8_,r_n_107__7_,r_n_107__6_,
  r_n_107__5_,r_n_107__4_,r_n_107__3_,r_n_107__2_,r_n_107__1_,r_n_107__0_,r_n_106__63_,
  r_n_106__62_,r_n_106__61_,r_n_106__60_,r_n_106__59_,r_n_106__58_,r_n_106__57_,
  r_n_106__56_,r_n_106__55_,r_n_106__54_,r_n_106__53_,r_n_106__52_,r_n_106__51_,
  r_n_106__50_,r_n_106__49_,r_n_106__48_,r_n_106__47_,r_n_106__46_,r_n_106__45_,
  r_n_106__44_,r_n_106__43_,r_n_106__42_,r_n_106__41_,r_n_106__40_,r_n_106__39_,
  r_n_106__38_,r_n_106__37_,r_n_106__36_,r_n_106__35_,r_n_106__34_,r_n_106__33_,
  r_n_106__32_,r_n_106__31_,r_n_106__30_,r_n_106__29_,r_n_106__28_,r_n_106__27_,r_n_106__26_,
  r_n_106__25_,r_n_106__24_,r_n_106__23_,r_n_106__22_,r_n_106__21_,r_n_106__20_,
  r_n_106__19_,r_n_106__18_,r_n_106__17_,r_n_106__16_,r_n_106__15_,r_n_106__14_,
  r_n_106__13_,r_n_106__12_,r_n_106__11_,r_n_106__10_,r_n_106__9_,r_n_106__8_,
  r_n_106__7_,r_n_106__6_,r_n_106__5_,r_n_106__4_,r_n_106__3_,r_n_106__2_,r_n_106__1_,
  r_n_106__0_,r_n_105__63_,r_n_105__62_,r_n_105__61_,r_n_105__60_,r_n_105__59_,
  r_n_105__58_,r_n_105__57_,r_n_105__56_,r_n_105__55_,r_n_105__54_,r_n_105__53_,
  r_n_105__52_,r_n_105__51_,r_n_105__50_,r_n_105__49_,r_n_105__48_,r_n_105__47_,
  r_n_105__46_,r_n_105__45_,r_n_105__44_,r_n_105__43_,r_n_105__42_,r_n_105__41_,r_n_105__40_,
  r_n_105__39_,r_n_105__38_,r_n_105__37_,r_n_105__36_,r_n_105__35_,r_n_105__34_,
  r_n_105__33_,r_n_105__32_,r_n_105__31_,r_n_105__30_,r_n_105__29_,r_n_105__28_,
  r_n_105__27_,r_n_105__26_,r_n_105__25_,r_n_105__24_,r_n_105__23_,r_n_105__22_,
  r_n_105__21_,r_n_105__20_,r_n_105__19_,r_n_105__18_,r_n_105__17_,r_n_105__16_,
  r_n_105__15_,r_n_105__14_,r_n_105__13_,r_n_105__12_,r_n_105__11_,r_n_105__10_,
  r_n_105__9_,r_n_105__8_,r_n_105__7_,r_n_105__6_,r_n_105__5_,r_n_105__4_,r_n_105__3_,
  r_n_105__2_,r_n_105__1_,r_n_105__0_,r_n_120__63_,r_n_120__62_,r_n_120__61_,
  r_n_120__60_,r_n_120__59_,r_n_120__58_,r_n_120__57_,r_n_120__56_,r_n_120__55_,r_n_120__54_,
  r_n_120__53_,r_n_120__52_,r_n_120__51_,r_n_120__50_,r_n_120__49_,r_n_120__48_,
  r_n_120__47_,r_n_120__46_,r_n_120__45_,r_n_120__44_,r_n_120__43_,r_n_120__42_,
  r_n_120__41_,r_n_120__40_,r_n_120__39_,r_n_120__38_,r_n_120__37_,r_n_120__36_,
  r_n_120__35_,r_n_120__34_,r_n_120__33_,r_n_120__32_,r_n_120__31_,r_n_120__30_,
  r_n_120__29_,r_n_120__28_,r_n_120__27_,r_n_120__26_,r_n_120__25_,r_n_120__24_,
  r_n_120__23_,r_n_120__22_,r_n_120__21_,r_n_120__20_,r_n_120__19_,r_n_120__18_,
  r_n_120__17_,r_n_120__16_,r_n_120__15_,r_n_120__14_,r_n_120__13_,r_n_120__12_,r_n_120__11_,
  r_n_120__10_,r_n_120__9_,r_n_120__8_,r_n_120__7_,r_n_120__6_,r_n_120__5_,
  r_n_120__4_,r_n_120__3_,r_n_120__2_,r_n_120__1_,r_n_120__0_,r_n_119__63_,r_n_119__62_,
  r_n_119__61_,r_n_119__60_,r_n_119__59_,r_n_119__58_,r_n_119__57_,r_n_119__56_,
  r_n_119__55_,r_n_119__54_,r_n_119__53_,r_n_119__52_,r_n_119__51_,r_n_119__50_,
  r_n_119__49_,r_n_119__48_,r_n_119__47_,r_n_119__46_,r_n_119__45_,r_n_119__44_,
  r_n_119__43_,r_n_119__42_,r_n_119__41_,r_n_119__40_,r_n_119__39_,r_n_119__38_,
  r_n_119__37_,r_n_119__36_,r_n_119__35_,r_n_119__34_,r_n_119__33_,r_n_119__32_,
  r_n_119__31_,r_n_119__30_,r_n_119__29_,r_n_119__28_,r_n_119__27_,r_n_119__26_,r_n_119__25_,
  r_n_119__24_,r_n_119__23_,r_n_119__22_,r_n_119__21_,r_n_119__20_,r_n_119__19_,
  r_n_119__18_,r_n_119__17_,r_n_119__16_,r_n_119__15_,r_n_119__14_,r_n_119__13_,
  r_n_119__12_,r_n_119__11_,r_n_119__10_,r_n_119__9_,r_n_119__8_,r_n_119__7_,
  r_n_119__6_,r_n_119__5_,r_n_119__4_,r_n_119__3_,r_n_119__2_,r_n_119__1_,r_n_119__0_,
  r_n_118__63_,r_n_118__62_,r_n_118__61_,r_n_118__60_,r_n_118__59_,r_n_118__58_,
  r_n_118__57_,r_n_118__56_,r_n_118__55_,r_n_118__54_,r_n_118__53_,r_n_118__52_,
  r_n_118__51_,r_n_118__50_,r_n_118__49_,r_n_118__48_,r_n_118__47_,r_n_118__46_,
  r_n_118__45_,r_n_118__44_,r_n_118__43_,r_n_118__42_,r_n_118__41_,r_n_118__40_,r_n_118__39_,
  r_n_118__38_,r_n_118__37_,r_n_118__36_,r_n_118__35_,r_n_118__34_,r_n_118__33_,
  r_n_118__32_,r_n_118__31_,r_n_118__30_,r_n_118__29_,r_n_118__28_,r_n_118__27_,
  r_n_118__26_,r_n_118__25_,r_n_118__24_,r_n_118__23_,r_n_118__22_,r_n_118__21_,
  r_n_118__20_,r_n_118__19_,r_n_118__18_,r_n_118__17_,r_n_118__16_,r_n_118__15_,
  r_n_118__14_,r_n_118__13_,r_n_118__12_,r_n_118__11_,r_n_118__10_,r_n_118__9_,r_n_118__8_,
  r_n_118__7_,r_n_118__6_,r_n_118__5_,r_n_118__4_,r_n_118__3_,r_n_118__2_,
  r_n_118__1_,r_n_118__0_,r_n_117__63_,r_n_117__62_,r_n_117__61_,r_n_117__60_,
  r_n_117__59_,r_n_117__58_,r_n_117__57_,r_n_117__56_,r_n_117__55_,r_n_117__54_,r_n_117__53_,
  r_n_117__52_,r_n_117__51_,r_n_117__50_,r_n_117__49_,r_n_117__48_,r_n_117__47_,
  r_n_117__46_,r_n_117__45_,r_n_117__44_,r_n_117__43_,r_n_117__42_,r_n_117__41_,
  r_n_117__40_,r_n_117__39_,r_n_117__38_,r_n_117__37_,r_n_117__36_,r_n_117__35_,
  r_n_117__34_,r_n_117__33_,r_n_117__32_,r_n_117__31_,r_n_117__30_,r_n_117__29_,
  r_n_117__28_,r_n_117__27_,r_n_117__26_,r_n_117__25_,r_n_117__24_,r_n_117__23_,
  r_n_117__22_,r_n_117__21_,r_n_117__20_,r_n_117__19_,r_n_117__18_,r_n_117__17_,r_n_117__16_,
  r_n_117__15_,r_n_117__14_,r_n_117__13_,r_n_117__12_,r_n_117__11_,r_n_117__10_,
  r_n_117__9_,r_n_117__8_,r_n_117__7_,r_n_117__6_,r_n_117__5_,r_n_117__4_,
  r_n_117__3_,r_n_117__2_,r_n_117__1_,r_n_117__0_,r_n_116__63_,r_n_116__62_,r_n_116__61_,
  r_n_116__60_,r_n_116__59_,r_n_116__58_,r_n_116__57_,r_n_116__56_,r_n_116__55_,
  r_n_116__54_,r_n_116__53_,r_n_116__52_,r_n_116__51_,r_n_116__50_,r_n_116__49_,
  r_n_116__48_,r_n_116__47_,r_n_116__46_,r_n_116__45_,r_n_116__44_,r_n_116__43_,
  r_n_116__42_,r_n_116__41_,r_n_116__40_,r_n_116__39_,r_n_116__38_,r_n_116__37_,
  r_n_116__36_,r_n_116__35_,r_n_116__34_,r_n_116__33_,r_n_116__32_,r_n_116__31_,r_n_116__30_,
  r_n_116__29_,r_n_116__28_,r_n_116__27_,r_n_116__26_,r_n_116__25_,r_n_116__24_,
  r_n_116__23_,r_n_116__22_,r_n_116__21_,r_n_116__20_,r_n_116__19_,r_n_116__18_,
  r_n_116__17_,r_n_116__16_,r_n_116__15_,r_n_116__14_,r_n_116__13_,r_n_116__12_,
  r_n_116__11_,r_n_116__10_,r_n_116__9_,r_n_116__8_,r_n_116__7_,r_n_116__6_,r_n_116__5_,
  r_n_116__4_,r_n_116__3_,r_n_116__2_,r_n_116__1_,r_n_116__0_,r_n_115__63_,
  r_n_115__62_,r_n_115__61_,r_n_115__60_,r_n_115__59_,r_n_115__58_,r_n_115__57_,
  r_n_115__56_,r_n_115__55_,r_n_115__54_,r_n_115__53_,r_n_115__52_,r_n_115__51_,
  r_n_115__50_,r_n_115__49_,r_n_115__48_,r_n_115__47_,r_n_115__46_,r_n_115__45_,r_n_115__44_,
  r_n_115__43_,r_n_115__42_,r_n_115__41_,r_n_115__40_,r_n_115__39_,r_n_115__38_,
  r_n_115__37_,r_n_115__36_,r_n_115__35_,r_n_115__34_,r_n_115__33_,r_n_115__32_,
  r_n_115__31_,r_n_115__30_,r_n_115__29_,r_n_115__28_,r_n_115__27_,r_n_115__26_,
  r_n_115__25_,r_n_115__24_,r_n_115__23_,r_n_115__22_,r_n_115__21_,r_n_115__20_,
  r_n_115__19_,r_n_115__18_,r_n_115__17_,r_n_115__16_,r_n_115__15_,r_n_115__14_,
  r_n_115__13_,r_n_115__12_,r_n_115__11_,r_n_115__10_,r_n_115__9_,r_n_115__8_,r_n_115__7_,
  r_n_115__6_,r_n_115__5_,r_n_115__4_,r_n_115__3_,r_n_115__2_,r_n_115__1_,
  r_n_115__0_,r_n_114__63_,r_n_114__62_,r_n_114__61_,r_n_114__60_,r_n_114__59_,r_n_114__58_,
  r_n_114__57_,r_n_114__56_,r_n_114__55_,r_n_114__54_,r_n_114__53_,r_n_114__52_,
  r_n_114__51_,r_n_114__50_,r_n_114__49_,r_n_114__48_,r_n_114__47_,r_n_114__46_,
  r_n_114__45_,r_n_114__44_,r_n_114__43_,r_n_114__42_,r_n_114__41_,r_n_114__40_,
  r_n_114__39_,r_n_114__38_,r_n_114__37_,r_n_114__36_,r_n_114__35_,r_n_114__34_,
  r_n_114__33_,r_n_114__32_,r_n_114__31_,r_n_114__30_,r_n_114__29_,r_n_114__28_,
  r_n_114__27_,r_n_114__26_,r_n_114__25_,r_n_114__24_,r_n_114__23_,r_n_114__22_,
  r_n_114__21_,r_n_114__20_,r_n_114__19_,r_n_114__18_,r_n_114__17_,r_n_114__16_,r_n_114__15_,
  r_n_114__14_,r_n_114__13_,r_n_114__12_,r_n_114__11_,r_n_114__10_,r_n_114__9_,
  r_n_114__8_,r_n_114__7_,r_n_114__6_,r_n_114__5_,r_n_114__4_,r_n_114__3_,r_n_114__2_,
  r_n_114__1_,r_n_114__0_,r_n_113__63_,r_n_113__62_,r_n_113__61_,r_n_113__60_,
  r_n_113__59_,r_n_113__58_,r_n_113__57_,r_n_113__56_,r_n_113__55_,r_n_113__54_,
  r_n_113__53_,r_n_113__52_,r_n_113__51_,r_n_113__50_,r_n_113__49_,r_n_113__48_,
  r_n_113__47_,r_n_113__46_,r_n_113__45_,r_n_113__44_,r_n_113__43_,r_n_113__42_,
  r_n_113__41_,r_n_113__40_,r_n_113__39_,r_n_113__38_,r_n_113__37_,r_n_113__36_,
  r_n_113__35_,r_n_113__34_,r_n_113__33_,r_n_113__32_,r_n_113__31_,r_n_113__30_,r_n_113__29_,
  r_n_113__28_,r_n_113__27_,r_n_113__26_,r_n_113__25_,r_n_113__24_,r_n_113__23_,
  r_n_113__22_,r_n_113__21_,r_n_113__20_,r_n_113__19_,r_n_113__18_,r_n_113__17_,
  r_n_113__16_,r_n_113__15_,r_n_113__14_,r_n_113__13_,r_n_113__12_,r_n_113__11_,
  r_n_113__10_,r_n_113__9_,r_n_113__8_,r_n_113__7_,r_n_113__6_,r_n_113__5_,r_n_113__4_,
  r_n_113__3_,r_n_113__2_,r_n_113__1_,r_n_113__0_,r_n_128__63_,r_n_128__62_,
  r_n_128__61_,r_n_128__60_,r_n_128__59_,r_n_128__58_,r_n_128__57_,r_n_128__56_,
  r_n_128__55_,r_n_128__54_,r_n_128__53_,r_n_128__52_,r_n_128__51_,r_n_128__50_,
  r_n_128__49_,r_n_128__48_,r_n_128__47_,r_n_128__46_,r_n_128__45_,r_n_128__44_,r_n_128__43_,
  r_n_128__42_,r_n_128__41_,r_n_128__40_,r_n_128__39_,r_n_128__38_,r_n_128__37_,
  r_n_128__36_,r_n_128__35_,r_n_128__34_,r_n_128__33_,r_n_128__32_,r_n_128__31_,
  r_n_128__30_,r_n_128__29_,r_n_128__28_,r_n_128__27_,r_n_128__26_,r_n_128__25_,
  r_n_128__24_,r_n_128__23_,r_n_128__22_,r_n_128__21_,r_n_128__20_,r_n_128__19_,
  r_n_128__18_,r_n_128__17_,r_n_128__16_,r_n_128__15_,r_n_128__14_,r_n_128__13_,
  r_n_128__12_,r_n_128__11_,r_n_128__10_,r_n_128__9_,r_n_128__8_,r_n_128__7_,r_n_128__6_,
  r_n_128__5_,r_n_128__4_,r_n_128__3_,r_n_128__2_,r_n_128__1_,r_n_128__0_,
  r_n_127__63_,r_n_127__62_,r_n_127__61_,r_n_127__60_,r_n_127__59_,r_n_127__58_,r_n_127__57_,
  r_n_127__56_,r_n_127__55_,r_n_127__54_,r_n_127__53_,r_n_127__52_,r_n_127__51_,
  r_n_127__50_,r_n_127__49_,r_n_127__48_,r_n_127__47_,r_n_127__46_,r_n_127__45_,
  r_n_127__44_,r_n_127__43_,r_n_127__42_,r_n_127__41_,r_n_127__40_,r_n_127__39_,
  r_n_127__38_,r_n_127__37_,r_n_127__36_,r_n_127__35_,r_n_127__34_,r_n_127__33_,
  r_n_127__32_,r_n_127__31_,r_n_127__30_,r_n_127__29_,r_n_127__28_,r_n_127__27_,
  r_n_127__26_,r_n_127__25_,r_n_127__24_,r_n_127__23_,r_n_127__22_,r_n_127__21_,r_n_127__20_,
  r_n_127__19_,r_n_127__18_,r_n_127__17_,r_n_127__16_,r_n_127__15_,r_n_127__14_,
  r_n_127__13_,r_n_127__12_,r_n_127__11_,r_n_127__10_,r_n_127__9_,r_n_127__8_,
  r_n_127__7_,r_n_127__6_,r_n_127__5_,r_n_127__4_,r_n_127__3_,r_n_127__2_,r_n_127__1_,
  r_n_127__0_,r_n_126__63_,r_n_126__62_,r_n_126__61_,r_n_126__60_,r_n_126__59_,
  r_n_126__58_,r_n_126__57_,r_n_126__56_,r_n_126__55_,r_n_126__54_,r_n_126__53_,
  r_n_126__52_,r_n_126__51_,r_n_126__50_,r_n_126__49_,r_n_126__48_,r_n_126__47_,
  r_n_126__46_,r_n_126__45_,r_n_126__44_,r_n_126__43_,r_n_126__42_,r_n_126__41_,
  r_n_126__40_,r_n_126__39_,r_n_126__38_,r_n_126__37_,r_n_126__36_,r_n_126__35_,r_n_126__34_,
  r_n_126__33_,r_n_126__32_,r_n_126__31_,r_n_126__30_,r_n_126__29_,r_n_126__28_,
  r_n_126__27_,r_n_126__26_,r_n_126__25_,r_n_126__24_,r_n_126__23_,r_n_126__22_,
  r_n_126__21_,r_n_126__20_,r_n_126__19_,r_n_126__18_,r_n_126__17_,r_n_126__16_,
  r_n_126__15_,r_n_126__14_,r_n_126__13_,r_n_126__12_,r_n_126__11_,r_n_126__10_,
  r_n_126__9_,r_n_126__8_,r_n_126__7_,r_n_126__6_,r_n_126__5_,r_n_126__4_,r_n_126__3_,
  r_n_126__2_,r_n_126__1_,r_n_126__0_,r_n_125__63_,r_n_125__62_,r_n_125__61_,
  r_n_125__60_,r_n_125__59_,r_n_125__58_,r_n_125__57_,r_n_125__56_,r_n_125__55_,
  r_n_125__54_,r_n_125__53_,r_n_125__52_,r_n_125__51_,r_n_125__50_,r_n_125__49_,r_n_125__48_,
  r_n_125__47_,r_n_125__46_,r_n_125__45_,r_n_125__44_,r_n_125__43_,r_n_125__42_,
  r_n_125__41_,r_n_125__40_,r_n_125__39_,r_n_125__38_,r_n_125__37_,r_n_125__36_,
  r_n_125__35_,r_n_125__34_,r_n_125__33_,r_n_125__32_,r_n_125__31_,r_n_125__30_,
  r_n_125__29_,r_n_125__28_,r_n_125__27_,r_n_125__26_,r_n_125__25_,r_n_125__24_,
  r_n_125__23_,r_n_125__22_,r_n_125__21_,r_n_125__20_,r_n_125__19_,r_n_125__18_,
  r_n_125__17_,r_n_125__16_,r_n_125__15_,r_n_125__14_,r_n_125__13_,r_n_125__12_,
  r_n_125__11_,r_n_125__10_,r_n_125__9_,r_n_125__8_,r_n_125__7_,r_n_125__6_,r_n_125__5_,
  r_n_125__4_,r_n_125__3_,r_n_125__2_,r_n_125__1_,r_n_125__0_,r_n_124__63_,r_n_124__62_,
  r_n_124__61_,r_n_124__60_,r_n_124__59_,r_n_124__58_,r_n_124__57_,r_n_124__56_,
  r_n_124__55_,r_n_124__54_,r_n_124__53_,r_n_124__52_,r_n_124__51_,r_n_124__50_,
  r_n_124__49_,r_n_124__48_,r_n_124__47_,r_n_124__46_,r_n_124__45_,r_n_124__44_,
  r_n_124__43_,r_n_124__42_,r_n_124__41_,r_n_124__40_,r_n_124__39_,r_n_124__38_,
  r_n_124__37_,r_n_124__36_,r_n_124__35_,r_n_124__34_,r_n_124__33_,r_n_124__32_,
  r_n_124__31_,r_n_124__30_,r_n_124__29_,r_n_124__28_,r_n_124__27_,r_n_124__26_,
  r_n_124__25_,r_n_124__24_,r_n_124__23_,r_n_124__22_,r_n_124__21_,r_n_124__20_,r_n_124__19_,
  r_n_124__18_,r_n_124__17_,r_n_124__16_,r_n_124__15_,r_n_124__14_,r_n_124__13_,
  r_n_124__12_,r_n_124__11_,r_n_124__10_,r_n_124__9_,r_n_124__8_,r_n_124__7_,
  r_n_124__6_,r_n_124__5_,r_n_124__4_,r_n_124__3_,r_n_124__2_,r_n_124__1_,r_n_124__0_,
  r_n_123__63_,r_n_123__62_,r_n_123__61_,r_n_123__60_,r_n_123__59_,r_n_123__58_,
  r_n_123__57_,r_n_123__56_,r_n_123__55_,r_n_123__54_,r_n_123__53_,r_n_123__52_,
  r_n_123__51_,r_n_123__50_,r_n_123__49_,r_n_123__48_,r_n_123__47_,r_n_123__46_,
  r_n_123__45_,r_n_123__44_,r_n_123__43_,r_n_123__42_,r_n_123__41_,r_n_123__40_,
  r_n_123__39_,r_n_123__38_,r_n_123__37_,r_n_123__36_,r_n_123__35_,r_n_123__34_,r_n_123__33_,
  r_n_123__32_,r_n_123__31_,r_n_123__30_,r_n_123__29_,r_n_123__28_,r_n_123__27_,
  r_n_123__26_,r_n_123__25_,r_n_123__24_,r_n_123__23_,r_n_123__22_,r_n_123__21_,
  r_n_123__20_,r_n_123__19_,r_n_123__18_,r_n_123__17_,r_n_123__16_,r_n_123__15_,
  r_n_123__14_,r_n_123__13_,r_n_123__12_,r_n_123__11_,r_n_123__10_,r_n_123__9_,
  r_n_123__8_,r_n_123__7_,r_n_123__6_,r_n_123__5_,r_n_123__4_,r_n_123__3_,r_n_123__2_,
  r_n_123__1_,r_n_123__0_,r_n_122__63_,r_n_122__62_,r_n_122__61_,r_n_122__60_,
  r_n_122__59_,r_n_122__58_,r_n_122__57_,r_n_122__56_,r_n_122__55_,r_n_122__54_,
  r_n_122__53_,r_n_122__52_,r_n_122__51_,r_n_122__50_,r_n_122__49_,r_n_122__48_,r_n_122__47_,
  r_n_122__46_,r_n_122__45_,r_n_122__44_,r_n_122__43_,r_n_122__42_,r_n_122__41_,
  r_n_122__40_,r_n_122__39_,r_n_122__38_,r_n_122__37_,r_n_122__36_,r_n_122__35_,
  r_n_122__34_,r_n_122__33_,r_n_122__32_,r_n_122__31_,r_n_122__30_,r_n_122__29_,
  r_n_122__28_,r_n_122__27_,r_n_122__26_,r_n_122__25_,r_n_122__24_,r_n_122__23_,
  r_n_122__22_,r_n_122__21_,r_n_122__20_,r_n_122__19_,r_n_122__18_,r_n_122__17_,
  r_n_122__16_,r_n_122__15_,r_n_122__14_,r_n_122__13_,r_n_122__12_,r_n_122__11_,r_n_122__10_,
  r_n_122__9_,r_n_122__8_,r_n_122__7_,r_n_122__6_,r_n_122__5_,r_n_122__4_,
  r_n_122__3_,r_n_122__2_,r_n_122__1_,r_n_122__0_,r_n_121__63_,r_n_121__62_,r_n_121__61_,
  r_n_121__60_,r_n_121__59_,r_n_121__58_,r_n_121__57_,r_n_121__56_,r_n_121__55_,
  r_n_121__54_,r_n_121__53_,r_n_121__52_,r_n_121__51_,r_n_121__50_,r_n_121__49_,
  r_n_121__48_,r_n_121__47_,r_n_121__46_,r_n_121__45_,r_n_121__44_,r_n_121__43_,
  r_n_121__42_,r_n_121__41_,r_n_121__40_,r_n_121__39_,r_n_121__38_,r_n_121__37_,
  r_n_121__36_,r_n_121__35_,r_n_121__34_,r_n_121__33_,r_n_121__32_,r_n_121__31_,
  r_n_121__30_,r_n_121__29_,r_n_121__28_,r_n_121__27_,r_n_121__26_,r_n_121__25_,r_n_121__24_,
  r_n_121__23_,r_n_121__22_,r_n_121__21_,r_n_121__20_,r_n_121__19_,r_n_121__18_,
  r_n_121__17_,r_n_121__16_,r_n_121__15_,r_n_121__14_,r_n_121__13_,r_n_121__12_,
  r_n_121__11_,r_n_121__10_,r_n_121__9_,r_n_121__8_,r_n_121__7_,r_n_121__6_,
  r_n_121__5_,r_n_121__4_,r_n_121__3_,r_n_121__2_,r_n_121__1_,r_n_121__0_,r_n_136__63_,
  r_n_136__62_,r_n_136__61_,r_n_136__60_,r_n_136__59_,r_n_136__58_,r_n_136__57_,
  r_n_136__56_,r_n_136__55_,r_n_136__54_,r_n_136__53_,r_n_136__52_,r_n_136__51_,
  r_n_136__50_,r_n_136__49_,r_n_136__48_,r_n_136__47_,r_n_136__46_,r_n_136__45_,
  r_n_136__44_,r_n_136__43_,r_n_136__42_,r_n_136__41_,r_n_136__40_,r_n_136__39_,r_n_136__38_,
  r_n_136__37_,r_n_136__36_,r_n_136__35_,r_n_136__34_,r_n_136__33_,r_n_136__32_,
  r_n_136__31_,r_n_136__30_,r_n_136__29_,r_n_136__28_,r_n_136__27_,r_n_136__26_,
  r_n_136__25_,r_n_136__24_,r_n_136__23_,r_n_136__22_,r_n_136__21_,r_n_136__20_,
  r_n_136__19_,r_n_136__18_,r_n_136__17_,r_n_136__16_,r_n_136__15_,r_n_136__14_,
  r_n_136__13_,r_n_136__12_,r_n_136__11_,r_n_136__10_,r_n_136__9_,r_n_136__8_,r_n_136__7_,
  r_n_136__6_,r_n_136__5_,r_n_136__4_,r_n_136__3_,r_n_136__2_,r_n_136__1_,
  r_n_136__0_,r_n_135__63_,r_n_135__62_,r_n_135__61_,r_n_135__60_,r_n_135__59_,
  r_n_135__58_,r_n_135__57_,r_n_135__56_,r_n_135__55_,r_n_135__54_,r_n_135__53_,r_n_135__52_,
  r_n_135__51_,r_n_135__50_,r_n_135__49_,r_n_135__48_,r_n_135__47_,r_n_135__46_,
  r_n_135__45_,r_n_135__44_,r_n_135__43_,r_n_135__42_,r_n_135__41_,r_n_135__40_,
  r_n_135__39_,r_n_135__38_,r_n_135__37_,r_n_135__36_,r_n_135__35_,r_n_135__34_,
  r_n_135__33_,r_n_135__32_,r_n_135__31_,r_n_135__30_,r_n_135__29_,r_n_135__28_,
  r_n_135__27_,r_n_135__26_,r_n_135__25_,r_n_135__24_,r_n_135__23_,r_n_135__22_,
  r_n_135__21_,r_n_135__20_,r_n_135__19_,r_n_135__18_,r_n_135__17_,r_n_135__16_,
  r_n_135__15_,r_n_135__14_,r_n_135__13_,r_n_135__12_,r_n_135__11_,r_n_135__10_,r_n_135__9_,
  r_n_135__8_,r_n_135__7_,r_n_135__6_,r_n_135__5_,r_n_135__4_,r_n_135__3_,
  r_n_135__2_,r_n_135__1_,r_n_135__0_,r_n_134__63_,r_n_134__62_,r_n_134__61_,r_n_134__60_,
  r_n_134__59_,r_n_134__58_,r_n_134__57_,r_n_134__56_,r_n_134__55_,r_n_134__54_,
  r_n_134__53_,r_n_134__52_,r_n_134__51_,r_n_134__50_,r_n_134__49_,r_n_134__48_,
  r_n_134__47_,r_n_134__46_,r_n_134__45_,r_n_134__44_,r_n_134__43_,r_n_134__42_,
  r_n_134__41_,r_n_134__40_,r_n_134__39_,r_n_134__38_,r_n_134__37_,r_n_134__36_,
  r_n_134__35_,r_n_134__34_,r_n_134__33_,r_n_134__32_,r_n_134__31_,r_n_134__30_,
  r_n_134__29_,r_n_134__28_,r_n_134__27_,r_n_134__26_,r_n_134__25_,r_n_134__24_,r_n_134__23_,
  r_n_134__22_,r_n_134__21_,r_n_134__20_,r_n_134__19_,r_n_134__18_,r_n_134__17_,
  r_n_134__16_,r_n_134__15_,r_n_134__14_,r_n_134__13_,r_n_134__12_,r_n_134__11_,
  r_n_134__10_,r_n_134__9_,r_n_134__8_,r_n_134__7_,r_n_134__6_,r_n_134__5_,r_n_134__4_,
  r_n_134__3_,r_n_134__2_,r_n_134__1_,r_n_134__0_,r_n_133__63_,r_n_133__62_,
  r_n_133__61_,r_n_133__60_,r_n_133__59_,r_n_133__58_,r_n_133__57_,r_n_133__56_,
  r_n_133__55_,r_n_133__54_,r_n_133__53_,r_n_133__52_,r_n_133__51_,r_n_133__50_,
  r_n_133__49_,r_n_133__48_,r_n_133__47_,r_n_133__46_,r_n_133__45_,r_n_133__44_,
  r_n_133__43_,r_n_133__42_,r_n_133__41_,r_n_133__40_,r_n_133__39_,r_n_133__38_,r_n_133__37_,
  r_n_133__36_,r_n_133__35_,r_n_133__34_,r_n_133__33_,r_n_133__32_,r_n_133__31_,
  r_n_133__30_,r_n_133__29_,r_n_133__28_,r_n_133__27_,r_n_133__26_,r_n_133__25_,
  r_n_133__24_,r_n_133__23_,r_n_133__22_,r_n_133__21_,r_n_133__20_,r_n_133__19_,
  r_n_133__18_,r_n_133__17_,r_n_133__16_,r_n_133__15_,r_n_133__14_,r_n_133__13_,
  r_n_133__12_,r_n_133__11_,r_n_133__10_,r_n_133__9_,r_n_133__8_,r_n_133__7_,r_n_133__6_,
  r_n_133__5_,r_n_133__4_,r_n_133__3_,r_n_133__2_,r_n_133__1_,r_n_133__0_,
  r_n_132__63_,r_n_132__62_,r_n_132__61_,r_n_132__60_,r_n_132__59_,r_n_132__58_,
  r_n_132__57_,r_n_132__56_,r_n_132__55_,r_n_132__54_,r_n_132__53_,r_n_132__52_,r_n_132__51_,
  r_n_132__50_,r_n_132__49_,r_n_132__48_,r_n_132__47_,r_n_132__46_,r_n_132__45_,
  r_n_132__44_,r_n_132__43_,r_n_132__42_,r_n_132__41_,r_n_132__40_,r_n_132__39_,
  r_n_132__38_,r_n_132__37_,r_n_132__36_,r_n_132__35_,r_n_132__34_,r_n_132__33_,
  r_n_132__32_,r_n_132__31_,r_n_132__30_,r_n_132__29_,r_n_132__28_,r_n_132__27_,
  r_n_132__26_,r_n_132__25_,r_n_132__24_,r_n_132__23_,r_n_132__22_,r_n_132__21_,
  r_n_132__20_,r_n_132__19_,r_n_132__18_,r_n_132__17_,r_n_132__16_,r_n_132__15_,r_n_132__14_,
  r_n_132__13_,r_n_132__12_,r_n_132__11_,r_n_132__10_,r_n_132__9_,r_n_132__8_,
  r_n_132__7_,r_n_132__6_,r_n_132__5_,r_n_132__4_,r_n_132__3_,r_n_132__2_,r_n_132__1_,
  r_n_132__0_,r_n_131__63_,r_n_131__62_,r_n_131__61_,r_n_131__60_,r_n_131__59_,
  r_n_131__58_,r_n_131__57_,r_n_131__56_,r_n_131__55_,r_n_131__54_,r_n_131__53_,
  r_n_131__52_,r_n_131__51_,r_n_131__50_,r_n_131__49_,r_n_131__48_,r_n_131__47_,
  r_n_131__46_,r_n_131__45_,r_n_131__44_,r_n_131__43_,r_n_131__42_,r_n_131__41_,
  r_n_131__40_,r_n_131__39_,r_n_131__38_,r_n_131__37_,r_n_131__36_,r_n_131__35_,
  r_n_131__34_,r_n_131__33_,r_n_131__32_,r_n_131__31_,r_n_131__30_,r_n_131__29_,r_n_131__28_,
  r_n_131__27_,r_n_131__26_,r_n_131__25_,r_n_131__24_,r_n_131__23_,r_n_131__22_,
  r_n_131__21_,r_n_131__20_,r_n_131__19_,r_n_131__18_,r_n_131__17_,r_n_131__16_,
  r_n_131__15_,r_n_131__14_,r_n_131__13_,r_n_131__12_,r_n_131__11_,r_n_131__10_,
  r_n_131__9_,r_n_131__8_,r_n_131__7_,r_n_131__6_,r_n_131__5_,r_n_131__4_,r_n_131__3_,
  r_n_131__2_,r_n_131__1_,r_n_131__0_,r_n_130__63_,r_n_130__62_,r_n_130__61_,
  r_n_130__60_,r_n_130__59_,r_n_130__58_,r_n_130__57_,r_n_130__56_,r_n_130__55_,
  r_n_130__54_,r_n_130__53_,r_n_130__52_,r_n_130__51_,r_n_130__50_,r_n_130__49_,
  r_n_130__48_,r_n_130__47_,r_n_130__46_,r_n_130__45_,r_n_130__44_,r_n_130__43_,r_n_130__42_,
  r_n_130__41_,r_n_130__40_,r_n_130__39_,r_n_130__38_,r_n_130__37_,r_n_130__36_,
  r_n_130__35_,r_n_130__34_,r_n_130__33_,r_n_130__32_,r_n_130__31_,r_n_130__30_,
  r_n_130__29_,r_n_130__28_,r_n_130__27_,r_n_130__26_,r_n_130__25_,r_n_130__24_,
  r_n_130__23_,r_n_130__22_,r_n_130__21_,r_n_130__20_,r_n_130__19_,r_n_130__18_,
  r_n_130__17_,r_n_130__16_,r_n_130__15_,r_n_130__14_,r_n_130__13_,r_n_130__12_,
  r_n_130__11_,r_n_130__10_,r_n_130__9_,r_n_130__8_,r_n_130__7_,r_n_130__6_,r_n_130__5_,
  r_n_130__4_,r_n_130__3_,r_n_130__2_,r_n_130__1_,r_n_130__0_,r_n_129__63_,
  r_n_129__62_,r_n_129__61_,r_n_129__60_,r_n_129__59_,r_n_129__58_,r_n_129__57_,r_n_129__56_,
  r_n_129__55_,r_n_129__54_,r_n_129__53_,r_n_129__52_,r_n_129__51_,r_n_129__50_,
  r_n_129__49_,r_n_129__48_,r_n_129__47_,r_n_129__46_,r_n_129__45_,r_n_129__44_,
  r_n_129__43_,r_n_129__42_,r_n_129__41_,r_n_129__40_,r_n_129__39_,r_n_129__38_,
  r_n_129__37_,r_n_129__36_,r_n_129__35_,r_n_129__34_,r_n_129__33_,r_n_129__32_,
  r_n_129__31_,r_n_129__30_,r_n_129__29_,r_n_129__28_,r_n_129__27_,r_n_129__26_,
  r_n_129__25_,r_n_129__24_,r_n_129__23_,r_n_129__22_,r_n_129__21_,r_n_129__20_,
  r_n_129__19_,r_n_129__18_,r_n_129__17_,r_n_129__16_,r_n_129__15_,r_n_129__14_,r_n_129__13_,
  r_n_129__12_,r_n_129__11_,r_n_129__10_,r_n_129__9_,r_n_129__8_,r_n_129__7_,
  r_n_129__6_,r_n_129__5_,r_n_129__4_,r_n_129__3_,r_n_129__2_,r_n_129__1_,r_n_129__0_,
  r_n_144__63_,r_n_144__62_,r_n_144__61_,r_n_144__60_,r_n_144__59_,r_n_144__58_,
  r_n_144__57_,r_n_144__56_,r_n_144__55_,r_n_144__54_,r_n_144__53_,r_n_144__52_,
  r_n_144__51_,r_n_144__50_,r_n_144__49_,r_n_144__48_,r_n_144__47_,r_n_144__46_,
  r_n_144__45_,r_n_144__44_,r_n_144__43_,r_n_144__42_,r_n_144__41_,r_n_144__40_,
  r_n_144__39_,r_n_144__38_,r_n_144__37_,r_n_144__36_,r_n_144__35_,r_n_144__34_,
  r_n_144__33_,r_n_144__32_,r_n_144__31_,r_n_144__30_,r_n_144__29_,r_n_144__28_,r_n_144__27_,
  r_n_144__26_,r_n_144__25_,r_n_144__24_,r_n_144__23_,r_n_144__22_,r_n_144__21_,
  r_n_144__20_,r_n_144__19_,r_n_144__18_,r_n_144__17_,r_n_144__16_,r_n_144__15_,
  r_n_144__14_,r_n_144__13_,r_n_144__12_,r_n_144__11_,r_n_144__10_,r_n_144__9_,
  r_n_144__8_,r_n_144__7_,r_n_144__6_,r_n_144__5_,r_n_144__4_,r_n_144__3_,r_n_144__2_,
  r_n_144__1_,r_n_144__0_,r_n_143__63_,r_n_143__62_,r_n_143__61_,r_n_143__60_,
  r_n_143__59_,r_n_143__58_,r_n_143__57_,r_n_143__56_,r_n_143__55_,r_n_143__54_,
  r_n_143__53_,r_n_143__52_,r_n_143__51_,r_n_143__50_,r_n_143__49_,r_n_143__48_,
  r_n_143__47_,r_n_143__46_,r_n_143__45_,r_n_143__44_,r_n_143__43_,r_n_143__42_,r_n_143__41_,
  r_n_143__40_,r_n_143__39_,r_n_143__38_,r_n_143__37_,r_n_143__36_,r_n_143__35_,
  r_n_143__34_,r_n_143__33_,r_n_143__32_,r_n_143__31_,r_n_143__30_,r_n_143__29_,
  r_n_143__28_,r_n_143__27_,r_n_143__26_,r_n_143__25_,r_n_143__24_,r_n_143__23_,
  r_n_143__22_,r_n_143__21_,r_n_143__20_,r_n_143__19_,r_n_143__18_,r_n_143__17_,
  r_n_143__16_,r_n_143__15_,r_n_143__14_,r_n_143__13_,r_n_143__12_,r_n_143__11_,
  r_n_143__10_,r_n_143__9_,r_n_143__8_,r_n_143__7_,r_n_143__6_,r_n_143__5_,r_n_143__4_,
  r_n_143__3_,r_n_143__2_,r_n_143__1_,r_n_143__0_,r_n_142__63_,r_n_142__62_,
  r_n_142__61_,r_n_142__60_,r_n_142__59_,r_n_142__58_,r_n_142__57_,r_n_142__56_,r_n_142__55_,
  r_n_142__54_,r_n_142__53_,r_n_142__52_,r_n_142__51_,r_n_142__50_,r_n_142__49_,
  r_n_142__48_,r_n_142__47_,r_n_142__46_,r_n_142__45_,r_n_142__44_,r_n_142__43_,
  r_n_142__42_,r_n_142__41_,r_n_142__40_,r_n_142__39_,r_n_142__38_,r_n_142__37_,
  r_n_142__36_,r_n_142__35_,r_n_142__34_,r_n_142__33_,r_n_142__32_,r_n_142__31_,
  r_n_142__30_,r_n_142__29_,r_n_142__28_,r_n_142__27_,r_n_142__26_,r_n_142__25_,
  r_n_142__24_,r_n_142__23_,r_n_142__22_,r_n_142__21_,r_n_142__20_,r_n_142__19_,r_n_142__18_,
  r_n_142__17_,r_n_142__16_,r_n_142__15_,r_n_142__14_,r_n_142__13_,r_n_142__12_,
  r_n_142__11_,r_n_142__10_,r_n_142__9_,r_n_142__8_,r_n_142__7_,r_n_142__6_,
  r_n_142__5_,r_n_142__4_,r_n_142__3_,r_n_142__2_,r_n_142__1_,r_n_142__0_,r_n_141__63_,
  r_n_141__62_,r_n_141__61_,r_n_141__60_,r_n_141__59_,r_n_141__58_,r_n_141__57_,
  r_n_141__56_,r_n_141__55_,r_n_141__54_,r_n_141__53_,r_n_141__52_,r_n_141__51_,
  r_n_141__50_,r_n_141__49_,r_n_141__48_,r_n_141__47_,r_n_141__46_,r_n_141__45_,
  r_n_141__44_,r_n_141__43_,r_n_141__42_,r_n_141__41_,r_n_141__40_,r_n_141__39_,
  r_n_141__38_,r_n_141__37_,r_n_141__36_,r_n_141__35_,r_n_141__34_,r_n_141__33_,r_n_141__32_,
  r_n_141__31_,r_n_141__30_,r_n_141__29_,r_n_141__28_,r_n_141__27_,r_n_141__26_,
  r_n_141__25_,r_n_141__24_,r_n_141__23_,r_n_141__22_,r_n_141__21_,r_n_141__20_,
  r_n_141__19_,r_n_141__18_,r_n_141__17_,r_n_141__16_,r_n_141__15_,r_n_141__14_,
  r_n_141__13_,r_n_141__12_,r_n_141__11_,r_n_141__10_,r_n_141__9_,r_n_141__8_,
  r_n_141__7_,r_n_141__6_,r_n_141__5_,r_n_141__4_,r_n_141__3_,r_n_141__2_,r_n_141__1_,
  r_n_141__0_,r_n_140__63_,r_n_140__62_,r_n_140__61_,r_n_140__60_,r_n_140__59_,
  r_n_140__58_,r_n_140__57_,r_n_140__56_,r_n_140__55_,r_n_140__54_,r_n_140__53_,
  r_n_140__52_,r_n_140__51_,r_n_140__50_,r_n_140__49_,r_n_140__48_,r_n_140__47_,r_n_140__46_,
  r_n_140__45_,r_n_140__44_,r_n_140__43_,r_n_140__42_,r_n_140__41_,r_n_140__40_,
  r_n_140__39_,r_n_140__38_,r_n_140__37_,r_n_140__36_,r_n_140__35_,r_n_140__34_,
  r_n_140__33_,r_n_140__32_,r_n_140__31_,r_n_140__30_,r_n_140__29_,r_n_140__28_,
  r_n_140__27_,r_n_140__26_,r_n_140__25_,r_n_140__24_,r_n_140__23_,r_n_140__22_,
  r_n_140__21_,r_n_140__20_,r_n_140__19_,r_n_140__18_,r_n_140__17_,r_n_140__16_,
  r_n_140__15_,r_n_140__14_,r_n_140__13_,r_n_140__12_,r_n_140__11_,r_n_140__10_,r_n_140__9_,
  r_n_140__8_,r_n_140__7_,r_n_140__6_,r_n_140__5_,r_n_140__4_,r_n_140__3_,
  r_n_140__2_,r_n_140__1_,r_n_140__0_,r_n_139__63_,r_n_139__62_,r_n_139__61_,r_n_139__60_,
  r_n_139__59_,r_n_139__58_,r_n_139__57_,r_n_139__56_,r_n_139__55_,r_n_139__54_,
  r_n_139__53_,r_n_139__52_,r_n_139__51_,r_n_139__50_,r_n_139__49_,r_n_139__48_,
  r_n_139__47_,r_n_139__46_,r_n_139__45_,r_n_139__44_,r_n_139__43_,r_n_139__42_,
  r_n_139__41_,r_n_139__40_,r_n_139__39_,r_n_139__38_,r_n_139__37_,r_n_139__36_,
  r_n_139__35_,r_n_139__34_,r_n_139__33_,r_n_139__32_,r_n_139__31_,r_n_139__30_,
  r_n_139__29_,r_n_139__28_,r_n_139__27_,r_n_139__26_,r_n_139__25_,r_n_139__24_,
  r_n_139__23_,r_n_139__22_,r_n_139__21_,r_n_139__20_,r_n_139__19_,r_n_139__18_,r_n_139__17_,
  r_n_139__16_,r_n_139__15_,r_n_139__14_,r_n_139__13_,r_n_139__12_,r_n_139__11_,
  r_n_139__10_,r_n_139__9_,r_n_139__8_,r_n_139__7_,r_n_139__6_,r_n_139__5_,
  r_n_139__4_,r_n_139__3_,r_n_139__2_,r_n_139__1_,r_n_139__0_,r_n_138__63_,r_n_138__62_,
  r_n_138__61_,r_n_138__60_,r_n_138__59_,r_n_138__58_,r_n_138__57_,r_n_138__56_,
  r_n_138__55_,r_n_138__54_,r_n_138__53_,r_n_138__52_,r_n_138__51_,r_n_138__50_,
  r_n_138__49_,r_n_138__48_,r_n_138__47_,r_n_138__46_,r_n_138__45_,r_n_138__44_,
  r_n_138__43_,r_n_138__42_,r_n_138__41_,r_n_138__40_,r_n_138__39_,r_n_138__38_,
  r_n_138__37_,r_n_138__36_,r_n_138__35_,r_n_138__34_,r_n_138__33_,r_n_138__32_,r_n_138__31_,
  r_n_138__30_,r_n_138__29_,r_n_138__28_,r_n_138__27_,r_n_138__26_,r_n_138__25_,
  r_n_138__24_,r_n_138__23_,r_n_138__22_,r_n_138__21_,r_n_138__20_,r_n_138__19_,
  r_n_138__18_,r_n_138__17_,r_n_138__16_,r_n_138__15_,r_n_138__14_,r_n_138__13_,
  r_n_138__12_,r_n_138__11_,r_n_138__10_,r_n_138__9_,r_n_138__8_,r_n_138__7_,r_n_138__6_,
  r_n_138__5_,r_n_138__4_,r_n_138__3_,r_n_138__2_,r_n_138__1_,r_n_138__0_,
  r_n_137__63_,r_n_137__62_,r_n_137__61_,r_n_137__60_,r_n_137__59_,r_n_137__58_,
  r_n_137__57_,r_n_137__56_,r_n_137__55_,r_n_137__54_,r_n_137__53_,r_n_137__52_,
  r_n_137__51_,r_n_137__50_,r_n_137__49_,r_n_137__48_,r_n_137__47_,r_n_137__46_,r_n_137__45_,
  r_n_137__44_,r_n_137__43_,r_n_137__42_,r_n_137__41_,r_n_137__40_,r_n_137__39_,
  r_n_137__38_,r_n_137__37_,r_n_137__36_,r_n_137__35_,r_n_137__34_,r_n_137__33_,
  r_n_137__32_,r_n_137__31_,r_n_137__30_,r_n_137__29_,r_n_137__28_,r_n_137__27_,
  r_n_137__26_,r_n_137__25_,r_n_137__24_,r_n_137__23_,r_n_137__22_,r_n_137__21_,
  r_n_137__20_,r_n_137__19_,r_n_137__18_,r_n_137__17_,r_n_137__16_,r_n_137__15_,
  r_n_137__14_,r_n_137__13_,r_n_137__12_,r_n_137__11_,r_n_137__10_,r_n_137__9_,r_n_137__8_,
  r_n_137__7_,r_n_137__6_,r_n_137__5_,r_n_137__4_,r_n_137__3_,r_n_137__2_,
  r_n_137__1_,r_n_137__0_,r_n_152__63_,r_n_152__62_,r_n_152__61_,r_n_152__60_,r_n_152__59_,
  r_n_152__58_,r_n_152__57_,r_n_152__56_,r_n_152__55_,r_n_152__54_,r_n_152__53_,
  r_n_152__52_,r_n_152__51_,r_n_152__50_,r_n_152__49_,r_n_152__48_,r_n_152__47_,
  r_n_152__46_,r_n_152__45_,r_n_152__44_,r_n_152__43_,r_n_152__42_,r_n_152__41_,
  r_n_152__40_,r_n_152__39_,r_n_152__38_,r_n_152__37_,r_n_152__36_,r_n_152__35_,
  r_n_152__34_,r_n_152__33_,r_n_152__32_,r_n_152__31_,r_n_152__30_,r_n_152__29_,
  r_n_152__28_,r_n_152__27_,r_n_152__26_,r_n_152__25_,r_n_152__24_,r_n_152__23_,r_n_152__22_,
  r_n_152__21_,r_n_152__20_,r_n_152__19_,r_n_152__18_,r_n_152__17_,r_n_152__16_,
  r_n_152__15_,r_n_152__14_,r_n_152__13_,r_n_152__12_,r_n_152__11_,r_n_152__10_,
  r_n_152__9_,r_n_152__8_,r_n_152__7_,r_n_152__6_,r_n_152__5_,r_n_152__4_,r_n_152__3_,
  r_n_152__2_,r_n_152__1_,r_n_152__0_,r_n_151__63_,r_n_151__62_,r_n_151__61_,
  r_n_151__60_,r_n_151__59_,r_n_151__58_,r_n_151__57_,r_n_151__56_,r_n_151__55_,
  r_n_151__54_,r_n_151__53_,r_n_151__52_,r_n_151__51_,r_n_151__50_,r_n_151__49_,
  r_n_151__48_,r_n_151__47_,r_n_151__46_,r_n_151__45_,r_n_151__44_,r_n_151__43_,
  r_n_151__42_,r_n_151__41_,r_n_151__40_,r_n_151__39_,r_n_151__38_,r_n_151__37_,r_n_151__36_,
  r_n_151__35_,r_n_151__34_,r_n_151__33_,r_n_151__32_,r_n_151__31_,r_n_151__30_,
  r_n_151__29_,r_n_151__28_,r_n_151__27_,r_n_151__26_,r_n_151__25_,r_n_151__24_,
  r_n_151__23_,r_n_151__22_,r_n_151__21_,r_n_151__20_,r_n_151__19_,r_n_151__18_,
  r_n_151__17_,r_n_151__16_,r_n_151__15_,r_n_151__14_,r_n_151__13_,r_n_151__12_,
  r_n_151__11_,r_n_151__10_,r_n_151__9_,r_n_151__8_,r_n_151__7_,r_n_151__6_,r_n_151__5_,
  r_n_151__4_,r_n_151__3_,r_n_151__2_,r_n_151__1_,r_n_151__0_,r_n_150__63_,
  r_n_150__62_,r_n_150__61_,r_n_150__60_,r_n_150__59_,r_n_150__58_,r_n_150__57_,
  r_n_150__56_,r_n_150__55_,r_n_150__54_,r_n_150__53_,r_n_150__52_,r_n_150__51_,r_n_150__50_,
  r_n_150__49_,r_n_150__48_,r_n_150__47_,r_n_150__46_,r_n_150__45_,r_n_150__44_,
  r_n_150__43_,r_n_150__42_,r_n_150__41_,r_n_150__40_,r_n_150__39_,r_n_150__38_,
  r_n_150__37_,r_n_150__36_,r_n_150__35_,r_n_150__34_,r_n_150__33_,r_n_150__32_,
  r_n_150__31_,r_n_150__30_,r_n_150__29_,r_n_150__28_,r_n_150__27_,r_n_150__26_,
  r_n_150__25_,r_n_150__24_,r_n_150__23_,r_n_150__22_,r_n_150__21_,r_n_150__20_,
  r_n_150__19_,r_n_150__18_,r_n_150__17_,r_n_150__16_,r_n_150__15_,r_n_150__14_,
  r_n_150__13_,r_n_150__12_,r_n_150__11_,r_n_150__10_,r_n_150__9_,r_n_150__8_,r_n_150__7_,
  r_n_150__6_,r_n_150__5_,r_n_150__4_,r_n_150__3_,r_n_150__2_,r_n_150__1_,r_n_150__0_,
  r_n_149__63_,r_n_149__62_,r_n_149__61_,r_n_149__60_,r_n_149__59_,r_n_149__58_,
  r_n_149__57_,r_n_149__56_,r_n_149__55_,r_n_149__54_,r_n_149__53_,r_n_149__52_,
  r_n_149__51_,r_n_149__50_,r_n_149__49_,r_n_149__48_,r_n_149__47_,r_n_149__46_,
  r_n_149__45_,r_n_149__44_,r_n_149__43_,r_n_149__42_,r_n_149__41_,r_n_149__40_,
  r_n_149__39_,r_n_149__38_,r_n_149__37_,r_n_149__36_,r_n_149__35_,r_n_149__34_,
  r_n_149__33_,r_n_149__32_,r_n_149__31_,r_n_149__30_,r_n_149__29_,r_n_149__28_,
  r_n_149__27_,r_n_149__26_,r_n_149__25_,r_n_149__24_,r_n_149__23_,r_n_149__22_,r_n_149__21_,
  r_n_149__20_,r_n_149__19_,r_n_149__18_,r_n_149__17_,r_n_149__16_,r_n_149__15_,
  r_n_149__14_,r_n_149__13_,r_n_149__12_,r_n_149__11_,r_n_149__10_,r_n_149__9_,
  r_n_149__8_,r_n_149__7_,r_n_149__6_,r_n_149__5_,r_n_149__4_,r_n_149__3_,r_n_149__2_,
  r_n_149__1_,r_n_149__0_,r_n_148__63_,r_n_148__62_,r_n_148__61_,r_n_148__60_,
  r_n_148__59_,r_n_148__58_,r_n_148__57_,r_n_148__56_,r_n_148__55_,r_n_148__54_,
  r_n_148__53_,r_n_148__52_,r_n_148__51_,r_n_148__50_,r_n_148__49_,r_n_148__48_,
  r_n_148__47_,r_n_148__46_,r_n_148__45_,r_n_148__44_,r_n_148__43_,r_n_148__42_,
  r_n_148__41_,r_n_148__40_,r_n_148__39_,r_n_148__38_,r_n_148__37_,r_n_148__36_,r_n_148__35_,
  r_n_148__34_,r_n_148__33_,r_n_148__32_,r_n_148__31_,r_n_148__30_,r_n_148__29_,
  r_n_148__28_,r_n_148__27_,r_n_148__26_,r_n_148__25_,r_n_148__24_,r_n_148__23_,
  r_n_148__22_,r_n_148__21_,r_n_148__20_,r_n_148__19_,r_n_148__18_,r_n_148__17_,
  r_n_148__16_,r_n_148__15_,r_n_148__14_,r_n_148__13_,r_n_148__12_,r_n_148__11_,
  r_n_148__10_,r_n_148__9_,r_n_148__8_,r_n_148__7_,r_n_148__6_,r_n_148__5_,r_n_148__4_,
  r_n_148__3_,r_n_148__2_,r_n_148__1_,r_n_148__0_,r_n_147__63_,r_n_147__62_,
  r_n_147__61_,r_n_147__60_,r_n_147__59_,r_n_147__58_,r_n_147__57_,r_n_147__56_,
  r_n_147__55_,r_n_147__54_,r_n_147__53_,r_n_147__52_,r_n_147__51_,r_n_147__50_,r_n_147__49_,
  r_n_147__48_,r_n_147__47_,r_n_147__46_,r_n_147__45_,r_n_147__44_,r_n_147__43_,
  r_n_147__42_,r_n_147__41_,r_n_147__40_,r_n_147__39_,r_n_147__38_,r_n_147__37_,
  r_n_147__36_,r_n_147__35_,r_n_147__34_,r_n_147__33_,r_n_147__32_,r_n_147__31_,
  r_n_147__30_,r_n_147__29_,r_n_147__28_,r_n_147__27_,r_n_147__26_,r_n_147__25_,
  r_n_147__24_,r_n_147__23_,r_n_147__22_,r_n_147__21_,r_n_147__20_,r_n_147__19_,
  r_n_147__18_,r_n_147__17_,r_n_147__16_,r_n_147__15_,r_n_147__14_,r_n_147__13_,r_n_147__12_,
  r_n_147__11_,r_n_147__10_,r_n_147__9_,r_n_147__8_,r_n_147__7_,r_n_147__6_,
  r_n_147__5_,r_n_147__4_,r_n_147__3_,r_n_147__2_,r_n_147__1_,r_n_147__0_,r_n_146__63_,
  r_n_146__62_,r_n_146__61_,r_n_146__60_,r_n_146__59_,r_n_146__58_,r_n_146__57_,
  r_n_146__56_,r_n_146__55_,r_n_146__54_,r_n_146__53_,r_n_146__52_,r_n_146__51_,
  r_n_146__50_,r_n_146__49_,r_n_146__48_,r_n_146__47_,r_n_146__46_,r_n_146__45_,
  r_n_146__44_,r_n_146__43_,r_n_146__42_,r_n_146__41_,r_n_146__40_,r_n_146__39_,
  r_n_146__38_,r_n_146__37_,r_n_146__36_,r_n_146__35_,r_n_146__34_,r_n_146__33_,
  r_n_146__32_,r_n_146__31_,r_n_146__30_,r_n_146__29_,r_n_146__28_,r_n_146__27_,r_n_146__26_,
  r_n_146__25_,r_n_146__24_,r_n_146__23_,r_n_146__22_,r_n_146__21_,r_n_146__20_,
  r_n_146__19_,r_n_146__18_,r_n_146__17_,r_n_146__16_,r_n_146__15_,r_n_146__14_,
  r_n_146__13_,r_n_146__12_,r_n_146__11_,r_n_146__10_,r_n_146__9_,r_n_146__8_,
  r_n_146__7_,r_n_146__6_,r_n_146__5_,r_n_146__4_,r_n_146__3_,r_n_146__2_,r_n_146__1_,
  r_n_146__0_,r_n_145__63_,r_n_145__62_,r_n_145__61_,r_n_145__60_,r_n_145__59_,
  r_n_145__58_,r_n_145__57_,r_n_145__56_,r_n_145__55_,r_n_145__54_,r_n_145__53_,
  r_n_145__52_,r_n_145__51_,r_n_145__50_,r_n_145__49_,r_n_145__48_,r_n_145__47_,
  r_n_145__46_,r_n_145__45_,r_n_145__44_,r_n_145__43_,r_n_145__42_,r_n_145__41_,r_n_145__40_,
  r_n_145__39_,r_n_145__38_,r_n_145__37_,r_n_145__36_,r_n_145__35_,r_n_145__34_,
  r_n_145__33_,r_n_145__32_,r_n_145__31_,r_n_145__30_,r_n_145__29_,r_n_145__28_,
  r_n_145__27_,r_n_145__26_,r_n_145__25_,r_n_145__24_,r_n_145__23_,r_n_145__22_,
  r_n_145__21_,r_n_145__20_,r_n_145__19_,r_n_145__18_,r_n_145__17_,r_n_145__16_,
  r_n_145__15_,r_n_145__14_,r_n_145__13_,r_n_145__12_,r_n_145__11_,r_n_145__10_,
  r_n_145__9_,r_n_145__8_,r_n_145__7_,r_n_145__6_,r_n_145__5_,r_n_145__4_,r_n_145__3_,
  r_n_145__2_,r_n_145__1_,r_n_145__0_,r_n_160__63_,r_n_160__62_,r_n_160__61_,
  r_n_160__60_,r_n_160__59_,r_n_160__58_,r_n_160__57_,r_n_160__56_,r_n_160__55_,r_n_160__54_,
  r_n_160__53_,r_n_160__52_,r_n_160__51_,r_n_160__50_,r_n_160__49_,r_n_160__48_,
  r_n_160__47_,r_n_160__46_,r_n_160__45_,r_n_160__44_,r_n_160__43_,r_n_160__42_,
  r_n_160__41_,r_n_160__40_,r_n_160__39_,r_n_160__38_,r_n_160__37_,r_n_160__36_,
  r_n_160__35_,r_n_160__34_,r_n_160__33_,r_n_160__32_,r_n_160__31_,r_n_160__30_,
  r_n_160__29_,r_n_160__28_,r_n_160__27_,r_n_160__26_,r_n_160__25_,r_n_160__24_,
  r_n_160__23_,r_n_160__22_,r_n_160__21_,r_n_160__20_,r_n_160__19_,r_n_160__18_,
  r_n_160__17_,r_n_160__16_,r_n_160__15_,r_n_160__14_,r_n_160__13_,r_n_160__12_,r_n_160__11_,
  r_n_160__10_,r_n_160__9_,r_n_160__8_,r_n_160__7_,r_n_160__6_,r_n_160__5_,
  r_n_160__4_,r_n_160__3_,r_n_160__2_,r_n_160__1_,r_n_160__0_,r_n_159__63_,r_n_159__62_,
  r_n_159__61_,r_n_159__60_,r_n_159__59_,r_n_159__58_,r_n_159__57_,r_n_159__56_,
  r_n_159__55_,r_n_159__54_,r_n_159__53_,r_n_159__52_,r_n_159__51_,r_n_159__50_,
  r_n_159__49_,r_n_159__48_,r_n_159__47_,r_n_159__46_,r_n_159__45_,r_n_159__44_,
  r_n_159__43_,r_n_159__42_,r_n_159__41_,r_n_159__40_,r_n_159__39_,r_n_159__38_,
  r_n_159__37_,r_n_159__36_,r_n_159__35_,r_n_159__34_,r_n_159__33_,r_n_159__32_,
  r_n_159__31_,r_n_159__30_,r_n_159__29_,r_n_159__28_,r_n_159__27_,r_n_159__26_,r_n_159__25_,
  r_n_159__24_,r_n_159__23_,r_n_159__22_,r_n_159__21_,r_n_159__20_,r_n_159__19_,
  r_n_159__18_,r_n_159__17_,r_n_159__16_,r_n_159__15_,r_n_159__14_,r_n_159__13_,
  r_n_159__12_,r_n_159__11_,r_n_159__10_,r_n_159__9_,r_n_159__8_,r_n_159__7_,
  r_n_159__6_,r_n_159__5_,r_n_159__4_,r_n_159__3_,r_n_159__2_,r_n_159__1_,r_n_159__0_,
  r_n_158__63_,r_n_158__62_,r_n_158__61_,r_n_158__60_,r_n_158__59_,r_n_158__58_,
  r_n_158__57_,r_n_158__56_,r_n_158__55_,r_n_158__54_,r_n_158__53_,r_n_158__52_,
  r_n_158__51_,r_n_158__50_,r_n_158__49_,r_n_158__48_,r_n_158__47_,r_n_158__46_,
  r_n_158__45_,r_n_158__44_,r_n_158__43_,r_n_158__42_,r_n_158__41_,r_n_158__40_,r_n_158__39_,
  r_n_158__38_,r_n_158__37_,r_n_158__36_,r_n_158__35_,r_n_158__34_,r_n_158__33_,
  r_n_158__32_,r_n_158__31_,r_n_158__30_,r_n_158__29_,r_n_158__28_,r_n_158__27_,
  r_n_158__26_,r_n_158__25_,r_n_158__24_,r_n_158__23_,r_n_158__22_,r_n_158__21_,
  r_n_158__20_,r_n_158__19_,r_n_158__18_,r_n_158__17_,r_n_158__16_,r_n_158__15_,
  r_n_158__14_,r_n_158__13_,r_n_158__12_,r_n_158__11_,r_n_158__10_,r_n_158__9_,r_n_158__8_,
  r_n_158__7_,r_n_158__6_,r_n_158__5_,r_n_158__4_,r_n_158__3_,r_n_158__2_,
  r_n_158__1_,r_n_158__0_,r_n_157__63_,r_n_157__62_,r_n_157__61_,r_n_157__60_,
  r_n_157__59_,r_n_157__58_,r_n_157__57_,r_n_157__56_,r_n_157__55_,r_n_157__54_,r_n_157__53_,
  r_n_157__52_,r_n_157__51_,r_n_157__50_,r_n_157__49_,r_n_157__48_,r_n_157__47_,
  r_n_157__46_,r_n_157__45_,r_n_157__44_,r_n_157__43_,r_n_157__42_,r_n_157__41_,
  r_n_157__40_,r_n_157__39_,r_n_157__38_,r_n_157__37_,r_n_157__36_,r_n_157__35_,
  r_n_157__34_,r_n_157__33_,r_n_157__32_,r_n_157__31_,r_n_157__30_,r_n_157__29_,
  r_n_157__28_,r_n_157__27_,r_n_157__26_,r_n_157__25_,r_n_157__24_,r_n_157__23_,
  r_n_157__22_,r_n_157__21_,r_n_157__20_,r_n_157__19_,r_n_157__18_,r_n_157__17_,r_n_157__16_,
  r_n_157__15_,r_n_157__14_,r_n_157__13_,r_n_157__12_,r_n_157__11_,r_n_157__10_,
  r_n_157__9_,r_n_157__8_,r_n_157__7_,r_n_157__6_,r_n_157__5_,r_n_157__4_,
  r_n_157__3_,r_n_157__2_,r_n_157__1_,r_n_157__0_,r_n_156__63_,r_n_156__62_,r_n_156__61_,
  r_n_156__60_,r_n_156__59_,r_n_156__58_,r_n_156__57_,r_n_156__56_,r_n_156__55_,
  r_n_156__54_,r_n_156__53_,r_n_156__52_,r_n_156__51_,r_n_156__50_,r_n_156__49_,
  r_n_156__48_,r_n_156__47_,r_n_156__46_,r_n_156__45_,r_n_156__44_,r_n_156__43_,
  r_n_156__42_,r_n_156__41_,r_n_156__40_,r_n_156__39_,r_n_156__38_,r_n_156__37_,
  r_n_156__36_,r_n_156__35_,r_n_156__34_,r_n_156__33_,r_n_156__32_,r_n_156__31_,r_n_156__30_,
  r_n_156__29_,r_n_156__28_,r_n_156__27_,r_n_156__26_,r_n_156__25_,r_n_156__24_,
  r_n_156__23_,r_n_156__22_,r_n_156__21_,r_n_156__20_,r_n_156__19_,r_n_156__18_,
  r_n_156__17_,r_n_156__16_,r_n_156__15_,r_n_156__14_,r_n_156__13_,r_n_156__12_,
  r_n_156__11_,r_n_156__10_,r_n_156__9_,r_n_156__8_,r_n_156__7_,r_n_156__6_,r_n_156__5_,
  r_n_156__4_,r_n_156__3_,r_n_156__2_,r_n_156__1_,r_n_156__0_,r_n_155__63_,
  r_n_155__62_,r_n_155__61_,r_n_155__60_,r_n_155__59_,r_n_155__58_,r_n_155__57_,
  r_n_155__56_,r_n_155__55_,r_n_155__54_,r_n_155__53_,r_n_155__52_,r_n_155__51_,
  r_n_155__50_,r_n_155__49_,r_n_155__48_,r_n_155__47_,r_n_155__46_,r_n_155__45_,r_n_155__44_,
  r_n_155__43_,r_n_155__42_,r_n_155__41_,r_n_155__40_,r_n_155__39_,r_n_155__38_,
  r_n_155__37_,r_n_155__36_,r_n_155__35_,r_n_155__34_,r_n_155__33_,r_n_155__32_,
  r_n_155__31_,r_n_155__30_,r_n_155__29_,r_n_155__28_,r_n_155__27_,r_n_155__26_,
  r_n_155__25_,r_n_155__24_,r_n_155__23_,r_n_155__22_,r_n_155__21_,r_n_155__20_,
  r_n_155__19_,r_n_155__18_,r_n_155__17_,r_n_155__16_,r_n_155__15_,r_n_155__14_,
  r_n_155__13_,r_n_155__12_,r_n_155__11_,r_n_155__10_,r_n_155__9_,r_n_155__8_,r_n_155__7_,
  r_n_155__6_,r_n_155__5_,r_n_155__4_,r_n_155__3_,r_n_155__2_,r_n_155__1_,
  r_n_155__0_,r_n_154__63_,r_n_154__62_,r_n_154__61_,r_n_154__60_,r_n_154__59_,r_n_154__58_,
  r_n_154__57_,r_n_154__56_,r_n_154__55_,r_n_154__54_,r_n_154__53_,r_n_154__52_,
  r_n_154__51_,r_n_154__50_,r_n_154__49_,r_n_154__48_,r_n_154__47_,r_n_154__46_,
  r_n_154__45_,r_n_154__44_,r_n_154__43_,r_n_154__42_,r_n_154__41_,r_n_154__40_,
  r_n_154__39_,r_n_154__38_,r_n_154__37_,r_n_154__36_,r_n_154__35_,r_n_154__34_,
  r_n_154__33_,r_n_154__32_,r_n_154__31_,r_n_154__30_,r_n_154__29_,r_n_154__28_,
  r_n_154__27_,r_n_154__26_,r_n_154__25_,r_n_154__24_,r_n_154__23_,r_n_154__22_,
  r_n_154__21_,r_n_154__20_,r_n_154__19_,r_n_154__18_,r_n_154__17_,r_n_154__16_,r_n_154__15_,
  r_n_154__14_,r_n_154__13_,r_n_154__12_,r_n_154__11_,r_n_154__10_,r_n_154__9_,
  r_n_154__8_,r_n_154__7_,r_n_154__6_,r_n_154__5_,r_n_154__4_,r_n_154__3_,r_n_154__2_,
  r_n_154__1_,r_n_154__0_,r_n_153__63_,r_n_153__62_,r_n_153__61_,r_n_153__60_,
  r_n_153__59_,r_n_153__58_,r_n_153__57_,r_n_153__56_,r_n_153__55_,r_n_153__54_,
  r_n_153__53_,r_n_153__52_,r_n_153__51_,r_n_153__50_,r_n_153__49_,r_n_153__48_,
  r_n_153__47_,r_n_153__46_,r_n_153__45_,r_n_153__44_,r_n_153__43_,r_n_153__42_,
  r_n_153__41_,r_n_153__40_,r_n_153__39_,r_n_153__38_,r_n_153__37_,r_n_153__36_,
  r_n_153__35_,r_n_153__34_,r_n_153__33_,r_n_153__32_,r_n_153__31_,r_n_153__30_,r_n_153__29_,
  r_n_153__28_,r_n_153__27_,r_n_153__26_,r_n_153__25_,r_n_153__24_,r_n_153__23_,
  r_n_153__22_,r_n_153__21_,r_n_153__20_,r_n_153__19_,r_n_153__18_,r_n_153__17_,
  r_n_153__16_,r_n_153__15_,r_n_153__14_,r_n_153__13_,r_n_153__12_,r_n_153__11_,
  r_n_153__10_,r_n_153__9_,r_n_153__8_,r_n_153__7_,r_n_153__6_,r_n_153__5_,r_n_153__4_,
  r_n_153__3_,r_n_153__2_,r_n_153__1_,r_n_153__0_,r_n_168__63_,r_n_168__62_,
  r_n_168__61_,r_n_168__60_,r_n_168__59_,r_n_168__58_,r_n_168__57_,r_n_168__56_,
  r_n_168__55_,r_n_168__54_,r_n_168__53_,r_n_168__52_,r_n_168__51_,r_n_168__50_,
  r_n_168__49_,r_n_168__48_,r_n_168__47_,r_n_168__46_,r_n_168__45_,r_n_168__44_,r_n_168__43_,
  r_n_168__42_,r_n_168__41_,r_n_168__40_,r_n_168__39_,r_n_168__38_,r_n_168__37_,
  r_n_168__36_,r_n_168__35_,r_n_168__34_,r_n_168__33_,r_n_168__32_,r_n_168__31_,
  r_n_168__30_,r_n_168__29_,r_n_168__28_,r_n_168__27_,r_n_168__26_,r_n_168__25_,
  r_n_168__24_,r_n_168__23_,r_n_168__22_,r_n_168__21_,r_n_168__20_,r_n_168__19_,
  r_n_168__18_,r_n_168__17_,r_n_168__16_,r_n_168__15_,r_n_168__14_,r_n_168__13_,
  r_n_168__12_,r_n_168__11_,r_n_168__10_,r_n_168__9_,r_n_168__8_,r_n_168__7_,r_n_168__6_,
  r_n_168__5_,r_n_168__4_,r_n_168__3_,r_n_168__2_,r_n_168__1_,r_n_168__0_,
  r_n_167__63_,r_n_167__62_,r_n_167__61_,r_n_167__60_,r_n_167__59_,r_n_167__58_,r_n_167__57_,
  r_n_167__56_,r_n_167__55_,r_n_167__54_,r_n_167__53_,r_n_167__52_,r_n_167__51_,
  r_n_167__50_,r_n_167__49_,r_n_167__48_,r_n_167__47_,r_n_167__46_,r_n_167__45_,
  r_n_167__44_,r_n_167__43_,r_n_167__42_,r_n_167__41_,r_n_167__40_,r_n_167__39_,
  r_n_167__38_,r_n_167__37_,r_n_167__36_,r_n_167__35_,r_n_167__34_,r_n_167__33_,
  r_n_167__32_,r_n_167__31_,r_n_167__30_,r_n_167__29_,r_n_167__28_,r_n_167__27_,
  r_n_167__26_,r_n_167__25_,r_n_167__24_,r_n_167__23_,r_n_167__22_,r_n_167__21_,r_n_167__20_,
  r_n_167__19_,r_n_167__18_,r_n_167__17_,r_n_167__16_,r_n_167__15_,r_n_167__14_,
  r_n_167__13_,r_n_167__12_,r_n_167__11_,r_n_167__10_,r_n_167__9_,r_n_167__8_,
  r_n_167__7_,r_n_167__6_,r_n_167__5_,r_n_167__4_,r_n_167__3_,r_n_167__2_,r_n_167__1_,
  r_n_167__0_,r_n_166__63_,r_n_166__62_,r_n_166__61_,r_n_166__60_,r_n_166__59_,
  r_n_166__58_,r_n_166__57_,r_n_166__56_,r_n_166__55_,r_n_166__54_,r_n_166__53_,
  r_n_166__52_,r_n_166__51_,r_n_166__50_,r_n_166__49_,r_n_166__48_,r_n_166__47_,
  r_n_166__46_,r_n_166__45_,r_n_166__44_,r_n_166__43_,r_n_166__42_,r_n_166__41_,
  r_n_166__40_,r_n_166__39_,r_n_166__38_,r_n_166__37_,r_n_166__36_,r_n_166__35_,r_n_166__34_,
  r_n_166__33_,r_n_166__32_,r_n_166__31_,r_n_166__30_,r_n_166__29_,r_n_166__28_,
  r_n_166__27_,r_n_166__26_,r_n_166__25_,r_n_166__24_,r_n_166__23_,r_n_166__22_,
  r_n_166__21_,r_n_166__20_,r_n_166__19_,r_n_166__18_,r_n_166__17_,r_n_166__16_,
  r_n_166__15_,r_n_166__14_,r_n_166__13_,r_n_166__12_,r_n_166__11_,r_n_166__10_,
  r_n_166__9_,r_n_166__8_,r_n_166__7_,r_n_166__6_,r_n_166__5_,r_n_166__4_,r_n_166__3_,
  r_n_166__2_,r_n_166__1_,r_n_166__0_,r_n_165__63_,r_n_165__62_,r_n_165__61_,
  r_n_165__60_,r_n_165__59_,r_n_165__58_,r_n_165__57_,r_n_165__56_,r_n_165__55_,
  r_n_165__54_,r_n_165__53_,r_n_165__52_,r_n_165__51_,r_n_165__50_,r_n_165__49_,r_n_165__48_,
  r_n_165__47_,r_n_165__46_,r_n_165__45_,r_n_165__44_,r_n_165__43_,r_n_165__42_,
  r_n_165__41_,r_n_165__40_,r_n_165__39_,r_n_165__38_,r_n_165__37_,r_n_165__36_,
  r_n_165__35_,r_n_165__34_,r_n_165__33_,r_n_165__32_,r_n_165__31_,r_n_165__30_,
  r_n_165__29_,r_n_165__28_,r_n_165__27_,r_n_165__26_,r_n_165__25_,r_n_165__24_,
  r_n_165__23_,r_n_165__22_,r_n_165__21_,r_n_165__20_,r_n_165__19_,r_n_165__18_,
  r_n_165__17_,r_n_165__16_,r_n_165__15_,r_n_165__14_,r_n_165__13_,r_n_165__12_,
  r_n_165__11_,r_n_165__10_,r_n_165__9_,r_n_165__8_,r_n_165__7_,r_n_165__6_,r_n_165__5_,
  r_n_165__4_,r_n_165__3_,r_n_165__2_,r_n_165__1_,r_n_165__0_,r_n_164__63_,r_n_164__62_,
  r_n_164__61_,r_n_164__60_,r_n_164__59_,r_n_164__58_,r_n_164__57_,r_n_164__56_,
  r_n_164__55_,r_n_164__54_,r_n_164__53_,r_n_164__52_,r_n_164__51_,r_n_164__50_,
  r_n_164__49_,r_n_164__48_,r_n_164__47_,r_n_164__46_,r_n_164__45_,r_n_164__44_,
  r_n_164__43_,r_n_164__42_,r_n_164__41_,r_n_164__40_,r_n_164__39_,r_n_164__38_,
  r_n_164__37_,r_n_164__36_,r_n_164__35_,r_n_164__34_,r_n_164__33_,r_n_164__32_,
  r_n_164__31_,r_n_164__30_,r_n_164__29_,r_n_164__28_,r_n_164__27_,r_n_164__26_,
  r_n_164__25_,r_n_164__24_,r_n_164__23_,r_n_164__22_,r_n_164__21_,r_n_164__20_,r_n_164__19_,
  r_n_164__18_,r_n_164__17_,r_n_164__16_,r_n_164__15_,r_n_164__14_,r_n_164__13_,
  r_n_164__12_,r_n_164__11_,r_n_164__10_,r_n_164__9_,r_n_164__8_,r_n_164__7_,
  r_n_164__6_,r_n_164__5_,r_n_164__4_,r_n_164__3_,r_n_164__2_,r_n_164__1_,r_n_164__0_,
  r_n_163__63_,r_n_163__62_,r_n_163__61_,r_n_163__60_,r_n_163__59_,r_n_163__58_,
  r_n_163__57_,r_n_163__56_,r_n_163__55_,r_n_163__54_,r_n_163__53_,r_n_163__52_,
  r_n_163__51_,r_n_163__50_,r_n_163__49_,r_n_163__48_,r_n_163__47_,r_n_163__46_,
  r_n_163__45_,r_n_163__44_,r_n_163__43_,r_n_163__42_,r_n_163__41_,r_n_163__40_,
  r_n_163__39_,r_n_163__38_,r_n_163__37_,r_n_163__36_,r_n_163__35_,r_n_163__34_,r_n_163__33_,
  r_n_163__32_,r_n_163__31_,r_n_163__30_,r_n_163__29_,r_n_163__28_,r_n_163__27_,
  r_n_163__26_,r_n_163__25_,r_n_163__24_,r_n_163__23_,r_n_163__22_,r_n_163__21_,
  r_n_163__20_,r_n_163__19_,r_n_163__18_,r_n_163__17_,r_n_163__16_,r_n_163__15_,
  r_n_163__14_,r_n_163__13_,r_n_163__12_,r_n_163__11_,r_n_163__10_,r_n_163__9_,
  r_n_163__8_,r_n_163__7_,r_n_163__6_,r_n_163__5_,r_n_163__4_,r_n_163__3_,r_n_163__2_,
  r_n_163__1_,r_n_163__0_,r_n_162__63_,r_n_162__62_,r_n_162__61_,r_n_162__60_,
  r_n_162__59_,r_n_162__58_,r_n_162__57_,r_n_162__56_,r_n_162__55_,r_n_162__54_,
  r_n_162__53_,r_n_162__52_,r_n_162__51_,r_n_162__50_,r_n_162__49_,r_n_162__48_,r_n_162__47_,
  r_n_162__46_,r_n_162__45_,r_n_162__44_,r_n_162__43_,r_n_162__42_,r_n_162__41_,
  r_n_162__40_,r_n_162__39_,r_n_162__38_,r_n_162__37_,r_n_162__36_,r_n_162__35_,
  r_n_162__34_,r_n_162__33_,r_n_162__32_,r_n_162__31_,r_n_162__30_,r_n_162__29_,
  r_n_162__28_,r_n_162__27_,r_n_162__26_,r_n_162__25_,r_n_162__24_,r_n_162__23_,
  r_n_162__22_,r_n_162__21_,r_n_162__20_,r_n_162__19_,r_n_162__18_,r_n_162__17_,
  r_n_162__16_,r_n_162__15_,r_n_162__14_,r_n_162__13_,r_n_162__12_,r_n_162__11_,r_n_162__10_,
  r_n_162__9_,r_n_162__8_,r_n_162__7_,r_n_162__6_,r_n_162__5_,r_n_162__4_,
  r_n_162__3_,r_n_162__2_,r_n_162__1_,r_n_162__0_,r_n_161__63_,r_n_161__62_,r_n_161__61_,
  r_n_161__60_,r_n_161__59_,r_n_161__58_,r_n_161__57_,r_n_161__56_,r_n_161__55_,
  r_n_161__54_,r_n_161__53_,r_n_161__52_,r_n_161__51_,r_n_161__50_,r_n_161__49_,
  r_n_161__48_,r_n_161__47_,r_n_161__46_,r_n_161__45_,r_n_161__44_,r_n_161__43_,
  r_n_161__42_,r_n_161__41_,r_n_161__40_,r_n_161__39_,r_n_161__38_,r_n_161__37_,
  r_n_161__36_,r_n_161__35_,r_n_161__34_,r_n_161__33_,r_n_161__32_,r_n_161__31_,
  r_n_161__30_,r_n_161__29_,r_n_161__28_,r_n_161__27_,r_n_161__26_,r_n_161__25_,r_n_161__24_,
  r_n_161__23_,r_n_161__22_,r_n_161__21_,r_n_161__20_,r_n_161__19_,r_n_161__18_,
  r_n_161__17_,r_n_161__16_,r_n_161__15_,r_n_161__14_,r_n_161__13_,r_n_161__12_,
  r_n_161__11_,r_n_161__10_,r_n_161__9_,r_n_161__8_,r_n_161__7_,r_n_161__6_,
  r_n_161__5_,r_n_161__4_,r_n_161__3_,r_n_161__2_,r_n_161__1_,r_n_161__0_,r_n_176__63_,
  r_n_176__62_,r_n_176__61_,r_n_176__60_,r_n_176__59_,r_n_176__58_,r_n_176__57_,
  r_n_176__56_,r_n_176__55_,r_n_176__54_,r_n_176__53_,r_n_176__52_,r_n_176__51_,
  r_n_176__50_,r_n_176__49_,r_n_176__48_,r_n_176__47_,r_n_176__46_,r_n_176__45_,
  r_n_176__44_,r_n_176__43_,r_n_176__42_,r_n_176__41_,r_n_176__40_,r_n_176__39_,r_n_176__38_,
  r_n_176__37_,r_n_176__36_,r_n_176__35_,r_n_176__34_,r_n_176__33_,r_n_176__32_,
  r_n_176__31_,r_n_176__30_,r_n_176__29_,r_n_176__28_,r_n_176__27_,r_n_176__26_,
  r_n_176__25_,r_n_176__24_,r_n_176__23_,r_n_176__22_,r_n_176__21_,r_n_176__20_,
  r_n_176__19_,r_n_176__18_,r_n_176__17_,r_n_176__16_,r_n_176__15_,r_n_176__14_,
  r_n_176__13_,r_n_176__12_,r_n_176__11_,r_n_176__10_,r_n_176__9_,r_n_176__8_,r_n_176__7_,
  r_n_176__6_,r_n_176__5_,r_n_176__4_,r_n_176__3_,r_n_176__2_,r_n_176__1_,
  r_n_176__0_,r_n_175__63_,r_n_175__62_,r_n_175__61_,r_n_175__60_,r_n_175__59_,
  r_n_175__58_,r_n_175__57_,r_n_175__56_,r_n_175__55_,r_n_175__54_,r_n_175__53_,r_n_175__52_,
  r_n_175__51_,r_n_175__50_,r_n_175__49_,r_n_175__48_,r_n_175__47_,r_n_175__46_,
  r_n_175__45_,r_n_175__44_,r_n_175__43_,r_n_175__42_,r_n_175__41_,r_n_175__40_,
  r_n_175__39_,r_n_175__38_,r_n_175__37_,r_n_175__36_,r_n_175__35_,r_n_175__34_,
  r_n_175__33_,r_n_175__32_,r_n_175__31_,r_n_175__30_,r_n_175__29_,r_n_175__28_,
  r_n_175__27_,r_n_175__26_,r_n_175__25_,r_n_175__24_,r_n_175__23_,r_n_175__22_,
  r_n_175__21_,r_n_175__20_,r_n_175__19_,r_n_175__18_,r_n_175__17_,r_n_175__16_,
  r_n_175__15_,r_n_175__14_,r_n_175__13_,r_n_175__12_,r_n_175__11_,r_n_175__10_,r_n_175__9_,
  r_n_175__8_,r_n_175__7_,r_n_175__6_,r_n_175__5_,r_n_175__4_,r_n_175__3_,
  r_n_175__2_,r_n_175__1_,r_n_175__0_,r_n_174__63_,r_n_174__62_,r_n_174__61_,r_n_174__60_,
  r_n_174__59_,r_n_174__58_,r_n_174__57_,r_n_174__56_,r_n_174__55_,r_n_174__54_,
  r_n_174__53_,r_n_174__52_,r_n_174__51_,r_n_174__50_,r_n_174__49_,r_n_174__48_,
  r_n_174__47_,r_n_174__46_,r_n_174__45_,r_n_174__44_,r_n_174__43_,r_n_174__42_,
  r_n_174__41_,r_n_174__40_,r_n_174__39_,r_n_174__38_,r_n_174__37_,r_n_174__36_,
  r_n_174__35_,r_n_174__34_,r_n_174__33_,r_n_174__32_,r_n_174__31_,r_n_174__30_,
  r_n_174__29_,r_n_174__28_,r_n_174__27_,r_n_174__26_,r_n_174__25_,r_n_174__24_,r_n_174__23_,
  r_n_174__22_,r_n_174__21_,r_n_174__20_,r_n_174__19_,r_n_174__18_,r_n_174__17_,
  r_n_174__16_,r_n_174__15_,r_n_174__14_,r_n_174__13_,r_n_174__12_,r_n_174__11_,
  r_n_174__10_,r_n_174__9_,r_n_174__8_,r_n_174__7_,r_n_174__6_,r_n_174__5_,r_n_174__4_,
  r_n_174__3_,r_n_174__2_,r_n_174__1_,r_n_174__0_,r_n_173__63_,r_n_173__62_,
  r_n_173__61_,r_n_173__60_,r_n_173__59_,r_n_173__58_,r_n_173__57_,r_n_173__56_,
  r_n_173__55_,r_n_173__54_,r_n_173__53_,r_n_173__52_,r_n_173__51_,r_n_173__50_,
  r_n_173__49_,r_n_173__48_,r_n_173__47_,r_n_173__46_,r_n_173__45_,r_n_173__44_,
  r_n_173__43_,r_n_173__42_,r_n_173__41_,r_n_173__40_,r_n_173__39_,r_n_173__38_,r_n_173__37_,
  r_n_173__36_,r_n_173__35_,r_n_173__34_,r_n_173__33_,r_n_173__32_,r_n_173__31_,
  r_n_173__30_,r_n_173__29_,r_n_173__28_,r_n_173__27_,r_n_173__26_,r_n_173__25_,
  r_n_173__24_,r_n_173__23_,r_n_173__22_,r_n_173__21_,r_n_173__20_,r_n_173__19_,
  r_n_173__18_,r_n_173__17_,r_n_173__16_,r_n_173__15_,r_n_173__14_,r_n_173__13_,
  r_n_173__12_,r_n_173__11_,r_n_173__10_,r_n_173__9_,r_n_173__8_,r_n_173__7_,r_n_173__6_,
  r_n_173__5_,r_n_173__4_,r_n_173__3_,r_n_173__2_,r_n_173__1_,r_n_173__0_,
  r_n_172__63_,r_n_172__62_,r_n_172__61_,r_n_172__60_,r_n_172__59_,r_n_172__58_,
  r_n_172__57_,r_n_172__56_,r_n_172__55_,r_n_172__54_,r_n_172__53_,r_n_172__52_,r_n_172__51_,
  r_n_172__50_,r_n_172__49_,r_n_172__48_,r_n_172__47_,r_n_172__46_,r_n_172__45_,
  r_n_172__44_,r_n_172__43_,r_n_172__42_,r_n_172__41_,r_n_172__40_,r_n_172__39_,
  r_n_172__38_,r_n_172__37_,r_n_172__36_,r_n_172__35_,r_n_172__34_,r_n_172__33_,
  r_n_172__32_,r_n_172__31_,r_n_172__30_,r_n_172__29_,r_n_172__28_,r_n_172__27_,
  r_n_172__26_,r_n_172__25_,r_n_172__24_,r_n_172__23_,r_n_172__22_,r_n_172__21_,
  r_n_172__20_,r_n_172__19_,r_n_172__18_,r_n_172__17_,r_n_172__16_,r_n_172__15_,r_n_172__14_,
  r_n_172__13_,r_n_172__12_,r_n_172__11_,r_n_172__10_,r_n_172__9_,r_n_172__8_,
  r_n_172__7_,r_n_172__6_,r_n_172__5_,r_n_172__4_,r_n_172__3_,r_n_172__2_,r_n_172__1_,
  r_n_172__0_,r_n_171__63_,r_n_171__62_,r_n_171__61_,r_n_171__60_,r_n_171__59_,
  r_n_171__58_,r_n_171__57_,r_n_171__56_,r_n_171__55_,r_n_171__54_,r_n_171__53_,
  r_n_171__52_,r_n_171__51_,r_n_171__50_,r_n_171__49_,r_n_171__48_,r_n_171__47_,
  r_n_171__46_,r_n_171__45_,r_n_171__44_,r_n_171__43_,r_n_171__42_,r_n_171__41_,
  r_n_171__40_,r_n_171__39_,r_n_171__38_,r_n_171__37_,r_n_171__36_,r_n_171__35_,
  r_n_171__34_,r_n_171__33_,r_n_171__32_,r_n_171__31_,r_n_171__30_,r_n_171__29_,r_n_171__28_,
  r_n_171__27_,r_n_171__26_,r_n_171__25_,r_n_171__24_,r_n_171__23_,r_n_171__22_,
  r_n_171__21_,r_n_171__20_,r_n_171__19_,r_n_171__18_,r_n_171__17_,r_n_171__16_,
  r_n_171__15_,r_n_171__14_,r_n_171__13_,r_n_171__12_,r_n_171__11_,r_n_171__10_,
  r_n_171__9_,r_n_171__8_,r_n_171__7_,r_n_171__6_,r_n_171__5_,r_n_171__4_,r_n_171__3_,
  r_n_171__2_,r_n_171__1_,r_n_171__0_,r_n_170__63_,r_n_170__62_,r_n_170__61_,
  r_n_170__60_,r_n_170__59_,r_n_170__58_,r_n_170__57_,r_n_170__56_,r_n_170__55_,
  r_n_170__54_,r_n_170__53_,r_n_170__52_,r_n_170__51_,r_n_170__50_,r_n_170__49_,
  r_n_170__48_,r_n_170__47_,r_n_170__46_,r_n_170__45_,r_n_170__44_,r_n_170__43_,r_n_170__42_,
  r_n_170__41_,r_n_170__40_,r_n_170__39_,r_n_170__38_,r_n_170__37_,r_n_170__36_,
  r_n_170__35_,r_n_170__34_,r_n_170__33_,r_n_170__32_,r_n_170__31_,r_n_170__30_,
  r_n_170__29_,r_n_170__28_,r_n_170__27_,r_n_170__26_,r_n_170__25_,r_n_170__24_,
  r_n_170__23_,r_n_170__22_,r_n_170__21_,r_n_170__20_,r_n_170__19_,r_n_170__18_,
  r_n_170__17_,r_n_170__16_,r_n_170__15_,r_n_170__14_,r_n_170__13_,r_n_170__12_,
  r_n_170__11_,r_n_170__10_,r_n_170__9_,r_n_170__8_,r_n_170__7_,r_n_170__6_,r_n_170__5_,
  r_n_170__4_,r_n_170__3_,r_n_170__2_,r_n_170__1_,r_n_170__0_,r_n_169__63_,
  r_n_169__62_,r_n_169__61_,r_n_169__60_,r_n_169__59_,r_n_169__58_,r_n_169__57_,r_n_169__56_,
  r_n_169__55_,r_n_169__54_,r_n_169__53_,r_n_169__52_,r_n_169__51_,r_n_169__50_,
  r_n_169__49_,r_n_169__48_,r_n_169__47_,r_n_169__46_,r_n_169__45_,r_n_169__44_,
  r_n_169__43_,r_n_169__42_,r_n_169__41_,r_n_169__40_,r_n_169__39_,r_n_169__38_,
  r_n_169__37_,r_n_169__36_,r_n_169__35_,r_n_169__34_,r_n_169__33_,r_n_169__32_,
  r_n_169__31_,r_n_169__30_,r_n_169__29_,r_n_169__28_,r_n_169__27_,r_n_169__26_,
  r_n_169__25_,r_n_169__24_,r_n_169__23_,r_n_169__22_,r_n_169__21_,r_n_169__20_,
  r_n_169__19_,r_n_169__18_,r_n_169__17_,r_n_169__16_,r_n_169__15_,r_n_169__14_,r_n_169__13_,
  r_n_169__12_,r_n_169__11_,r_n_169__10_,r_n_169__9_,r_n_169__8_,r_n_169__7_,
  r_n_169__6_,r_n_169__5_,r_n_169__4_,r_n_169__3_,r_n_169__2_,r_n_169__1_,r_n_169__0_,
  r_n_184__63_,r_n_184__62_,r_n_184__61_,r_n_184__60_,r_n_184__59_,r_n_184__58_,
  r_n_184__57_,r_n_184__56_,r_n_184__55_,r_n_184__54_,r_n_184__53_,r_n_184__52_,
  r_n_184__51_,r_n_184__50_,r_n_184__49_,r_n_184__48_,r_n_184__47_,r_n_184__46_,
  r_n_184__45_,r_n_184__44_,r_n_184__43_,r_n_184__42_,r_n_184__41_,r_n_184__40_,
  r_n_184__39_,r_n_184__38_,r_n_184__37_,r_n_184__36_,r_n_184__35_,r_n_184__34_,
  r_n_184__33_,r_n_184__32_,r_n_184__31_,r_n_184__30_,r_n_184__29_,r_n_184__28_,r_n_184__27_,
  r_n_184__26_,r_n_184__25_,r_n_184__24_,r_n_184__23_,r_n_184__22_,r_n_184__21_,
  r_n_184__20_,r_n_184__19_,r_n_184__18_,r_n_184__17_,r_n_184__16_,r_n_184__15_,
  r_n_184__14_,r_n_184__13_,r_n_184__12_,r_n_184__11_,r_n_184__10_,r_n_184__9_,
  r_n_184__8_,r_n_184__7_,r_n_184__6_,r_n_184__5_,r_n_184__4_,r_n_184__3_,r_n_184__2_,
  r_n_184__1_,r_n_184__0_,r_n_183__63_,r_n_183__62_,r_n_183__61_,r_n_183__60_,
  r_n_183__59_,r_n_183__58_,r_n_183__57_,r_n_183__56_,r_n_183__55_,r_n_183__54_,
  r_n_183__53_,r_n_183__52_,r_n_183__51_,r_n_183__50_,r_n_183__49_,r_n_183__48_,
  r_n_183__47_,r_n_183__46_,r_n_183__45_,r_n_183__44_,r_n_183__43_,r_n_183__42_,r_n_183__41_,
  r_n_183__40_,r_n_183__39_,r_n_183__38_,r_n_183__37_,r_n_183__36_,r_n_183__35_,
  r_n_183__34_,r_n_183__33_,r_n_183__32_,r_n_183__31_,r_n_183__30_,r_n_183__29_,
  r_n_183__28_,r_n_183__27_,r_n_183__26_,r_n_183__25_,r_n_183__24_,r_n_183__23_,
  r_n_183__22_,r_n_183__21_,r_n_183__20_,r_n_183__19_,r_n_183__18_,r_n_183__17_,
  r_n_183__16_,r_n_183__15_,r_n_183__14_,r_n_183__13_,r_n_183__12_,r_n_183__11_,
  r_n_183__10_,r_n_183__9_,r_n_183__8_,r_n_183__7_,r_n_183__6_,r_n_183__5_,r_n_183__4_,
  r_n_183__3_,r_n_183__2_,r_n_183__1_,r_n_183__0_,r_n_182__63_,r_n_182__62_,
  r_n_182__61_,r_n_182__60_,r_n_182__59_,r_n_182__58_,r_n_182__57_,r_n_182__56_,r_n_182__55_,
  r_n_182__54_,r_n_182__53_,r_n_182__52_,r_n_182__51_,r_n_182__50_,r_n_182__49_,
  r_n_182__48_,r_n_182__47_,r_n_182__46_,r_n_182__45_,r_n_182__44_,r_n_182__43_,
  r_n_182__42_,r_n_182__41_,r_n_182__40_,r_n_182__39_,r_n_182__38_,r_n_182__37_,
  r_n_182__36_,r_n_182__35_,r_n_182__34_,r_n_182__33_,r_n_182__32_,r_n_182__31_,
  r_n_182__30_,r_n_182__29_,r_n_182__28_,r_n_182__27_,r_n_182__26_,r_n_182__25_,
  r_n_182__24_,r_n_182__23_,r_n_182__22_,r_n_182__21_,r_n_182__20_,r_n_182__19_,r_n_182__18_,
  r_n_182__17_,r_n_182__16_,r_n_182__15_,r_n_182__14_,r_n_182__13_,r_n_182__12_,
  r_n_182__11_,r_n_182__10_,r_n_182__9_,r_n_182__8_,r_n_182__7_,r_n_182__6_,
  r_n_182__5_,r_n_182__4_,r_n_182__3_,r_n_182__2_,r_n_182__1_,r_n_182__0_,r_n_181__63_,
  r_n_181__62_,r_n_181__61_,r_n_181__60_,r_n_181__59_,r_n_181__58_,r_n_181__57_,
  r_n_181__56_,r_n_181__55_,r_n_181__54_,r_n_181__53_,r_n_181__52_,r_n_181__51_,
  r_n_181__50_,r_n_181__49_,r_n_181__48_,r_n_181__47_,r_n_181__46_,r_n_181__45_,
  r_n_181__44_,r_n_181__43_,r_n_181__42_,r_n_181__41_,r_n_181__40_,r_n_181__39_,
  r_n_181__38_,r_n_181__37_,r_n_181__36_,r_n_181__35_,r_n_181__34_,r_n_181__33_,r_n_181__32_,
  r_n_181__31_,r_n_181__30_,r_n_181__29_,r_n_181__28_,r_n_181__27_,r_n_181__26_,
  r_n_181__25_,r_n_181__24_,r_n_181__23_,r_n_181__22_,r_n_181__21_,r_n_181__20_,
  r_n_181__19_,r_n_181__18_,r_n_181__17_,r_n_181__16_,r_n_181__15_,r_n_181__14_,
  r_n_181__13_,r_n_181__12_,r_n_181__11_,r_n_181__10_,r_n_181__9_,r_n_181__8_,
  r_n_181__7_,r_n_181__6_,r_n_181__5_,r_n_181__4_,r_n_181__3_,r_n_181__2_,r_n_181__1_,
  r_n_181__0_,r_n_180__63_,r_n_180__62_,r_n_180__61_,r_n_180__60_,r_n_180__59_,
  r_n_180__58_,r_n_180__57_,r_n_180__56_,r_n_180__55_,r_n_180__54_,r_n_180__53_,
  r_n_180__52_,r_n_180__51_,r_n_180__50_,r_n_180__49_,r_n_180__48_,r_n_180__47_,r_n_180__46_,
  r_n_180__45_,r_n_180__44_,r_n_180__43_,r_n_180__42_,r_n_180__41_,r_n_180__40_,
  r_n_180__39_,r_n_180__38_,r_n_180__37_,r_n_180__36_,r_n_180__35_,r_n_180__34_,
  r_n_180__33_,r_n_180__32_,r_n_180__31_,r_n_180__30_,r_n_180__29_,r_n_180__28_,
  r_n_180__27_,r_n_180__26_,r_n_180__25_,r_n_180__24_,r_n_180__23_,r_n_180__22_,
  r_n_180__21_,r_n_180__20_,r_n_180__19_,r_n_180__18_,r_n_180__17_,r_n_180__16_,
  r_n_180__15_,r_n_180__14_,r_n_180__13_,r_n_180__12_,r_n_180__11_,r_n_180__10_,r_n_180__9_,
  r_n_180__8_,r_n_180__7_,r_n_180__6_,r_n_180__5_,r_n_180__4_,r_n_180__3_,
  r_n_180__2_,r_n_180__1_,r_n_180__0_,r_n_179__63_,r_n_179__62_,r_n_179__61_,r_n_179__60_,
  r_n_179__59_,r_n_179__58_,r_n_179__57_,r_n_179__56_,r_n_179__55_,r_n_179__54_,
  r_n_179__53_,r_n_179__52_,r_n_179__51_,r_n_179__50_,r_n_179__49_,r_n_179__48_,
  r_n_179__47_,r_n_179__46_,r_n_179__45_,r_n_179__44_,r_n_179__43_,r_n_179__42_,
  r_n_179__41_,r_n_179__40_,r_n_179__39_,r_n_179__38_,r_n_179__37_,r_n_179__36_,
  r_n_179__35_,r_n_179__34_,r_n_179__33_,r_n_179__32_,r_n_179__31_,r_n_179__30_,
  r_n_179__29_,r_n_179__28_,r_n_179__27_,r_n_179__26_,r_n_179__25_,r_n_179__24_,
  r_n_179__23_,r_n_179__22_,r_n_179__21_,r_n_179__20_,r_n_179__19_,r_n_179__18_,r_n_179__17_,
  r_n_179__16_,r_n_179__15_,r_n_179__14_,r_n_179__13_,r_n_179__12_,r_n_179__11_,
  r_n_179__10_,r_n_179__9_,r_n_179__8_,r_n_179__7_,r_n_179__6_,r_n_179__5_,
  r_n_179__4_,r_n_179__3_,r_n_179__2_,r_n_179__1_,r_n_179__0_,r_n_178__63_,r_n_178__62_,
  r_n_178__61_,r_n_178__60_,r_n_178__59_,r_n_178__58_,r_n_178__57_,r_n_178__56_,
  r_n_178__55_,r_n_178__54_,r_n_178__53_,r_n_178__52_,r_n_178__51_,r_n_178__50_,
  r_n_178__49_,r_n_178__48_,r_n_178__47_,r_n_178__46_,r_n_178__45_,r_n_178__44_,
  r_n_178__43_,r_n_178__42_,r_n_178__41_,r_n_178__40_,r_n_178__39_,r_n_178__38_,
  r_n_178__37_,r_n_178__36_,r_n_178__35_,r_n_178__34_,r_n_178__33_,r_n_178__32_,r_n_178__31_,
  r_n_178__30_,r_n_178__29_,r_n_178__28_,r_n_178__27_,r_n_178__26_,r_n_178__25_,
  r_n_178__24_,r_n_178__23_,r_n_178__22_,r_n_178__21_,r_n_178__20_,r_n_178__19_,
  r_n_178__18_,r_n_178__17_,r_n_178__16_,r_n_178__15_,r_n_178__14_,r_n_178__13_,
  r_n_178__12_,r_n_178__11_,r_n_178__10_,r_n_178__9_,r_n_178__8_,r_n_178__7_,r_n_178__6_,
  r_n_178__5_,r_n_178__4_,r_n_178__3_,r_n_178__2_,r_n_178__1_,r_n_178__0_,
  r_n_177__63_,r_n_177__62_,r_n_177__61_,r_n_177__60_,r_n_177__59_,r_n_177__58_,
  r_n_177__57_,r_n_177__56_,r_n_177__55_,r_n_177__54_,r_n_177__53_,r_n_177__52_,
  r_n_177__51_,r_n_177__50_,r_n_177__49_,r_n_177__48_,r_n_177__47_,r_n_177__46_,r_n_177__45_,
  r_n_177__44_,r_n_177__43_,r_n_177__42_,r_n_177__41_,r_n_177__40_,r_n_177__39_,
  r_n_177__38_,r_n_177__37_,r_n_177__36_,r_n_177__35_,r_n_177__34_,r_n_177__33_,
  r_n_177__32_,r_n_177__31_,r_n_177__30_,r_n_177__29_,r_n_177__28_,r_n_177__27_,
  r_n_177__26_,r_n_177__25_,r_n_177__24_,r_n_177__23_,r_n_177__22_,r_n_177__21_,
  r_n_177__20_,r_n_177__19_,r_n_177__18_,r_n_177__17_,r_n_177__16_,r_n_177__15_,
  r_n_177__14_,r_n_177__13_,r_n_177__12_,r_n_177__11_,r_n_177__10_,r_n_177__9_,r_n_177__8_,
  r_n_177__7_,r_n_177__6_,r_n_177__5_,r_n_177__4_,r_n_177__3_,r_n_177__2_,
  r_n_177__1_,r_n_177__0_,r_n_192__63_,r_n_192__62_,r_n_192__61_,r_n_192__60_,r_n_192__59_,
  r_n_192__58_,r_n_192__57_,r_n_192__56_,r_n_192__55_,r_n_192__54_,r_n_192__53_,
  r_n_192__52_,r_n_192__51_,r_n_192__50_,r_n_192__49_,r_n_192__48_,r_n_192__47_,
  r_n_192__46_,r_n_192__45_,r_n_192__44_,r_n_192__43_,r_n_192__42_,r_n_192__41_,
  r_n_192__40_,r_n_192__39_,r_n_192__38_,r_n_192__37_,r_n_192__36_,r_n_192__35_,
  r_n_192__34_,r_n_192__33_,r_n_192__32_,r_n_192__31_,r_n_192__30_,r_n_192__29_,
  r_n_192__28_,r_n_192__27_,r_n_192__26_,r_n_192__25_,r_n_192__24_,r_n_192__23_,r_n_192__22_,
  r_n_192__21_,r_n_192__20_,r_n_192__19_,r_n_192__18_,r_n_192__17_,r_n_192__16_,
  r_n_192__15_,r_n_192__14_,r_n_192__13_,r_n_192__12_,r_n_192__11_,r_n_192__10_,
  r_n_192__9_,r_n_192__8_,r_n_192__7_,r_n_192__6_,r_n_192__5_,r_n_192__4_,r_n_192__3_,
  r_n_192__2_,r_n_192__1_,r_n_192__0_,r_n_191__63_,r_n_191__62_,r_n_191__61_,
  r_n_191__60_,r_n_191__59_,r_n_191__58_,r_n_191__57_,r_n_191__56_,r_n_191__55_,
  r_n_191__54_,r_n_191__53_,r_n_191__52_,r_n_191__51_,r_n_191__50_,r_n_191__49_,
  r_n_191__48_,r_n_191__47_,r_n_191__46_,r_n_191__45_,r_n_191__44_,r_n_191__43_,
  r_n_191__42_,r_n_191__41_,r_n_191__40_,r_n_191__39_,r_n_191__38_,r_n_191__37_,r_n_191__36_,
  r_n_191__35_,r_n_191__34_,r_n_191__33_,r_n_191__32_,r_n_191__31_,r_n_191__30_,
  r_n_191__29_,r_n_191__28_,r_n_191__27_,r_n_191__26_,r_n_191__25_,r_n_191__24_,
  r_n_191__23_,r_n_191__22_,r_n_191__21_,r_n_191__20_,r_n_191__19_,r_n_191__18_,
  r_n_191__17_,r_n_191__16_,r_n_191__15_,r_n_191__14_,r_n_191__13_,r_n_191__12_,
  r_n_191__11_,r_n_191__10_,r_n_191__9_,r_n_191__8_,r_n_191__7_,r_n_191__6_,r_n_191__5_,
  r_n_191__4_,r_n_191__3_,r_n_191__2_,r_n_191__1_,r_n_191__0_,r_n_190__63_,
  r_n_190__62_,r_n_190__61_,r_n_190__60_,r_n_190__59_,r_n_190__58_,r_n_190__57_,
  r_n_190__56_,r_n_190__55_,r_n_190__54_,r_n_190__53_,r_n_190__52_,r_n_190__51_,r_n_190__50_,
  r_n_190__49_,r_n_190__48_,r_n_190__47_,r_n_190__46_,r_n_190__45_,r_n_190__44_,
  r_n_190__43_,r_n_190__42_,r_n_190__41_,r_n_190__40_,r_n_190__39_,r_n_190__38_,
  r_n_190__37_,r_n_190__36_,r_n_190__35_,r_n_190__34_,r_n_190__33_,r_n_190__32_,
  r_n_190__31_,r_n_190__30_,r_n_190__29_,r_n_190__28_,r_n_190__27_,r_n_190__26_,
  r_n_190__25_,r_n_190__24_,r_n_190__23_,r_n_190__22_,r_n_190__21_,r_n_190__20_,
  r_n_190__19_,r_n_190__18_,r_n_190__17_,r_n_190__16_,r_n_190__15_,r_n_190__14_,
  r_n_190__13_,r_n_190__12_,r_n_190__11_,r_n_190__10_,r_n_190__9_,r_n_190__8_,r_n_190__7_,
  r_n_190__6_,r_n_190__5_,r_n_190__4_,r_n_190__3_,r_n_190__2_,r_n_190__1_,r_n_190__0_,
  r_n_189__63_,r_n_189__62_,r_n_189__61_,r_n_189__60_,r_n_189__59_,r_n_189__58_,
  r_n_189__57_,r_n_189__56_,r_n_189__55_,r_n_189__54_,r_n_189__53_,r_n_189__52_,
  r_n_189__51_,r_n_189__50_,r_n_189__49_,r_n_189__48_,r_n_189__47_,r_n_189__46_,
  r_n_189__45_,r_n_189__44_,r_n_189__43_,r_n_189__42_,r_n_189__41_,r_n_189__40_,
  r_n_189__39_,r_n_189__38_,r_n_189__37_,r_n_189__36_,r_n_189__35_,r_n_189__34_,
  r_n_189__33_,r_n_189__32_,r_n_189__31_,r_n_189__30_,r_n_189__29_,r_n_189__28_,
  r_n_189__27_,r_n_189__26_,r_n_189__25_,r_n_189__24_,r_n_189__23_,r_n_189__22_,r_n_189__21_,
  r_n_189__20_,r_n_189__19_,r_n_189__18_,r_n_189__17_,r_n_189__16_,r_n_189__15_,
  r_n_189__14_,r_n_189__13_,r_n_189__12_,r_n_189__11_,r_n_189__10_,r_n_189__9_,
  r_n_189__8_,r_n_189__7_,r_n_189__6_,r_n_189__5_,r_n_189__4_,r_n_189__3_,r_n_189__2_,
  r_n_189__1_,r_n_189__0_,r_n_188__63_,r_n_188__62_,r_n_188__61_,r_n_188__60_,
  r_n_188__59_,r_n_188__58_,r_n_188__57_,r_n_188__56_,r_n_188__55_,r_n_188__54_,
  r_n_188__53_,r_n_188__52_,r_n_188__51_,r_n_188__50_,r_n_188__49_,r_n_188__48_,
  r_n_188__47_,r_n_188__46_,r_n_188__45_,r_n_188__44_,r_n_188__43_,r_n_188__42_,
  r_n_188__41_,r_n_188__40_,r_n_188__39_,r_n_188__38_,r_n_188__37_,r_n_188__36_,r_n_188__35_,
  r_n_188__34_,r_n_188__33_,r_n_188__32_,r_n_188__31_,r_n_188__30_,r_n_188__29_,
  r_n_188__28_,r_n_188__27_,r_n_188__26_,r_n_188__25_,r_n_188__24_,r_n_188__23_,
  r_n_188__22_,r_n_188__21_,r_n_188__20_,r_n_188__19_,r_n_188__18_,r_n_188__17_,
  r_n_188__16_,r_n_188__15_,r_n_188__14_,r_n_188__13_,r_n_188__12_,r_n_188__11_,
  r_n_188__10_,r_n_188__9_,r_n_188__8_,r_n_188__7_,r_n_188__6_,r_n_188__5_,r_n_188__4_,
  r_n_188__3_,r_n_188__2_,r_n_188__1_,r_n_188__0_,r_n_187__63_,r_n_187__62_,
  r_n_187__61_,r_n_187__60_,r_n_187__59_,r_n_187__58_,r_n_187__57_,r_n_187__56_,
  r_n_187__55_,r_n_187__54_,r_n_187__53_,r_n_187__52_,r_n_187__51_,r_n_187__50_,r_n_187__49_,
  r_n_187__48_,r_n_187__47_,r_n_187__46_,r_n_187__45_,r_n_187__44_,r_n_187__43_,
  r_n_187__42_,r_n_187__41_,r_n_187__40_,r_n_187__39_,r_n_187__38_,r_n_187__37_,
  r_n_187__36_,r_n_187__35_,r_n_187__34_,r_n_187__33_,r_n_187__32_,r_n_187__31_,
  r_n_187__30_,r_n_187__29_,r_n_187__28_,r_n_187__27_,r_n_187__26_,r_n_187__25_,
  r_n_187__24_,r_n_187__23_,r_n_187__22_,r_n_187__21_,r_n_187__20_,r_n_187__19_,
  r_n_187__18_,r_n_187__17_,r_n_187__16_,r_n_187__15_,r_n_187__14_,r_n_187__13_,r_n_187__12_,
  r_n_187__11_,r_n_187__10_,r_n_187__9_,r_n_187__8_,r_n_187__7_,r_n_187__6_,
  r_n_187__5_,r_n_187__4_,r_n_187__3_,r_n_187__2_,r_n_187__1_,r_n_187__0_,r_n_186__63_,
  r_n_186__62_,r_n_186__61_,r_n_186__60_,r_n_186__59_,r_n_186__58_,r_n_186__57_,
  r_n_186__56_,r_n_186__55_,r_n_186__54_,r_n_186__53_,r_n_186__52_,r_n_186__51_,
  r_n_186__50_,r_n_186__49_,r_n_186__48_,r_n_186__47_,r_n_186__46_,r_n_186__45_,
  r_n_186__44_,r_n_186__43_,r_n_186__42_,r_n_186__41_,r_n_186__40_,r_n_186__39_,
  r_n_186__38_,r_n_186__37_,r_n_186__36_,r_n_186__35_,r_n_186__34_,r_n_186__33_,
  r_n_186__32_,r_n_186__31_,r_n_186__30_,r_n_186__29_,r_n_186__28_,r_n_186__27_,r_n_186__26_,
  r_n_186__25_,r_n_186__24_,r_n_186__23_,r_n_186__22_,r_n_186__21_,r_n_186__20_,
  r_n_186__19_,r_n_186__18_,r_n_186__17_,r_n_186__16_,r_n_186__15_,r_n_186__14_,
  r_n_186__13_,r_n_186__12_,r_n_186__11_,r_n_186__10_,r_n_186__9_,r_n_186__8_,
  r_n_186__7_,r_n_186__6_,r_n_186__5_,r_n_186__4_,r_n_186__3_,r_n_186__2_,r_n_186__1_,
  r_n_186__0_,r_n_185__63_,r_n_185__62_,r_n_185__61_,r_n_185__60_,r_n_185__59_,
  r_n_185__58_,r_n_185__57_,r_n_185__56_,r_n_185__55_,r_n_185__54_,r_n_185__53_,
  r_n_185__52_,r_n_185__51_,r_n_185__50_,r_n_185__49_,r_n_185__48_,r_n_185__47_,
  r_n_185__46_,r_n_185__45_,r_n_185__44_,r_n_185__43_,r_n_185__42_,r_n_185__41_,r_n_185__40_,
  r_n_185__39_,r_n_185__38_,r_n_185__37_,r_n_185__36_,r_n_185__35_,r_n_185__34_,
  r_n_185__33_,r_n_185__32_,r_n_185__31_,r_n_185__30_,r_n_185__29_,r_n_185__28_,
  r_n_185__27_,r_n_185__26_,r_n_185__25_,r_n_185__24_,r_n_185__23_,r_n_185__22_,
  r_n_185__21_,r_n_185__20_,r_n_185__19_,r_n_185__18_,r_n_185__17_,r_n_185__16_,
  r_n_185__15_,r_n_185__14_,r_n_185__13_,r_n_185__12_,r_n_185__11_,r_n_185__10_,
  r_n_185__9_,r_n_185__8_,r_n_185__7_,r_n_185__6_,r_n_185__5_,r_n_185__4_,r_n_185__3_,
  r_n_185__2_,r_n_185__1_,r_n_185__0_,r_n_200__63_,r_n_200__62_,r_n_200__61_,
  r_n_200__60_,r_n_200__59_,r_n_200__58_,r_n_200__57_,r_n_200__56_,r_n_200__55_,r_n_200__54_,
  r_n_200__53_,r_n_200__52_,r_n_200__51_,r_n_200__50_,r_n_200__49_,r_n_200__48_,
  r_n_200__47_,r_n_200__46_,r_n_200__45_,r_n_200__44_,r_n_200__43_,r_n_200__42_,
  r_n_200__41_,r_n_200__40_,r_n_200__39_,r_n_200__38_,r_n_200__37_,r_n_200__36_,
  r_n_200__35_,r_n_200__34_,r_n_200__33_,r_n_200__32_,r_n_200__31_,r_n_200__30_,
  r_n_200__29_,r_n_200__28_,r_n_200__27_,r_n_200__26_,r_n_200__25_,r_n_200__24_,
  r_n_200__23_,r_n_200__22_,r_n_200__21_,r_n_200__20_,r_n_200__19_,r_n_200__18_,
  r_n_200__17_,r_n_200__16_,r_n_200__15_,r_n_200__14_,r_n_200__13_,r_n_200__12_,r_n_200__11_,
  r_n_200__10_,r_n_200__9_,r_n_200__8_,r_n_200__7_,r_n_200__6_,r_n_200__5_,
  r_n_200__4_,r_n_200__3_,r_n_200__2_,r_n_200__1_,r_n_200__0_,r_n_199__63_,r_n_199__62_,
  r_n_199__61_,r_n_199__60_,r_n_199__59_,r_n_199__58_,r_n_199__57_,r_n_199__56_,
  r_n_199__55_,r_n_199__54_,r_n_199__53_,r_n_199__52_,r_n_199__51_,r_n_199__50_,
  r_n_199__49_,r_n_199__48_,r_n_199__47_,r_n_199__46_,r_n_199__45_,r_n_199__44_,
  r_n_199__43_,r_n_199__42_,r_n_199__41_,r_n_199__40_,r_n_199__39_,r_n_199__38_,
  r_n_199__37_,r_n_199__36_,r_n_199__35_,r_n_199__34_,r_n_199__33_,r_n_199__32_,
  r_n_199__31_,r_n_199__30_,r_n_199__29_,r_n_199__28_,r_n_199__27_,r_n_199__26_,r_n_199__25_,
  r_n_199__24_,r_n_199__23_,r_n_199__22_,r_n_199__21_,r_n_199__20_,r_n_199__19_,
  r_n_199__18_,r_n_199__17_,r_n_199__16_,r_n_199__15_,r_n_199__14_,r_n_199__13_,
  r_n_199__12_,r_n_199__11_,r_n_199__10_,r_n_199__9_,r_n_199__8_,r_n_199__7_,
  r_n_199__6_,r_n_199__5_,r_n_199__4_,r_n_199__3_,r_n_199__2_,r_n_199__1_,r_n_199__0_,
  r_n_198__63_,r_n_198__62_,r_n_198__61_,r_n_198__60_,r_n_198__59_,r_n_198__58_,
  r_n_198__57_,r_n_198__56_,r_n_198__55_,r_n_198__54_,r_n_198__53_,r_n_198__52_,
  r_n_198__51_,r_n_198__50_,r_n_198__49_,r_n_198__48_,r_n_198__47_,r_n_198__46_,
  r_n_198__45_,r_n_198__44_,r_n_198__43_,r_n_198__42_,r_n_198__41_,r_n_198__40_,r_n_198__39_,
  r_n_198__38_,r_n_198__37_,r_n_198__36_,r_n_198__35_,r_n_198__34_,r_n_198__33_,
  r_n_198__32_,r_n_198__31_,r_n_198__30_,r_n_198__29_,r_n_198__28_,r_n_198__27_,
  r_n_198__26_,r_n_198__25_,r_n_198__24_,r_n_198__23_,r_n_198__22_,r_n_198__21_,
  r_n_198__20_,r_n_198__19_,r_n_198__18_,r_n_198__17_,r_n_198__16_,r_n_198__15_,
  r_n_198__14_,r_n_198__13_,r_n_198__12_,r_n_198__11_,r_n_198__10_,r_n_198__9_,r_n_198__8_,
  r_n_198__7_,r_n_198__6_,r_n_198__5_,r_n_198__4_,r_n_198__3_,r_n_198__2_,
  r_n_198__1_,r_n_198__0_,r_n_197__63_,r_n_197__62_,r_n_197__61_,r_n_197__60_,
  r_n_197__59_,r_n_197__58_,r_n_197__57_,r_n_197__56_,r_n_197__55_,r_n_197__54_,r_n_197__53_,
  r_n_197__52_,r_n_197__51_,r_n_197__50_,r_n_197__49_,r_n_197__48_,r_n_197__47_,
  r_n_197__46_,r_n_197__45_,r_n_197__44_,r_n_197__43_,r_n_197__42_,r_n_197__41_,
  r_n_197__40_,r_n_197__39_,r_n_197__38_,r_n_197__37_,r_n_197__36_,r_n_197__35_,
  r_n_197__34_,r_n_197__33_,r_n_197__32_,r_n_197__31_,r_n_197__30_,r_n_197__29_,
  r_n_197__28_,r_n_197__27_,r_n_197__26_,r_n_197__25_,r_n_197__24_,r_n_197__23_,
  r_n_197__22_,r_n_197__21_,r_n_197__20_,r_n_197__19_,r_n_197__18_,r_n_197__17_,r_n_197__16_,
  r_n_197__15_,r_n_197__14_,r_n_197__13_,r_n_197__12_,r_n_197__11_,r_n_197__10_,
  r_n_197__9_,r_n_197__8_,r_n_197__7_,r_n_197__6_,r_n_197__5_,r_n_197__4_,
  r_n_197__3_,r_n_197__2_,r_n_197__1_,r_n_197__0_,r_n_196__63_,r_n_196__62_,r_n_196__61_,
  r_n_196__60_,r_n_196__59_,r_n_196__58_,r_n_196__57_,r_n_196__56_,r_n_196__55_,
  r_n_196__54_,r_n_196__53_,r_n_196__52_,r_n_196__51_,r_n_196__50_,r_n_196__49_,
  r_n_196__48_,r_n_196__47_,r_n_196__46_,r_n_196__45_,r_n_196__44_,r_n_196__43_,
  r_n_196__42_,r_n_196__41_,r_n_196__40_,r_n_196__39_,r_n_196__38_,r_n_196__37_,
  r_n_196__36_,r_n_196__35_,r_n_196__34_,r_n_196__33_,r_n_196__32_,r_n_196__31_,r_n_196__30_,
  r_n_196__29_,r_n_196__28_,r_n_196__27_,r_n_196__26_,r_n_196__25_,r_n_196__24_,
  r_n_196__23_,r_n_196__22_,r_n_196__21_,r_n_196__20_,r_n_196__19_,r_n_196__18_,
  r_n_196__17_,r_n_196__16_,r_n_196__15_,r_n_196__14_,r_n_196__13_,r_n_196__12_,
  r_n_196__11_,r_n_196__10_,r_n_196__9_,r_n_196__8_,r_n_196__7_,r_n_196__6_,r_n_196__5_,
  r_n_196__4_,r_n_196__3_,r_n_196__2_,r_n_196__1_,r_n_196__0_,r_n_195__63_,
  r_n_195__62_,r_n_195__61_,r_n_195__60_,r_n_195__59_,r_n_195__58_,r_n_195__57_,
  r_n_195__56_,r_n_195__55_,r_n_195__54_,r_n_195__53_,r_n_195__52_,r_n_195__51_,
  r_n_195__50_,r_n_195__49_,r_n_195__48_,r_n_195__47_,r_n_195__46_,r_n_195__45_,r_n_195__44_,
  r_n_195__43_,r_n_195__42_,r_n_195__41_,r_n_195__40_,r_n_195__39_,r_n_195__38_,
  r_n_195__37_,r_n_195__36_,r_n_195__35_,r_n_195__34_,r_n_195__33_,r_n_195__32_,
  r_n_195__31_,r_n_195__30_,r_n_195__29_,r_n_195__28_,r_n_195__27_,r_n_195__26_,
  r_n_195__25_,r_n_195__24_,r_n_195__23_,r_n_195__22_,r_n_195__21_,r_n_195__20_,
  r_n_195__19_,r_n_195__18_,r_n_195__17_,r_n_195__16_,r_n_195__15_,r_n_195__14_,
  r_n_195__13_,r_n_195__12_,r_n_195__11_,r_n_195__10_,r_n_195__9_,r_n_195__8_,r_n_195__7_,
  r_n_195__6_,r_n_195__5_,r_n_195__4_,r_n_195__3_,r_n_195__2_,r_n_195__1_,
  r_n_195__0_,r_n_194__63_,r_n_194__62_,r_n_194__61_,r_n_194__60_,r_n_194__59_,r_n_194__58_,
  r_n_194__57_,r_n_194__56_,r_n_194__55_,r_n_194__54_,r_n_194__53_,r_n_194__52_,
  r_n_194__51_,r_n_194__50_,r_n_194__49_,r_n_194__48_,r_n_194__47_,r_n_194__46_,
  r_n_194__45_,r_n_194__44_,r_n_194__43_,r_n_194__42_,r_n_194__41_,r_n_194__40_,
  r_n_194__39_,r_n_194__38_,r_n_194__37_,r_n_194__36_,r_n_194__35_,r_n_194__34_,
  r_n_194__33_,r_n_194__32_,r_n_194__31_,r_n_194__30_,r_n_194__29_,r_n_194__28_,
  r_n_194__27_,r_n_194__26_,r_n_194__25_,r_n_194__24_,r_n_194__23_,r_n_194__22_,
  r_n_194__21_,r_n_194__20_,r_n_194__19_,r_n_194__18_,r_n_194__17_,r_n_194__16_,r_n_194__15_,
  r_n_194__14_,r_n_194__13_,r_n_194__12_,r_n_194__11_,r_n_194__10_,r_n_194__9_,
  r_n_194__8_,r_n_194__7_,r_n_194__6_,r_n_194__5_,r_n_194__4_,r_n_194__3_,r_n_194__2_,
  r_n_194__1_,r_n_194__0_,r_n_193__63_,r_n_193__62_,r_n_193__61_,r_n_193__60_,
  r_n_193__59_,r_n_193__58_,r_n_193__57_,r_n_193__56_,r_n_193__55_,r_n_193__54_,
  r_n_193__53_,r_n_193__52_,r_n_193__51_,r_n_193__50_,r_n_193__49_,r_n_193__48_,
  r_n_193__47_,r_n_193__46_,r_n_193__45_,r_n_193__44_,r_n_193__43_,r_n_193__42_,
  r_n_193__41_,r_n_193__40_,r_n_193__39_,r_n_193__38_,r_n_193__37_,r_n_193__36_,
  r_n_193__35_,r_n_193__34_,r_n_193__33_,r_n_193__32_,r_n_193__31_,r_n_193__30_,r_n_193__29_,
  r_n_193__28_,r_n_193__27_,r_n_193__26_,r_n_193__25_,r_n_193__24_,r_n_193__23_,
  r_n_193__22_,r_n_193__21_,r_n_193__20_,r_n_193__19_,r_n_193__18_,r_n_193__17_,
  r_n_193__16_,r_n_193__15_,r_n_193__14_,r_n_193__13_,r_n_193__12_,r_n_193__11_,
  r_n_193__10_,r_n_193__9_,r_n_193__8_,r_n_193__7_,r_n_193__6_,r_n_193__5_,r_n_193__4_,
  r_n_193__3_,r_n_193__2_,r_n_193__1_,r_n_193__0_,r_n_208__63_,r_n_208__62_,
  r_n_208__61_,r_n_208__60_,r_n_208__59_,r_n_208__58_,r_n_208__57_,r_n_208__56_,
  r_n_208__55_,r_n_208__54_,r_n_208__53_,r_n_208__52_,r_n_208__51_,r_n_208__50_,
  r_n_208__49_,r_n_208__48_,r_n_208__47_,r_n_208__46_,r_n_208__45_,r_n_208__44_,r_n_208__43_,
  r_n_208__42_,r_n_208__41_,r_n_208__40_,r_n_208__39_,r_n_208__38_,r_n_208__37_,
  r_n_208__36_,r_n_208__35_,r_n_208__34_,r_n_208__33_,r_n_208__32_,r_n_208__31_,
  r_n_208__30_,r_n_208__29_,r_n_208__28_,r_n_208__27_,r_n_208__26_,r_n_208__25_,
  r_n_208__24_,r_n_208__23_,r_n_208__22_,r_n_208__21_,r_n_208__20_,r_n_208__19_,
  r_n_208__18_,r_n_208__17_,r_n_208__16_,r_n_208__15_,r_n_208__14_,r_n_208__13_,
  r_n_208__12_,r_n_208__11_,r_n_208__10_,r_n_208__9_,r_n_208__8_,r_n_208__7_,r_n_208__6_,
  r_n_208__5_,r_n_208__4_,r_n_208__3_,r_n_208__2_,r_n_208__1_,r_n_208__0_,
  r_n_207__63_,r_n_207__62_,r_n_207__61_,r_n_207__60_,r_n_207__59_,r_n_207__58_,r_n_207__57_,
  r_n_207__56_,r_n_207__55_,r_n_207__54_,r_n_207__53_,r_n_207__52_,r_n_207__51_,
  r_n_207__50_,r_n_207__49_,r_n_207__48_,r_n_207__47_,r_n_207__46_,r_n_207__45_,
  r_n_207__44_,r_n_207__43_,r_n_207__42_,r_n_207__41_,r_n_207__40_,r_n_207__39_,
  r_n_207__38_,r_n_207__37_,r_n_207__36_,r_n_207__35_,r_n_207__34_,r_n_207__33_,
  r_n_207__32_,r_n_207__31_,r_n_207__30_,r_n_207__29_,r_n_207__28_,r_n_207__27_,
  r_n_207__26_,r_n_207__25_,r_n_207__24_,r_n_207__23_,r_n_207__22_,r_n_207__21_,r_n_207__20_,
  r_n_207__19_,r_n_207__18_,r_n_207__17_,r_n_207__16_,r_n_207__15_,r_n_207__14_,
  r_n_207__13_,r_n_207__12_,r_n_207__11_,r_n_207__10_,r_n_207__9_,r_n_207__8_,
  r_n_207__7_,r_n_207__6_,r_n_207__5_,r_n_207__4_,r_n_207__3_,r_n_207__2_,r_n_207__1_,
  r_n_207__0_,r_n_206__63_,r_n_206__62_,r_n_206__61_,r_n_206__60_,r_n_206__59_,
  r_n_206__58_,r_n_206__57_,r_n_206__56_,r_n_206__55_,r_n_206__54_,r_n_206__53_,
  r_n_206__52_,r_n_206__51_,r_n_206__50_,r_n_206__49_,r_n_206__48_,r_n_206__47_,
  r_n_206__46_,r_n_206__45_,r_n_206__44_,r_n_206__43_,r_n_206__42_,r_n_206__41_,
  r_n_206__40_,r_n_206__39_,r_n_206__38_,r_n_206__37_,r_n_206__36_,r_n_206__35_,r_n_206__34_,
  r_n_206__33_,r_n_206__32_,r_n_206__31_,r_n_206__30_,r_n_206__29_,r_n_206__28_,
  r_n_206__27_,r_n_206__26_,r_n_206__25_,r_n_206__24_,r_n_206__23_,r_n_206__22_,
  r_n_206__21_,r_n_206__20_,r_n_206__19_,r_n_206__18_,r_n_206__17_,r_n_206__16_,
  r_n_206__15_,r_n_206__14_,r_n_206__13_,r_n_206__12_,r_n_206__11_,r_n_206__10_,
  r_n_206__9_,r_n_206__8_,r_n_206__7_,r_n_206__6_,r_n_206__5_,r_n_206__4_,r_n_206__3_,
  r_n_206__2_,r_n_206__1_,r_n_206__0_,r_n_205__63_,r_n_205__62_,r_n_205__61_,
  r_n_205__60_,r_n_205__59_,r_n_205__58_,r_n_205__57_,r_n_205__56_,r_n_205__55_,
  r_n_205__54_,r_n_205__53_,r_n_205__52_,r_n_205__51_,r_n_205__50_,r_n_205__49_,r_n_205__48_,
  r_n_205__47_,r_n_205__46_,r_n_205__45_,r_n_205__44_,r_n_205__43_,r_n_205__42_,
  r_n_205__41_,r_n_205__40_,r_n_205__39_,r_n_205__38_,r_n_205__37_,r_n_205__36_,
  r_n_205__35_,r_n_205__34_,r_n_205__33_,r_n_205__32_,r_n_205__31_,r_n_205__30_,
  r_n_205__29_,r_n_205__28_,r_n_205__27_,r_n_205__26_,r_n_205__25_,r_n_205__24_,
  r_n_205__23_,r_n_205__22_,r_n_205__21_,r_n_205__20_,r_n_205__19_,r_n_205__18_,
  r_n_205__17_,r_n_205__16_,r_n_205__15_,r_n_205__14_,r_n_205__13_,r_n_205__12_,
  r_n_205__11_,r_n_205__10_,r_n_205__9_,r_n_205__8_,r_n_205__7_,r_n_205__6_,r_n_205__5_,
  r_n_205__4_,r_n_205__3_,r_n_205__2_,r_n_205__1_,r_n_205__0_,r_n_204__63_,r_n_204__62_,
  r_n_204__61_,r_n_204__60_,r_n_204__59_,r_n_204__58_,r_n_204__57_,r_n_204__56_,
  r_n_204__55_,r_n_204__54_,r_n_204__53_,r_n_204__52_,r_n_204__51_,r_n_204__50_,
  r_n_204__49_,r_n_204__48_,r_n_204__47_,r_n_204__46_,r_n_204__45_,r_n_204__44_,
  r_n_204__43_,r_n_204__42_,r_n_204__41_,r_n_204__40_,r_n_204__39_,r_n_204__38_,
  r_n_204__37_,r_n_204__36_,r_n_204__35_,r_n_204__34_,r_n_204__33_,r_n_204__32_,
  r_n_204__31_,r_n_204__30_,r_n_204__29_,r_n_204__28_,r_n_204__27_,r_n_204__26_,
  r_n_204__25_,r_n_204__24_,r_n_204__23_,r_n_204__22_,r_n_204__21_,r_n_204__20_,r_n_204__19_,
  r_n_204__18_,r_n_204__17_,r_n_204__16_,r_n_204__15_,r_n_204__14_,r_n_204__13_,
  r_n_204__12_,r_n_204__11_,r_n_204__10_,r_n_204__9_,r_n_204__8_,r_n_204__7_,
  r_n_204__6_,r_n_204__5_,r_n_204__4_,r_n_204__3_,r_n_204__2_,r_n_204__1_,r_n_204__0_,
  r_n_203__63_,r_n_203__62_,r_n_203__61_,r_n_203__60_,r_n_203__59_,r_n_203__58_,
  r_n_203__57_,r_n_203__56_,r_n_203__55_,r_n_203__54_,r_n_203__53_,r_n_203__52_,
  r_n_203__51_,r_n_203__50_,r_n_203__49_,r_n_203__48_,r_n_203__47_,r_n_203__46_,
  r_n_203__45_,r_n_203__44_,r_n_203__43_,r_n_203__42_,r_n_203__41_,r_n_203__40_,
  r_n_203__39_,r_n_203__38_,r_n_203__37_,r_n_203__36_,r_n_203__35_,r_n_203__34_,r_n_203__33_,
  r_n_203__32_,r_n_203__31_,r_n_203__30_,r_n_203__29_,r_n_203__28_,r_n_203__27_,
  r_n_203__26_,r_n_203__25_,r_n_203__24_,r_n_203__23_,r_n_203__22_,r_n_203__21_,
  r_n_203__20_,r_n_203__19_,r_n_203__18_,r_n_203__17_,r_n_203__16_,r_n_203__15_,
  r_n_203__14_,r_n_203__13_,r_n_203__12_,r_n_203__11_,r_n_203__10_,r_n_203__9_,
  r_n_203__8_,r_n_203__7_,r_n_203__6_,r_n_203__5_,r_n_203__4_,r_n_203__3_,r_n_203__2_,
  r_n_203__1_,r_n_203__0_,r_n_202__63_,r_n_202__62_,r_n_202__61_,r_n_202__60_,
  r_n_202__59_,r_n_202__58_,r_n_202__57_,r_n_202__56_,r_n_202__55_,r_n_202__54_,
  r_n_202__53_,r_n_202__52_,r_n_202__51_,r_n_202__50_,r_n_202__49_,r_n_202__48_,r_n_202__47_,
  r_n_202__46_,r_n_202__45_,r_n_202__44_,r_n_202__43_,r_n_202__42_,r_n_202__41_,
  r_n_202__40_,r_n_202__39_,r_n_202__38_,r_n_202__37_,r_n_202__36_,r_n_202__35_,
  r_n_202__34_,r_n_202__33_,r_n_202__32_,r_n_202__31_,r_n_202__30_,r_n_202__29_,
  r_n_202__28_,r_n_202__27_,r_n_202__26_,r_n_202__25_,r_n_202__24_,r_n_202__23_,
  r_n_202__22_,r_n_202__21_,r_n_202__20_,r_n_202__19_,r_n_202__18_,r_n_202__17_,
  r_n_202__16_,r_n_202__15_,r_n_202__14_,r_n_202__13_,r_n_202__12_,r_n_202__11_,r_n_202__10_,
  r_n_202__9_,r_n_202__8_,r_n_202__7_,r_n_202__6_,r_n_202__5_,r_n_202__4_,
  r_n_202__3_,r_n_202__2_,r_n_202__1_,r_n_202__0_,r_n_201__63_,r_n_201__62_,r_n_201__61_,
  r_n_201__60_,r_n_201__59_,r_n_201__58_,r_n_201__57_,r_n_201__56_,r_n_201__55_,
  r_n_201__54_,r_n_201__53_,r_n_201__52_,r_n_201__51_,r_n_201__50_,r_n_201__49_,
  r_n_201__48_,r_n_201__47_,r_n_201__46_,r_n_201__45_,r_n_201__44_,r_n_201__43_,
  r_n_201__42_,r_n_201__41_,r_n_201__40_,r_n_201__39_,r_n_201__38_,r_n_201__37_,
  r_n_201__36_,r_n_201__35_,r_n_201__34_,r_n_201__33_,r_n_201__32_,r_n_201__31_,
  r_n_201__30_,r_n_201__29_,r_n_201__28_,r_n_201__27_,r_n_201__26_,r_n_201__25_,r_n_201__24_,
  r_n_201__23_,r_n_201__22_,r_n_201__21_,r_n_201__20_,r_n_201__19_,r_n_201__18_,
  r_n_201__17_,r_n_201__16_,r_n_201__15_,r_n_201__14_,r_n_201__13_,r_n_201__12_,
  r_n_201__11_,r_n_201__10_,r_n_201__9_,r_n_201__8_,r_n_201__7_,r_n_201__6_,
  r_n_201__5_,r_n_201__4_,r_n_201__3_,r_n_201__2_,r_n_201__1_,r_n_201__0_,r_n_216__63_,
  r_n_216__62_,r_n_216__61_,r_n_216__60_,r_n_216__59_,r_n_216__58_,r_n_216__57_,
  r_n_216__56_,r_n_216__55_,r_n_216__54_,r_n_216__53_,r_n_216__52_,r_n_216__51_,
  r_n_216__50_,r_n_216__49_,r_n_216__48_,r_n_216__47_,r_n_216__46_,r_n_216__45_,
  r_n_216__44_,r_n_216__43_,r_n_216__42_,r_n_216__41_,r_n_216__40_,r_n_216__39_,r_n_216__38_,
  r_n_216__37_,r_n_216__36_,r_n_216__35_,r_n_216__34_,r_n_216__33_,r_n_216__32_,
  r_n_216__31_,r_n_216__30_,r_n_216__29_,r_n_216__28_,r_n_216__27_,r_n_216__26_,
  r_n_216__25_,r_n_216__24_,r_n_216__23_,r_n_216__22_,r_n_216__21_,r_n_216__20_,
  r_n_216__19_,r_n_216__18_,r_n_216__17_,r_n_216__16_,r_n_216__15_,r_n_216__14_,
  r_n_216__13_,r_n_216__12_,r_n_216__11_,r_n_216__10_,r_n_216__9_,r_n_216__8_,r_n_216__7_,
  r_n_216__6_,r_n_216__5_,r_n_216__4_,r_n_216__3_,r_n_216__2_,r_n_216__1_,
  r_n_216__0_,r_n_215__63_,r_n_215__62_,r_n_215__61_,r_n_215__60_,r_n_215__59_,
  r_n_215__58_,r_n_215__57_,r_n_215__56_,r_n_215__55_,r_n_215__54_,r_n_215__53_,r_n_215__52_,
  r_n_215__51_,r_n_215__50_,r_n_215__49_,r_n_215__48_,r_n_215__47_,r_n_215__46_,
  r_n_215__45_,r_n_215__44_,r_n_215__43_,r_n_215__42_,r_n_215__41_,r_n_215__40_,
  r_n_215__39_,r_n_215__38_,r_n_215__37_,r_n_215__36_,r_n_215__35_,r_n_215__34_,
  r_n_215__33_,r_n_215__32_,r_n_215__31_,r_n_215__30_,r_n_215__29_,r_n_215__28_,
  r_n_215__27_,r_n_215__26_,r_n_215__25_,r_n_215__24_,r_n_215__23_,r_n_215__22_,
  r_n_215__21_,r_n_215__20_,r_n_215__19_,r_n_215__18_,r_n_215__17_,r_n_215__16_,
  r_n_215__15_,r_n_215__14_,r_n_215__13_,r_n_215__12_,r_n_215__11_,r_n_215__10_,r_n_215__9_,
  r_n_215__8_,r_n_215__7_,r_n_215__6_,r_n_215__5_,r_n_215__4_,r_n_215__3_,
  r_n_215__2_,r_n_215__1_,r_n_215__0_,r_n_214__63_,r_n_214__62_,r_n_214__61_,r_n_214__60_,
  r_n_214__59_,r_n_214__58_,r_n_214__57_,r_n_214__56_,r_n_214__55_,r_n_214__54_,
  r_n_214__53_,r_n_214__52_,r_n_214__51_,r_n_214__50_,r_n_214__49_,r_n_214__48_,
  r_n_214__47_,r_n_214__46_,r_n_214__45_,r_n_214__44_,r_n_214__43_,r_n_214__42_,
  r_n_214__41_,r_n_214__40_,r_n_214__39_,r_n_214__38_,r_n_214__37_,r_n_214__36_,
  r_n_214__35_,r_n_214__34_,r_n_214__33_,r_n_214__32_,r_n_214__31_,r_n_214__30_,
  r_n_214__29_,r_n_214__28_,r_n_214__27_,r_n_214__26_,r_n_214__25_,r_n_214__24_,r_n_214__23_,
  r_n_214__22_,r_n_214__21_,r_n_214__20_,r_n_214__19_,r_n_214__18_,r_n_214__17_,
  r_n_214__16_,r_n_214__15_,r_n_214__14_,r_n_214__13_,r_n_214__12_,r_n_214__11_,
  r_n_214__10_,r_n_214__9_,r_n_214__8_,r_n_214__7_,r_n_214__6_,r_n_214__5_,r_n_214__4_,
  r_n_214__3_,r_n_214__2_,r_n_214__1_,r_n_214__0_,r_n_213__63_,r_n_213__62_,
  r_n_213__61_,r_n_213__60_,r_n_213__59_,r_n_213__58_,r_n_213__57_,r_n_213__56_,
  r_n_213__55_,r_n_213__54_,r_n_213__53_,r_n_213__52_,r_n_213__51_,r_n_213__50_,
  r_n_213__49_,r_n_213__48_,r_n_213__47_,r_n_213__46_,r_n_213__45_,r_n_213__44_,
  r_n_213__43_,r_n_213__42_,r_n_213__41_,r_n_213__40_,r_n_213__39_,r_n_213__38_,r_n_213__37_,
  r_n_213__36_,r_n_213__35_,r_n_213__34_,r_n_213__33_,r_n_213__32_,r_n_213__31_,
  r_n_213__30_,r_n_213__29_,r_n_213__28_,r_n_213__27_,r_n_213__26_,r_n_213__25_,
  r_n_213__24_,r_n_213__23_,r_n_213__22_,r_n_213__21_,r_n_213__20_,r_n_213__19_,
  r_n_213__18_,r_n_213__17_,r_n_213__16_,r_n_213__15_,r_n_213__14_,r_n_213__13_,
  r_n_213__12_,r_n_213__11_,r_n_213__10_,r_n_213__9_,r_n_213__8_,r_n_213__7_,r_n_213__6_,
  r_n_213__5_,r_n_213__4_,r_n_213__3_,r_n_213__2_,r_n_213__1_,r_n_213__0_,
  r_n_212__63_,r_n_212__62_,r_n_212__61_,r_n_212__60_,r_n_212__59_,r_n_212__58_,
  r_n_212__57_,r_n_212__56_,r_n_212__55_,r_n_212__54_,r_n_212__53_,r_n_212__52_,r_n_212__51_,
  r_n_212__50_,r_n_212__49_,r_n_212__48_,r_n_212__47_,r_n_212__46_,r_n_212__45_,
  r_n_212__44_,r_n_212__43_,r_n_212__42_,r_n_212__41_,r_n_212__40_,r_n_212__39_,
  r_n_212__38_,r_n_212__37_,r_n_212__36_,r_n_212__35_,r_n_212__34_,r_n_212__33_,
  r_n_212__32_,r_n_212__31_,r_n_212__30_,r_n_212__29_,r_n_212__28_,r_n_212__27_,
  r_n_212__26_,r_n_212__25_,r_n_212__24_,r_n_212__23_,r_n_212__22_,r_n_212__21_,
  r_n_212__20_,r_n_212__19_,r_n_212__18_,r_n_212__17_,r_n_212__16_,r_n_212__15_,r_n_212__14_,
  r_n_212__13_,r_n_212__12_,r_n_212__11_,r_n_212__10_,r_n_212__9_,r_n_212__8_,
  r_n_212__7_,r_n_212__6_,r_n_212__5_,r_n_212__4_,r_n_212__3_,r_n_212__2_,r_n_212__1_,
  r_n_212__0_,r_n_211__63_,r_n_211__62_,r_n_211__61_,r_n_211__60_,r_n_211__59_,
  r_n_211__58_,r_n_211__57_,r_n_211__56_,r_n_211__55_,r_n_211__54_,r_n_211__53_,
  r_n_211__52_,r_n_211__51_,r_n_211__50_,r_n_211__49_,r_n_211__48_,r_n_211__47_,
  r_n_211__46_,r_n_211__45_,r_n_211__44_,r_n_211__43_,r_n_211__42_,r_n_211__41_,
  r_n_211__40_,r_n_211__39_,r_n_211__38_,r_n_211__37_,r_n_211__36_,r_n_211__35_,
  r_n_211__34_,r_n_211__33_,r_n_211__32_,r_n_211__31_,r_n_211__30_,r_n_211__29_,r_n_211__28_,
  r_n_211__27_,r_n_211__26_,r_n_211__25_,r_n_211__24_,r_n_211__23_,r_n_211__22_,
  r_n_211__21_,r_n_211__20_,r_n_211__19_,r_n_211__18_,r_n_211__17_,r_n_211__16_,
  r_n_211__15_,r_n_211__14_,r_n_211__13_,r_n_211__12_,r_n_211__11_,r_n_211__10_,
  r_n_211__9_,r_n_211__8_,r_n_211__7_,r_n_211__6_,r_n_211__5_,r_n_211__4_,r_n_211__3_,
  r_n_211__2_,r_n_211__1_,r_n_211__0_,r_n_210__63_,r_n_210__62_,r_n_210__61_,
  r_n_210__60_,r_n_210__59_,r_n_210__58_,r_n_210__57_,r_n_210__56_,r_n_210__55_,
  r_n_210__54_,r_n_210__53_,r_n_210__52_,r_n_210__51_,r_n_210__50_,r_n_210__49_,
  r_n_210__48_,r_n_210__47_,r_n_210__46_,r_n_210__45_,r_n_210__44_,r_n_210__43_,r_n_210__42_,
  r_n_210__41_,r_n_210__40_,r_n_210__39_,r_n_210__38_,r_n_210__37_,r_n_210__36_,
  r_n_210__35_,r_n_210__34_,r_n_210__33_,r_n_210__32_,r_n_210__31_,r_n_210__30_,
  r_n_210__29_,r_n_210__28_,r_n_210__27_,r_n_210__26_,r_n_210__25_,r_n_210__24_,
  r_n_210__23_,r_n_210__22_,r_n_210__21_,r_n_210__20_,r_n_210__19_,r_n_210__18_,
  r_n_210__17_,r_n_210__16_,r_n_210__15_,r_n_210__14_,r_n_210__13_,r_n_210__12_,
  r_n_210__11_,r_n_210__10_,r_n_210__9_,r_n_210__8_,r_n_210__7_,r_n_210__6_,r_n_210__5_,
  r_n_210__4_,r_n_210__3_,r_n_210__2_,r_n_210__1_,r_n_210__0_,r_n_209__63_,
  r_n_209__62_,r_n_209__61_,r_n_209__60_,r_n_209__59_,r_n_209__58_,r_n_209__57_,r_n_209__56_,
  r_n_209__55_,r_n_209__54_,r_n_209__53_,r_n_209__52_,r_n_209__51_,r_n_209__50_,
  r_n_209__49_,r_n_209__48_,r_n_209__47_,r_n_209__46_,r_n_209__45_,r_n_209__44_,
  r_n_209__43_,r_n_209__42_,r_n_209__41_,r_n_209__40_,r_n_209__39_,r_n_209__38_,
  r_n_209__37_,r_n_209__36_,r_n_209__35_,r_n_209__34_,r_n_209__33_,r_n_209__32_,
  r_n_209__31_,r_n_209__30_,r_n_209__29_,r_n_209__28_,r_n_209__27_,r_n_209__26_,
  r_n_209__25_,r_n_209__24_,r_n_209__23_,r_n_209__22_,r_n_209__21_,r_n_209__20_,
  r_n_209__19_,r_n_209__18_,r_n_209__17_,r_n_209__16_,r_n_209__15_,r_n_209__14_,r_n_209__13_,
  r_n_209__12_,r_n_209__11_,r_n_209__10_,r_n_209__9_,r_n_209__8_,r_n_209__7_,
  r_n_209__6_,r_n_209__5_,r_n_209__4_,r_n_209__3_,r_n_209__2_,r_n_209__1_,r_n_209__0_,
  r_n_224__63_,r_n_224__62_,r_n_224__61_,r_n_224__60_,r_n_224__59_,r_n_224__58_,
  r_n_224__57_,r_n_224__56_,r_n_224__55_,r_n_224__54_,r_n_224__53_,r_n_224__52_,
  r_n_224__51_,r_n_224__50_,r_n_224__49_,r_n_224__48_,r_n_224__47_,r_n_224__46_,
  r_n_224__45_,r_n_224__44_,r_n_224__43_,r_n_224__42_,r_n_224__41_,r_n_224__40_,
  r_n_224__39_,r_n_224__38_,r_n_224__37_,r_n_224__36_,r_n_224__35_,r_n_224__34_,
  r_n_224__33_,r_n_224__32_,r_n_224__31_,r_n_224__30_,r_n_224__29_,r_n_224__28_,r_n_224__27_,
  r_n_224__26_,r_n_224__25_,r_n_224__24_,r_n_224__23_,r_n_224__22_,r_n_224__21_,
  r_n_224__20_,r_n_224__19_,r_n_224__18_,r_n_224__17_,r_n_224__16_,r_n_224__15_,
  r_n_224__14_,r_n_224__13_,r_n_224__12_,r_n_224__11_,r_n_224__10_,r_n_224__9_,
  r_n_224__8_,r_n_224__7_,r_n_224__6_,r_n_224__5_,r_n_224__4_,r_n_224__3_,r_n_224__2_,
  r_n_224__1_,r_n_224__0_,r_n_223__63_,r_n_223__62_,r_n_223__61_,r_n_223__60_,
  r_n_223__59_,r_n_223__58_,r_n_223__57_,r_n_223__56_,r_n_223__55_,r_n_223__54_,
  r_n_223__53_,r_n_223__52_,r_n_223__51_,r_n_223__50_,r_n_223__49_,r_n_223__48_,
  r_n_223__47_,r_n_223__46_,r_n_223__45_,r_n_223__44_,r_n_223__43_,r_n_223__42_,r_n_223__41_,
  r_n_223__40_,r_n_223__39_,r_n_223__38_,r_n_223__37_,r_n_223__36_,r_n_223__35_,
  r_n_223__34_,r_n_223__33_,r_n_223__32_,r_n_223__31_,r_n_223__30_,r_n_223__29_,
  r_n_223__28_,r_n_223__27_,r_n_223__26_,r_n_223__25_,r_n_223__24_,r_n_223__23_,
  r_n_223__22_,r_n_223__21_,r_n_223__20_,r_n_223__19_,r_n_223__18_,r_n_223__17_,
  r_n_223__16_,r_n_223__15_,r_n_223__14_,r_n_223__13_,r_n_223__12_,r_n_223__11_,
  r_n_223__10_,r_n_223__9_,r_n_223__8_,r_n_223__7_,r_n_223__6_,r_n_223__5_,r_n_223__4_,
  r_n_223__3_,r_n_223__2_,r_n_223__1_,r_n_223__0_,r_n_222__63_,r_n_222__62_,
  r_n_222__61_,r_n_222__60_,r_n_222__59_,r_n_222__58_,r_n_222__57_,r_n_222__56_,r_n_222__55_,
  r_n_222__54_,r_n_222__53_,r_n_222__52_,r_n_222__51_,r_n_222__50_,r_n_222__49_,
  r_n_222__48_,r_n_222__47_,r_n_222__46_,r_n_222__45_,r_n_222__44_,r_n_222__43_,
  r_n_222__42_,r_n_222__41_,r_n_222__40_,r_n_222__39_,r_n_222__38_,r_n_222__37_,
  r_n_222__36_,r_n_222__35_,r_n_222__34_,r_n_222__33_,r_n_222__32_,r_n_222__31_,
  r_n_222__30_,r_n_222__29_,r_n_222__28_,r_n_222__27_,r_n_222__26_,r_n_222__25_,
  r_n_222__24_,r_n_222__23_,r_n_222__22_,r_n_222__21_,r_n_222__20_,r_n_222__19_,r_n_222__18_,
  r_n_222__17_,r_n_222__16_,r_n_222__15_,r_n_222__14_,r_n_222__13_,r_n_222__12_,
  r_n_222__11_,r_n_222__10_,r_n_222__9_,r_n_222__8_,r_n_222__7_,r_n_222__6_,
  r_n_222__5_,r_n_222__4_,r_n_222__3_,r_n_222__2_,r_n_222__1_,r_n_222__0_,r_n_221__63_,
  r_n_221__62_,r_n_221__61_,r_n_221__60_,r_n_221__59_,r_n_221__58_,r_n_221__57_,
  r_n_221__56_,r_n_221__55_,r_n_221__54_,r_n_221__53_,r_n_221__52_,r_n_221__51_,
  r_n_221__50_,r_n_221__49_,r_n_221__48_,r_n_221__47_,r_n_221__46_,r_n_221__45_,
  r_n_221__44_,r_n_221__43_,r_n_221__42_,r_n_221__41_,r_n_221__40_,r_n_221__39_,
  r_n_221__38_,r_n_221__37_,r_n_221__36_,r_n_221__35_,r_n_221__34_,r_n_221__33_,r_n_221__32_,
  r_n_221__31_,r_n_221__30_,r_n_221__29_,r_n_221__28_,r_n_221__27_,r_n_221__26_,
  r_n_221__25_,r_n_221__24_,r_n_221__23_,r_n_221__22_,r_n_221__21_,r_n_221__20_,
  r_n_221__19_,r_n_221__18_,r_n_221__17_,r_n_221__16_,r_n_221__15_,r_n_221__14_,
  r_n_221__13_,r_n_221__12_,r_n_221__11_,r_n_221__10_,r_n_221__9_,r_n_221__8_,
  r_n_221__7_,r_n_221__6_,r_n_221__5_,r_n_221__4_,r_n_221__3_,r_n_221__2_,r_n_221__1_,
  r_n_221__0_,r_n_220__63_,r_n_220__62_,r_n_220__61_,r_n_220__60_,r_n_220__59_,
  r_n_220__58_,r_n_220__57_,r_n_220__56_,r_n_220__55_,r_n_220__54_,r_n_220__53_,
  r_n_220__52_,r_n_220__51_,r_n_220__50_,r_n_220__49_,r_n_220__48_,r_n_220__47_,r_n_220__46_,
  r_n_220__45_,r_n_220__44_,r_n_220__43_,r_n_220__42_,r_n_220__41_,r_n_220__40_,
  r_n_220__39_,r_n_220__38_,r_n_220__37_,r_n_220__36_,r_n_220__35_,r_n_220__34_,
  r_n_220__33_,r_n_220__32_,r_n_220__31_,r_n_220__30_,r_n_220__29_,r_n_220__28_,
  r_n_220__27_,r_n_220__26_,r_n_220__25_,r_n_220__24_,r_n_220__23_,r_n_220__22_,
  r_n_220__21_,r_n_220__20_,r_n_220__19_,r_n_220__18_,r_n_220__17_,r_n_220__16_,
  r_n_220__15_,r_n_220__14_,r_n_220__13_,r_n_220__12_,r_n_220__11_,r_n_220__10_,r_n_220__9_,
  r_n_220__8_,r_n_220__7_,r_n_220__6_,r_n_220__5_,r_n_220__4_,r_n_220__3_,
  r_n_220__2_,r_n_220__1_,r_n_220__0_,r_n_219__63_,r_n_219__62_,r_n_219__61_,r_n_219__60_,
  r_n_219__59_,r_n_219__58_,r_n_219__57_,r_n_219__56_,r_n_219__55_,r_n_219__54_,
  r_n_219__53_,r_n_219__52_,r_n_219__51_,r_n_219__50_,r_n_219__49_,r_n_219__48_,
  r_n_219__47_,r_n_219__46_,r_n_219__45_,r_n_219__44_,r_n_219__43_,r_n_219__42_,
  r_n_219__41_,r_n_219__40_,r_n_219__39_,r_n_219__38_,r_n_219__37_,r_n_219__36_,
  r_n_219__35_,r_n_219__34_,r_n_219__33_,r_n_219__32_,r_n_219__31_,r_n_219__30_,
  r_n_219__29_,r_n_219__28_,r_n_219__27_,r_n_219__26_,r_n_219__25_,r_n_219__24_,
  r_n_219__23_,r_n_219__22_,r_n_219__21_,r_n_219__20_,r_n_219__19_,r_n_219__18_,r_n_219__17_,
  r_n_219__16_,r_n_219__15_,r_n_219__14_,r_n_219__13_,r_n_219__12_,r_n_219__11_,
  r_n_219__10_,r_n_219__9_,r_n_219__8_,r_n_219__7_,r_n_219__6_,r_n_219__5_,
  r_n_219__4_,r_n_219__3_,r_n_219__2_,r_n_219__1_,r_n_219__0_,r_n_218__63_,r_n_218__62_,
  r_n_218__61_,r_n_218__60_,r_n_218__59_,r_n_218__58_,r_n_218__57_,r_n_218__56_,
  r_n_218__55_,r_n_218__54_,r_n_218__53_,r_n_218__52_,r_n_218__51_,r_n_218__50_,
  r_n_218__49_,r_n_218__48_,r_n_218__47_,r_n_218__46_,r_n_218__45_,r_n_218__44_,
  r_n_218__43_,r_n_218__42_,r_n_218__41_,r_n_218__40_,r_n_218__39_,r_n_218__38_,
  r_n_218__37_,r_n_218__36_,r_n_218__35_,r_n_218__34_,r_n_218__33_,r_n_218__32_,r_n_218__31_,
  r_n_218__30_,r_n_218__29_,r_n_218__28_,r_n_218__27_,r_n_218__26_,r_n_218__25_,
  r_n_218__24_,r_n_218__23_,r_n_218__22_,r_n_218__21_,r_n_218__20_,r_n_218__19_,
  r_n_218__18_,r_n_218__17_,r_n_218__16_,r_n_218__15_,r_n_218__14_,r_n_218__13_,
  r_n_218__12_,r_n_218__11_,r_n_218__10_,r_n_218__9_,r_n_218__8_,r_n_218__7_,r_n_218__6_,
  r_n_218__5_,r_n_218__4_,r_n_218__3_,r_n_218__2_,r_n_218__1_,r_n_218__0_,
  r_n_217__63_,r_n_217__62_,r_n_217__61_,r_n_217__60_,r_n_217__59_,r_n_217__58_,
  r_n_217__57_,r_n_217__56_,r_n_217__55_,r_n_217__54_,r_n_217__53_,r_n_217__52_,
  r_n_217__51_,r_n_217__50_,r_n_217__49_,r_n_217__48_,r_n_217__47_,r_n_217__46_,r_n_217__45_,
  r_n_217__44_,r_n_217__43_,r_n_217__42_,r_n_217__41_,r_n_217__40_,r_n_217__39_,
  r_n_217__38_,r_n_217__37_,r_n_217__36_,r_n_217__35_,r_n_217__34_,r_n_217__33_,
  r_n_217__32_,r_n_217__31_,r_n_217__30_,r_n_217__29_,r_n_217__28_,r_n_217__27_,
  r_n_217__26_,r_n_217__25_,r_n_217__24_,r_n_217__23_,r_n_217__22_,r_n_217__21_,
  r_n_217__20_,r_n_217__19_,r_n_217__18_,r_n_217__17_,r_n_217__16_,r_n_217__15_,
  r_n_217__14_,r_n_217__13_,r_n_217__12_,r_n_217__11_,r_n_217__10_,r_n_217__9_,r_n_217__8_,
  r_n_217__7_,r_n_217__6_,r_n_217__5_,r_n_217__4_,r_n_217__3_,r_n_217__2_,
  r_n_217__1_,r_n_217__0_,r_n_232__63_,r_n_232__62_,r_n_232__61_,r_n_232__60_,r_n_232__59_,
  r_n_232__58_,r_n_232__57_,r_n_232__56_,r_n_232__55_,r_n_232__54_,r_n_232__53_,
  r_n_232__52_,r_n_232__51_,r_n_232__50_,r_n_232__49_,r_n_232__48_,r_n_232__47_,
  r_n_232__46_,r_n_232__45_,r_n_232__44_,r_n_232__43_,r_n_232__42_,r_n_232__41_,
  r_n_232__40_,r_n_232__39_,r_n_232__38_,r_n_232__37_,r_n_232__36_,r_n_232__35_,
  r_n_232__34_,r_n_232__33_,r_n_232__32_,r_n_232__31_,r_n_232__30_,r_n_232__29_,
  r_n_232__28_,r_n_232__27_,r_n_232__26_,r_n_232__25_,r_n_232__24_,r_n_232__23_,r_n_232__22_,
  r_n_232__21_,r_n_232__20_,r_n_232__19_,r_n_232__18_,r_n_232__17_,r_n_232__16_,
  r_n_232__15_,r_n_232__14_,r_n_232__13_,r_n_232__12_,r_n_232__11_,r_n_232__10_,
  r_n_232__9_,r_n_232__8_,r_n_232__7_,r_n_232__6_,r_n_232__5_,r_n_232__4_,r_n_232__3_,
  r_n_232__2_,r_n_232__1_,r_n_232__0_,r_n_231__63_,r_n_231__62_,r_n_231__61_,
  r_n_231__60_,r_n_231__59_,r_n_231__58_,r_n_231__57_,r_n_231__56_,r_n_231__55_,
  r_n_231__54_,r_n_231__53_,r_n_231__52_,r_n_231__51_,r_n_231__50_,r_n_231__49_,
  r_n_231__48_,r_n_231__47_,r_n_231__46_,r_n_231__45_,r_n_231__44_,r_n_231__43_,
  r_n_231__42_,r_n_231__41_,r_n_231__40_,r_n_231__39_,r_n_231__38_,r_n_231__37_,r_n_231__36_,
  r_n_231__35_,r_n_231__34_,r_n_231__33_,r_n_231__32_,r_n_231__31_,r_n_231__30_,
  r_n_231__29_,r_n_231__28_,r_n_231__27_,r_n_231__26_,r_n_231__25_,r_n_231__24_,
  r_n_231__23_,r_n_231__22_,r_n_231__21_,r_n_231__20_,r_n_231__19_,r_n_231__18_,
  r_n_231__17_,r_n_231__16_,r_n_231__15_,r_n_231__14_,r_n_231__13_,r_n_231__12_,
  r_n_231__11_,r_n_231__10_,r_n_231__9_,r_n_231__8_,r_n_231__7_,r_n_231__6_,r_n_231__5_,
  r_n_231__4_,r_n_231__3_,r_n_231__2_,r_n_231__1_,r_n_231__0_,r_n_230__63_,
  r_n_230__62_,r_n_230__61_,r_n_230__60_,r_n_230__59_,r_n_230__58_,r_n_230__57_,
  r_n_230__56_,r_n_230__55_,r_n_230__54_,r_n_230__53_,r_n_230__52_,r_n_230__51_,r_n_230__50_,
  r_n_230__49_,r_n_230__48_,r_n_230__47_,r_n_230__46_,r_n_230__45_,r_n_230__44_,
  r_n_230__43_,r_n_230__42_,r_n_230__41_,r_n_230__40_,r_n_230__39_,r_n_230__38_,
  r_n_230__37_,r_n_230__36_,r_n_230__35_,r_n_230__34_,r_n_230__33_,r_n_230__32_,
  r_n_230__31_,r_n_230__30_,r_n_230__29_,r_n_230__28_,r_n_230__27_,r_n_230__26_,
  r_n_230__25_,r_n_230__24_,r_n_230__23_,r_n_230__22_,r_n_230__21_,r_n_230__20_,
  r_n_230__19_,r_n_230__18_,r_n_230__17_,r_n_230__16_,r_n_230__15_,r_n_230__14_,
  r_n_230__13_,r_n_230__12_,r_n_230__11_,r_n_230__10_,r_n_230__9_,r_n_230__8_,r_n_230__7_,
  r_n_230__6_,r_n_230__5_,r_n_230__4_,r_n_230__3_,r_n_230__2_,r_n_230__1_,r_n_230__0_,
  r_n_229__63_,r_n_229__62_,r_n_229__61_,r_n_229__60_,r_n_229__59_,r_n_229__58_,
  r_n_229__57_,r_n_229__56_,r_n_229__55_,r_n_229__54_,r_n_229__53_,r_n_229__52_,
  r_n_229__51_,r_n_229__50_,r_n_229__49_,r_n_229__48_,r_n_229__47_,r_n_229__46_,
  r_n_229__45_,r_n_229__44_,r_n_229__43_,r_n_229__42_,r_n_229__41_,r_n_229__40_,
  r_n_229__39_,r_n_229__38_,r_n_229__37_,r_n_229__36_,r_n_229__35_,r_n_229__34_,
  r_n_229__33_,r_n_229__32_,r_n_229__31_,r_n_229__30_,r_n_229__29_,r_n_229__28_,
  r_n_229__27_,r_n_229__26_,r_n_229__25_,r_n_229__24_,r_n_229__23_,r_n_229__22_,r_n_229__21_,
  r_n_229__20_,r_n_229__19_,r_n_229__18_,r_n_229__17_,r_n_229__16_,r_n_229__15_,
  r_n_229__14_,r_n_229__13_,r_n_229__12_,r_n_229__11_,r_n_229__10_,r_n_229__9_,
  r_n_229__8_,r_n_229__7_,r_n_229__6_,r_n_229__5_,r_n_229__4_,r_n_229__3_,r_n_229__2_,
  r_n_229__1_,r_n_229__0_,r_n_228__63_,r_n_228__62_,r_n_228__61_,r_n_228__60_,
  r_n_228__59_,r_n_228__58_,r_n_228__57_,r_n_228__56_,r_n_228__55_,r_n_228__54_,
  r_n_228__53_,r_n_228__52_,r_n_228__51_,r_n_228__50_,r_n_228__49_,r_n_228__48_,
  r_n_228__47_,r_n_228__46_,r_n_228__45_,r_n_228__44_,r_n_228__43_,r_n_228__42_,
  r_n_228__41_,r_n_228__40_,r_n_228__39_,r_n_228__38_,r_n_228__37_,r_n_228__36_,r_n_228__35_,
  r_n_228__34_,r_n_228__33_,r_n_228__32_,r_n_228__31_,r_n_228__30_,r_n_228__29_,
  r_n_228__28_,r_n_228__27_,r_n_228__26_,r_n_228__25_,r_n_228__24_,r_n_228__23_,
  r_n_228__22_,r_n_228__21_,r_n_228__20_,r_n_228__19_,r_n_228__18_,r_n_228__17_,
  r_n_228__16_,r_n_228__15_,r_n_228__14_,r_n_228__13_,r_n_228__12_,r_n_228__11_,
  r_n_228__10_,r_n_228__9_,r_n_228__8_,r_n_228__7_,r_n_228__6_,r_n_228__5_,r_n_228__4_,
  r_n_228__3_,r_n_228__2_,r_n_228__1_,r_n_228__0_,r_n_227__63_,r_n_227__62_,
  r_n_227__61_,r_n_227__60_,r_n_227__59_,r_n_227__58_,r_n_227__57_,r_n_227__56_,
  r_n_227__55_,r_n_227__54_,r_n_227__53_,r_n_227__52_,r_n_227__51_,r_n_227__50_,r_n_227__49_,
  r_n_227__48_,r_n_227__47_,r_n_227__46_,r_n_227__45_,r_n_227__44_,r_n_227__43_,
  r_n_227__42_,r_n_227__41_,r_n_227__40_,r_n_227__39_,r_n_227__38_,r_n_227__37_,
  r_n_227__36_,r_n_227__35_,r_n_227__34_,r_n_227__33_,r_n_227__32_,r_n_227__31_,
  r_n_227__30_,r_n_227__29_,r_n_227__28_,r_n_227__27_,r_n_227__26_,r_n_227__25_,
  r_n_227__24_,r_n_227__23_,r_n_227__22_,r_n_227__21_,r_n_227__20_,r_n_227__19_,
  r_n_227__18_,r_n_227__17_,r_n_227__16_,r_n_227__15_,r_n_227__14_,r_n_227__13_,r_n_227__12_,
  r_n_227__11_,r_n_227__10_,r_n_227__9_,r_n_227__8_,r_n_227__7_,r_n_227__6_,
  r_n_227__5_,r_n_227__4_,r_n_227__3_,r_n_227__2_,r_n_227__1_,r_n_227__0_,r_n_226__63_,
  r_n_226__62_,r_n_226__61_,r_n_226__60_,r_n_226__59_,r_n_226__58_,r_n_226__57_,
  r_n_226__56_,r_n_226__55_,r_n_226__54_,r_n_226__53_,r_n_226__52_,r_n_226__51_,
  r_n_226__50_,r_n_226__49_,r_n_226__48_,r_n_226__47_,r_n_226__46_,r_n_226__45_,
  r_n_226__44_,r_n_226__43_,r_n_226__42_,r_n_226__41_,r_n_226__40_,r_n_226__39_,
  r_n_226__38_,r_n_226__37_,r_n_226__36_,r_n_226__35_,r_n_226__34_,r_n_226__33_,
  r_n_226__32_,r_n_226__31_,r_n_226__30_,r_n_226__29_,r_n_226__28_,r_n_226__27_,r_n_226__26_,
  r_n_226__25_,r_n_226__24_,r_n_226__23_,r_n_226__22_,r_n_226__21_,r_n_226__20_,
  r_n_226__19_,r_n_226__18_,r_n_226__17_,r_n_226__16_,r_n_226__15_,r_n_226__14_,
  r_n_226__13_,r_n_226__12_,r_n_226__11_,r_n_226__10_,r_n_226__9_,r_n_226__8_,
  r_n_226__7_,r_n_226__6_,r_n_226__5_,r_n_226__4_,r_n_226__3_,r_n_226__2_,r_n_226__1_,
  r_n_226__0_,r_n_225__63_,r_n_225__62_,r_n_225__61_,r_n_225__60_,r_n_225__59_,
  r_n_225__58_,r_n_225__57_,r_n_225__56_,r_n_225__55_,r_n_225__54_,r_n_225__53_,
  r_n_225__52_,r_n_225__51_,r_n_225__50_,r_n_225__49_,r_n_225__48_,r_n_225__47_,
  r_n_225__46_,r_n_225__45_,r_n_225__44_,r_n_225__43_,r_n_225__42_,r_n_225__41_,r_n_225__40_,
  r_n_225__39_,r_n_225__38_,r_n_225__37_,r_n_225__36_,r_n_225__35_,r_n_225__34_,
  r_n_225__33_,r_n_225__32_,r_n_225__31_,r_n_225__30_,r_n_225__29_,r_n_225__28_,
  r_n_225__27_,r_n_225__26_,r_n_225__25_,r_n_225__24_,r_n_225__23_,r_n_225__22_,
  r_n_225__21_,r_n_225__20_,r_n_225__19_,r_n_225__18_,r_n_225__17_,r_n_225__16_,
  r_n_225__15_,r_n_225__14_,r_n_225__13_,r_n_225__12_,r_n_225__11_,r_n_225__10_,
  r_n_225__9_,r_n_225__8_,r_n_225__7_,r_n_225__6_,r_n_225__5_,r_n_225__4_,r_n_225__3_,
  r_n_225__2_,r_n_225__1_,r_n_225__0_,r_n_240__63_,r_n_240__62_,r_n_240__61_,
  r_n_240__60_,r_n_240__59_,r_n_240__58_,r_n_240__57_,r_n_240__56_,r_n_240__55_,r_n_240__54_,
  r_n_240__53_,r_n_240__52_,r_n_240__51_,r_n_240__50_,r_n_240__49_,r_n_240__48_,
  r_n_240__47_,r_n_240__46_,r_n_240__45_,r_n_240__44_,r_n_240__43_,r_n_240__42_,
  r_n_240__41_,r_n_240__40_,r_n_240__39_,r_n_240__38_,r_n_240__37_,r_n_240__36_,
  r_n_240__35_,r_n_240__34_,r_n_240__33_,r_n_240__32_,r_n_240__31_,r_n_240__30_,
  r_n_240__29_,r_n_240__28_,r_n_240__27_,r_n_240__26_,r_n_240__25_,r_n_240__24_,
  r_n_240__23_,r_n_240__22_,r_n_240__21_,r_n_240__20_,r_n_240__19_,r_n_240__18_,
  r_n_240__17_,r_n_240__16_,r_n_240__15_,r_n_240__14_,r_n_240__13_,r_n_240__12_,r_n_240__11_,
  r_n_240__10_,r_n_240__9_,r_n_240__8_,r_n_240__7_,r_n_240__6_,r_n_240__5_,
  r_n_240__4_,r_n_240__3_,r_n_240__2_,r_n_240__1_,r_n_240__0_,r_n_239__63_,r_n_239__62_,
  r_n_239__61_,r_n_239__60_,r_n_239__59_,r_n_239__58_,r_n_239__57_,r_n_239__56_,
  r_n_239__55_,r_n_239__54_,r_n_239__53_,r_n_239__52_,r_n_239__51_,r_n_239__50_,
  r_n_239__49_,r_n_239__48_,r_n_239__47_,r_n_239__46_,r_n_239__45_,r_n_239__44_,
  r_n_239__43_,r_n_239__42_,r_n_239__41_,r_n_239__40_,r_n_239__39_,r_n_239__38_,
  r_n_239__37_,r_n_239__36_,r_n_239__35_,r_n_239__34_,r_n_239__33_,r_n_239__32_,
  r_n_239__31_,r_n_239__30_,r_n_239__29_,r_n_239__28_,r_n_239__27_,r_n_239__26_,r_n_239__25_,
  r_n_239__24_,r_n_239__23_,r_n_239__22_,r_n_239__21_,r_n_239__20_,r_n_239__19_,
  r_n_239__18_,r_n_239__17_,r_n_239__16_,r_n_239__15_,r_n_239__14_,r_n_239__13_,
  r_n_239__12_,r_n_239__11_,r_n_239__10_,r_n_239__9_,r_n_239__8_,r_n_239__7_,
  r_n_239__6_,r_n_239__5_,r_n_239__4_,r_n_239__3_,r_n_239__2_,r_n_239__1_,r_n_239__0_,
  r_n_238__63_,r_n_238__62_,r_n_238__61_,r_n_238__60_,r_n_238__59_,r_n_238__58_,
  r_n_238__57_,r_n_238__56_,r_n_238__55_,r_n_238__54_,r_n_238__53_,r_n_238__52_,
  r_n_238__51_,r_n_238__50_,r_n_238__49_,r_n_238__48_,r_n_238__47_,r_n_238__46_,
  r_n_238__45_,r_n_238__44_,r_n_238__43_,r_n_238__42_,r_n_238__41_,r_n_238__40_,r_n_238__39_,
  r_n_238__38_,r_n_238__37_,r_n_238__36_,r_n_238__35_,r_n_238__34_,r_n_238__33_,
  r_n_238__32_,r_n_238__31_,r_n_238__30_,r_n_238__29_,r_n_238__28_,r_n_238__27_,
  r_n_238__26_,r_n_238__25_,r_n_238__24_,r_n_238__23_,r_n_238__22_,r_n_238__21_,
  r_n_238__20_,r_n_238__19_,r_n_238__18_,r_n_238__17_,r_n_238__16_,r_n_238__15_,
  r_n_238__14_,r_n_238__13_,r_n_238__12_,r_n_238__11_,r_n_238__10_,r_n_238__9_,r_n_238__8_,
  r_n_238__7_,r_n_238__6_,r_n_238__5_,r_n_238__4_,r_n_238__3_,r_n_238__2_,
  r_n_238__1_,r_n_238__0_,r_n_237__63_,r_n_237__62_,r_n_237__61_,r_n_237__60_,
  r_n_237__59_,r_n_237__58_,r_n_237__57_,r_n_237__56_,r_n_237__55_,r_n_237__54_,r_n_237__53_,
  r_n_237__52_,r_n_237__51_,r_n_237__50_,r_n_237__49_,r_n_237__48_,r_n_237__47_,
  r_n_237__46_,r_n_237__45_,r_n_237__44_,r_n_237__43_,r_n_237__42_,r_n_237__41_,
  r_n_237__40_,r_n_237__39_,r_n_237__38_,r_n_237__37_,r_n_237__36_,r_n_237__35_,
  r_n_237__34_,r_n_237__33_,r_n_237__32_,r_n_237__31_,r_n_237__30_,r_n_237__29_,
  r_n_237__28_,r_n_237__27_,r_n_237__26_,r_n_237__25_,r_n_237__24_,r_n_237__23_,
  r_n_237__22_,r_n_237__21_,r_n_237__20_,r_n_237__19_,r_n_237__18_,r_n_237__17_,r_n_237__16_,
  r_n_237__15_,r_n_237__14_,r_n_237__13_,r_n_237__12_,r_n_237__11_,r_n_237__10_,
  r_n_237__9_,r_n_237__8_,r_n_237__7_,r_n_237__6_,r_n_237__5_,r_n_237__4_,
  r_n_237__3_,r_n_237__2_,r_n_237__1_,r_n_237__0_,r_n_236__63_,r_n_236__62_,r_n_236__61_,
  r_n_236__60_,r_n_236__59_,r_n_236__58_,r_n_236__57_,r_n_236__56_,r_n_236__55_,
  r_n_236__54_,r_n_236__53_,r_n_236__52_,r_n_236__51_,r_n_236__50_,r_n_236__49_,
  r_n_236__48_,r_n_236__47_,r_n_236__46_,r_n_236__45_,r_n_236__44_,r_n_236__43_,
  r_n_236__42_,r_n_236__41_,r_n_236__40_,r_n_236__39_,r_n_236__38_,r_n_236__37_,
  r_n_236__36_,r_n_236__35_,r_n_236__34_,r_n_236__33_,r_n_236__32_,r_n_236__31_,r_n_236__30_,
  r_n_236__29_,r_n_236__28_,r_n_236__27_,r_n_236__26_,r_n_236__25_,r_n_236__24_,
  r_n_236__23_,r_n_236__22_,r_n_236__21_,r_n_236__20_,r_n_236__19_,r_n_236__18_,
  r_n_236__17_,r_n_236__16_,r_n_236__15_,r_n_236__14_,r_n_236__13_,r_n_236__12_,
  r_n_236__11_,r_n_236__10_,r_n_236__9_,r_n_236__8_,r_n_236__7_,r_n_236__6_,r_n_236__5_,
  r_n_236__4_,r_n_236__3_,r_n_236__2_,r_n_236__1_,r_n_236__0_,r_n_235__63_,
  r_n_235__62_,r_n_235__61_,r_n_235__60_,r_n_235__59_,r_n_235__58_,r_n_235__57_,
  r_n_235__56_,r_n_235__55_,r_n_235__54_,r_n_235__53_,r_n_235__52_,r_n_235__51_,
  r_n_235__50_,r_n_235__49_,r_n_235__48_,r_n_235__47_,r_n_235__46_,r_n_235__45_,r_n_235__44_,
  r_n_235__43_,r_n_235__42_,r_n_235__41_,r_n_235__40_,r_n_235__39_,r_n_235__38_,
  r_n_235__37_,r_n_235__36_,r_n_235__35_,r_n_235__34_,r_n_235__33_,r_n_235__32_,
  r_n_235__31_,r_n_235__30_,r_n_235__29_,r_n_235__28_,r_n_235__27_,r_n_235__26_,
  r_n_235__25_,r_n_235__24_,r_n_235__23_,r_n_235__22_,r_n_235__21_,r_n_235__20_,
  r_n_235__19_,r_n_235__18_,r_n_235__17_,r_n_235__16_,r_n_235__15_,r_n_235__14_,
  r_n_235__13_,r_n_235__12_,r_n_235__11_,r_n_235__10_,r_n_235__9_,r_n_235__8_,r_n_235__7_,
  r_n_235__6_,r_n_235__5_,r_n_235__4_,r_n_235__3_,r_n_235__2_,r_n_235__1_,
  r_n_235__0_,r_n_234__63_,r_n_234__62_,r_n_234__61_,r_n_234__60_,r_n_234__59_,r_n_234__58_,
  r_n_234__57_,r_n_234__56_,r_n_234__55_,r_n_234__54_,r_n_234__53_,r_n_234__52_,
  r_n_234__51_,r_n_234__50_,r_n_234__49_,r_n_234__48_,r_n_234__47_,r_n_234__46_,
  r_n_234__45_,r_n_234__44_,r_n_234__43_,r_n_234__42_,r_n_234__41_,r_n_234__40_,
  r_n_234__39_,r_n_234__38_,r_n_234__37_,r_n_234__36_,r_n_234__35_,r_n_234__34_,
  r_n_234__33_,r_n_234__32_,r_n_234__31_,r_n_234__30_,r_n_234__29_,r_n_234__28_,
  r_n_234__27_,r_n_234__26_,r_n_234__25_,r_n_234__24_,r_n_234__23_,r_n_234__22_,
  r_n_234__21_,r_n_234__20_,r_n_234__19_,r_n_234__18_,r_n_234__17_,r_n_234__16_,r_n_234__15_,
  r_n_234__14_,r_n_234__13_,r_n_234__12_,r_n_234__11_,r_n_234__10_,r_n_234__9_,
  r_n_234__8_,r_n_234__7_,r_n_234__6_,r_n_234__5_,r_n_234__4_,r_n_234__3_,r_n_234__2_,
  r_n_234__1_,r_n_234__0_,r_n_233__63_,r_n_233__62_,r_n_233__61_,r_n_233__60_,
  r_n_233__59_,r_n_233__58_,r_n_233__57_,r_n_233__56_,r_n_233__55_,r_n_233__54_,
  r_n_233__53_,r_n_233__52_,r_n_233__51_,r_n_233__50_,r_n_233__49_,r_n_233__48_,
  r_n_233__47_,r_n_233__46_,r_n_233__45_,r_n_233__44_,r_n_233__43_,r_n_233__42_,
  r_n_233__41_,r_n_233__40_,r_n_233__39_,r_n_233__38_,r_n_233__37_,r_n_233__36_,
  r_n_233__35_,r_n_233__34_,r_n_233__33_,r_n_233__32_,r_n_233__31_,r_n_233__30_,r_n_233__29_,
  r_n_233__28_,r_n_233__27_,r_n_233__26_,r_n_233__25_,r_n_233__24_,r_n_233__23_,
  r_n_233__22_,r_n_233__21_,r_n_233__20_,r_n_233__19_,r_n_233__18_,r_n_233__17_,
  r_n_233__16_,r_n_233__15_,r_n_233__14_,r_n_233__13_,r_n_233__12_,r_n_233__11_,
  r_n_233__10_,r_n_233__9_,r_n_233__8_,r_n_233__7_,r_n_233__6_,r_n_233__5_,r_n_233__4_,
  r_n_233__3_,r_n_233__2_,r_n_233__1_,r_n_233__0_,r_n_248__63_,r_n_248__62_,
  r_n_248__61_,r_n_248__60_,r_n_248__59_,r_n_248__58_,r_n_248__57_,r_n_248__56_,
  r_n_248__55_,r_n_248__54_,r_n_248__53_,r_n_248__52_,r_n_248__51_,r_n_248__50_,
  r_n_248__49_,r_n_248__48_,r_n_248__47_,r_n_248__46_,r_n_248__45_,r_n_248__44_,r_n_248__43_,
  r_n_248__42_,r_n_248__41_,r_n_248__40_,r_n_248__39_,r_n_248__38_,r_n_248__37_,
  r_n_248__36_,r_n_248__35_,r_n_248__34_,r_n_248__33_,r_n_248__32_,r_n_248__31_,
  r_n_248__30_,r_n_248__29_,r_n_248__28_,r_n_248__27_,r_n_248__26_,r_n_248__25_,
  r_n_248__24_,r_n_248__23_,r_n_248__22_,r_n_248__21_,r_n_248__20_,r_n_248__19_,
  r_n_248__18_,r_n_248__17_,r_n_248__16_,r_n_248__15_,r_n_248__14_,r_n_248__13_,
  r_n_248__12_,r_n_248__11_,r_n_248__10_,r_n_248__9_,r_n_248__8_,r_n_248__7_,r_n_248__6_,
  r_n_248__5_,r_n_248__4_,r_n_248__3_,r_n_248__2_,r_n_248__1_,r_n_248__0_,
  r_n_247__63_,r_n_247__62_,r_n_247__61_,r_n_247__60_,r_n_247__59_,r_n_247__58_,r_n_247__57_,
  r_n_247__56_,r_n_247__55_,r_n_247__54_,r_n_247__53_,r_n_247__52_,r_n_247__51_,
  r_n_247__50_,r_n_247__49_,r_n_247__48_,r_n_247__47_,r_n_247__46_,r_n_247__45_,
  r_n_247__44_,r_n_247__43_,r_n_247__42_,r_n_247__41_,r_n_247__40_,r_n_247__39_,
  r_n_247__38_,r_n_247__37_,r_n_247__36_,r_n_247__35_,r_n_247__34_,r_n_247__33_,
  r_n_247__32_,r_n_247__31_,r_n_247__30_,r_n_247__29_,r_n_247__28_,r_n_247__27_,
  r_n_247__26_,r_n_247__25_,r_n_247__24_,r_n_247__23_,r_n_247__22_,r_n_247__21_,r_n_247__20_,
  r_n_247__19_,r_n_247__18_,r_n_247__17_,r_n_247__16_,r_n_247__15_,r_n_247__14_,
  r_n_247__13_,r_n_247__12_,r_n_247__11_,r_n_247__10_,r_n_247__9_,r_n_247__8_,
  r_n_247__7_,r_n_247__6_,r_n_247__5_,r_n_247__4_,r_n_247__3_,r_n_247__2_,r_n_247__1_,
  r_n_247__0_,r_n_246__63_,r_n_246__62_,r_n_246__61_,r_n_246__60_,r_n_246__59_,
  r_n_246__58_,r_n_246__57_,r_n_246__56_,r_n_246__55_,r_n_246__54_,r_n_246__53_,
  r_n_246__52_,r_n_246__51_,r_n_246__50_,r_n_246__49_,r_n_246__48_,r_n_246__47_,
  r_n_246__46_,r_n_246__45_,r_n_246__44_,r_n_246__43_,r_n_246__42_,r_n_246__41_,
  r_n_246__40_,r_n_246__39_,r_n_246__38_,r_n_246__37_,r_n_246__36_,r_n_246__35_,r_n_246__34_,
  r_n_246__33_,r_n_246__32_,r_n_246__31_,r_n_246__30_,r_n_246__29_,r_n_246__28_,
  r_n_246__27_,r_n_246__26_,r_n_246__25_,r_n_246__24_,r_n_246__23_,r_n_246__22_,
  r_n_246__21_,r_n_246__20_,r_n_246__19_,r_n_246__18_,r_n_246__17_,r_n_246__16_,
  r_n_246__15_,r_n_246__14_,r_n_246__13_,r_n_246__12_,r_n_246__11_,r_n_246__10_,
  r_n_246__9_,r_n_246__8_,r_n_246__7_,r_n_246__6_,r_n_246__5_,r_n_246__4_,r_n_246__3_,
  r_n_246__2_,r_n_246__1_,r_n_246__0_,r_n_245__63_,r_n_245__62_,r_n_245__61_,
  r_n_245__60_,r_n_245__59_,r_n_245__58_,r_n_245__57_,r_n_245__56_,r_n_245__55_,
  r_n_245__54_,r_n_245__53_,r_n_245__52_,r_n_245__51_,r_n_245__50_,r_n_245__49_,r_n_245__48_,
  r_n_245__47_,r_n_245__46_,r_n_245__45_,r_n_245__44_,r_n_245__43_,r_n_245__42_,
  r_n_245__41_,r_n_245__40_,r_n_245__39_,r_n_245__38_,r_n_245__37_,r_n_245__36_,
  r_n_245__35_,r_n_245__34_,r_n_245__33_,r_n_245__32_,r_n_245__31_,r_n_245__30_,
  r_n_245__29_,r_n_245__28_,r_n_245__27_,r_n_245__26_,r_n_245__25_,r_n_245__24_,
  r_n_245__23_,r_n_245__22_,r_n_245__21_,r_n_245__20_,r_n_245__19_,r_n_245__18_,
  r_n_245__17_,r_n_245__16_,r_n_245__15_,r_n_245__14_,r_n_245__13_,r_n_245__12_,
  r_n_245__11_,r_n_245__10_,r_n_245__9_,r_n_245__8_,r_n_245__7_,r_n_245__6_,r_n_245__5_,
  r_n_245__4_,r_n_245__3_,r_n_245__2_,r_n_245__1_,r_n_245__0_,r_n_244__63_,r_n_244__62_,
  r_n_244__61_,r_n_244__60_,r_n_244__59_,r_n_244__58_,r_n_244__57_,r_n_244__56_,
  r_n_244__55_,r_n_244__54_,r_n_244__53_,r_n_244__52_,r_n_244__51_,r_n_244__50_,
  r_n_244__49_,r_n_244__48_,r_n_244__47_,r_n_244__46_,r_n_244__45_,r_n_244__44_,
  r_n_244__43_,r_n_244__42_,r_n_244__41_,r_n_244__40_,r_n_244__39_,r_n_244__38_,
  r_n_244__37_,r_n_244__36_,r_n_244__35_,r_n_244__34_,r_n_244__33_,r_n_244__32_,
  r_n_244__31_,r_n_244__30_,r_n_244__29_,r_n_244__28_,r_n_244__27_,r_n_244__26_,
  r_n_244__25_,r_n_244__24_,r_n_244__23_,r_n_244__22_,r_n_244__21_,r_n_244__20_,r_n_244__19_,
  r_n_244__18_,r_n_244__17_,r_n_244__16_,r_n_244__15_,r_n_244__14_,r_n_244__13_,
  r_n_244__12_,r_n_244__11_,r_n_244__10_,r_n_244__9_,r_n_244__8_,r_n_244__7_,
  r_n_244__6_,r_n_244__5_,r_n_244__4_,r_n_244__3_,r_n_244__2_,r_n_244__1_,r_n_244__0_,
  r_n_243__63_,r_n_243__62_,r_n_243__61_,r_n_243__60_,r_n_243__59_,r_n_243__58_,
  r_n_243__57_,r_n_243__56_,r_n_243__55_,r_n_243__54_,r_n_243__53_,r_n_243__52_,
  r_n_243__51_,r_n_243__50_,r_n_243__49_,r_n_243__48_,r_n_243__47_,r_n_243__46_,
  r_n_243__45_,r_n_243__44_,r_n_243__43_,r_n_243__42_,r_n_243__41_,r_n_243__40_,
  r_n_243__39_,r_n_243__38_,r_n_243__37_,r_n_243__36_,r_n_243__35_,r_n_243__34_,r_n_243__33_,
  r_n_243__32_,r_n_243__31_,r_n_243__30_,r_n_243__29_,r_n_243__28_,r_n_243__27_,
  r_n_243__26_,r_n_243__25_,r_n_243__24_,r_n_243__23_,r_n_243__22_,r_n_243__21_,
  r_n_243__20_,r_n_243__19_,r_n_243__18_,r_n_243__17_,r_n_243__16_,r_n_243__15_,
  r_n_243__14_,r_n_243__13_,r_n_243__12_,r_n_243__11_,r_n_243__10_,r_n_243__9_,
  r_n_243__8_,r_n_243__7_,r_n_243__6_,r_n_243__5_,r_n_243__4_,r_n_243__3_,r_n_243__2_,
  r_n_243__1_,r_n_243__0_,r_n_242__63_,r_n_242__62_,r_n_242__61_,r_n_242__60_,
  r_n_242__59_,r_n_242__58_,r_n_242__57_,r_n_242__56_,r_n_242__55_,r_n_242__54_,
  r_n_242__53_,r_n_242__52_,r_n_242__51_,r_n_242__50_,r_n_242__49_,r_n_242__48_,r_n_242__47_,
  r_n_242__46_,r_n_242__45_,r_n_242__44_,r_n_242__43_,r_n_242__42_,r_n_242__41_,
  r_n_242__40_,r_n_242__39_,r_n_242__38_,r_n_242__37_,r_n_242__36_,r_n_242__35_,
  r_n_242__34_,r_n_242__33_,r_n_242__32_,r_n_242__31_,r_n_242__30_,r_n_242__29_,
  r_n_242__28_,r_n_242__27_,r_n_242__26_,r_n_242__25_,r_n_242__24_,r_n_242__23_,
  r_n_242__22_,r_n_242__21_,r_n_242__20_,r_n_242__19_,r_n_242__18_,r_n_242__17_,
  r_n_242__16_,r_n_242__15_,r_n_242__14_,r_n_242__13_,r_n_242__12_,r_n_242__11_,r_n_242__10_,
  r_n_242__9_,r_n_242__8_,r_n_242__7_,r_n_242__6_,r_n_242__5_,r_n_242__4_,
  r_n_242__3_,r_n_242__2_,r_n_242__1_,r_n_242__0_,r_n_241__63_,r_n_241__62_,r_n_241__61_,
  r_n_241__60_,r_n_241__59_,r_n_241__58_,r_n_241__57_,r_n_241__56_,r_n_241__55_,
  r_n_241__54_,r_n_241__53_,r_n_241__52_,r_n_241__51_,r_n_241__50_,r_n_241__49_,
  r_n_241__48_,r_n_241__47_,r_n_241__46_,r_n_241__45_,r_n_241__44_,r_n_241__43_,
  r_n_241__42_,r_n_241__41_,r_n_241__40_,r_n_241__39_,r_n_241__38_,r_n_241__37_,
  r_n_241__36_,r_n_241__35_,r_n_241__34_,r_n_241__33_,r_n_241__32_,r_n_241__31_,
  r_n_241__30_,r_n_241__29_,r_n_241__28_,r_n_241__27_,r_n_241__26_,r_n_241__25_,r_n_241__24_,
  r_n_241__23_,r_n_241__22_,r_n_241__21_,r_n_241__20_,r_n_241__19_,r_n_241__18_,
  r_n_241__17_,r_n_241__16_,r_n_241__15_,r_n_241__14_,r_n_241__13_,r_n_241__12_,
  r_n_241__11_,r_n_241__10_,r_n_241__9_,r_n_241__8_,r_n_241__7_,r_n_241__6_,
  r_n_241__5_,r_n_241__4_,r_n_241__3_,r_n_241__2_,r_n_241__1_,r_n_241__0_,r_n_256__63_,
  r_n_256__62_,r_n_256__61_,r_n_256__60_,r_n_256__59_,r_n_256__58_,r_n_256__57_,
  r_n_256__56_,r_n_256__55_,r_n_256__54_,r_n_256__53_,r_n_256__52_,r_n_256__51_,
  r_n_256__50_,r_n_256__49_,r_n_256__48_,r_n_256__47_,r_n_256__46_,r_n_256__45_,
  r_n_256__44_,r_n_256__43_,r_n_256__42_,r_n_256__41_,r_n_256__40_,r_n_256__39_,r_n_256__38_,
  r_n_256__37_,r_n_256__36_,r_n_256__35_,r_n_256__34_,r_n_256__33_,r_n_256__32_,
  r_n_256__31_,r_n_256__30_,r_n_256__29_,r_n_256__28_,r_n_256__27_,r_n_256__26_,
  r_n_256__25_,r_n_256__24_,r_n_256__23_,r_n_256__22_,r_n_256__21_,r_n_256__20_,
  r_n_256__19_,r_n_256__18_,r_n_256__17_,r_n_256__16_,r_n_256__15_,r_n_256__14_,
  r_n_256__13_,r_n_256__12_,r_n_256__11_,r_n_256__10_,r_n_256__9_,r_n_256__8_,r_n_256__7_,
  r_n_256__6_,r_n_256__5_,r_n_256__4_,r_n_256__3_,r_n_256__2_,r_n_256__1_,
  r_n_256__0_,r_n_255__63_,r_n_255__62_,r_n_255__61_,r_n_255__60_,r_n_255__59_,
  r_n_255__58_,r_n_255__57_,r_n_255__56_,r_n_255__55_,r_n_255__54_,r_n_255__53_,r_n_255__52_,
  r_n_255__51_,r_n_255__50_,r_n_255__49_,r_n_255__48_,r_n_255__47_,r_n_255__46_,
  r_n_255__45_,r_n_255__44_,r_n_255__43_,r_n_255__42_,r_n_255__41_,r_n_255__40_,
  r_n_255__39_,r_n_255__38_,r_n_255__37_,r_n_255__36_,r_n_255__35_,r_n_255__34_,
  r_n_255__33_,r_n_255__32_,r_n_255__31_,r_n_255__30_,r_n_255__29_,r_n_255__28_,
  r_n_255__27_,r_n_255__26_,r_n_255__25_,r_n_255__24_,r_n_255__23_,r_n_255__22_,
  r_n_255__21_,r_n_255__20_,r_n_255__19_,r_n_255__18_,r_n_255__17_,r_n_255__16_,
  r_n_255__15_,r_n_255__14_,r_n_255__13_,r_n_255__12_,r_n_255__11_,r_n_255__10_,r_n_255__9_,
  r_n_255__8_,r_n_255__7_,r_n_255__6_,r_n_255__5_,r_n_255__4_,r_n_255__3_,
  r_n_255__2_,r_n_255__1_,r_n_255__0_,r_n_254__63_,r_n_254__62_,r_n_254__61_,r_n_254__60_,
  r_n_254__59_,r_n_254__58_,r_n_254__57_,r_n_254__56_,r_n_254__55_,r_n_254__54_,
  r_n_254__53_,r_n_254__52_,r_n_254__51_,r_n_254__50_,r_n_254__49_,r_n_254__48_,
  r_n_254__47_,r_n_254__46_,r_n_254__45_,r_n_254__44_,r_n_254__43_,r_n_254__42_,
  r_n_254__41_,r_n_254__40_,r_n_254__39_,r_n_254__38_,r_n_254__37_,r_n_254__36_,
  r_n_254__35_,r_n_254__34_,r_n_254__33_,r_n_254__32_,r_n_254__31_,r_n_254__30_,
  r_n_254__29_,r_n_254__28_,r_n_254__27_,r_n_254__26_,r_n_254__25_,r_n_254__24_,r_n_254__23_,
  r_n_254__22_,r_n_254__21_,r_n_254__20_,r_n_254__19_,r_n_254__18_,r_n_254__17_,
  r_n_254__16_,r_n_254__15_,r_n_254__14_,r_n_254__13_,r_n_254__12_,r_n_254__11_,
  r_n_254__10_,r_n_254__9_,r_n_254__8_,r_n_254__7_,r_n_254__6_,r_n_254__5_,r_n_254__4_,
  r_n_254__3_,r_n_254__2_,r_n_254__1_,r_n_254__0_,r_n_253__63_,r_n_253__62_,
  r_n_253__61_,r_n_253__60_,r_n_253__59_,r_n_253__58_,r_n_253__57_,r_n_253__56_,
  r_n_253__55_,r_n_253__54_,r_n_253__53_,r_n_253__52_,r_n_253__51_,r_n_253__50_,
  r_n_253__49_,r_n_253__48_,r_n_253__47_,r_n_253__46_,r_n_253__45_,r_n_253__44_,
  r_n_253__43_,r_n_253__42_,r_n_253__41_,r_n_253__40_,r_n_253__39_,r_n_253__38_,r_n_253__37_,
  r_n_253__36_,r_n_253__35_,r_n_253__34_,r_n_253__33_,r_n_253__32_,r_n_253__31_,
  r_n_253__30_,r_n_253__29_,r_n_253__28_,r_n_253__27_,r_n_253__26_,r_n_253__25_,
  r_n_253__24_,r_n_253__23_,r_n_253__22_,r_n_253__21_,r_n_253__20_,r_n_253__19_,
  r_n_253__18_,r_n_253__17_,r_n_253__16_,r_n_253__15_,r_n_253__14_,r_n_253__13_,
  r_n_253__12_,r_n_253__11_,r_n_253__10_,r_n_253__9_,r_n_253__8_,r_n_253__7_,r_n_253__6_,
  r_n_253__5_,r_n_253__4_,r_n_253__3_,r_n_253__2_,r_n_253__1_,r_n_253__0_,
  r_n_252__63_,r_n_252__62_,r_n_252__61_,r_n_252__60_,r_n_252__59_,r_n_252__58_,
  r_n_252__57_,r_n_252__56_,r_n_252__55_,r_n_252__54_,r_n_252__53_,r_n_252__52_,r_n_252__51_,
  r_n_252__50_,r_n_252__49_,r_n_252__48_,r_n_252__47_,r_n_252__46_,r_n_252__45_,
  r_n_252__44_,r_n_252__43_,r_n_252__42_,r_n_252__41_,r_n_252__40_,r_n_252__39_,
  r_n_252__38_,r_n_252__37_,r_n_252__36_,r_n_252__35_,r_n_252__34_,r_n_252__33_,
  r_n_252__32_,r_n_252__31_,r_n_252__30_,r_n_252__29_,r_n_252__28_,r_n_252__27_,
  r_n_252__26_,r_n_252__25_,r_n_252__24_,r_n_252__23_,r_n_252__22_,r_n_252__21_,
  r_n_252__20_,r_n_252__19_,r_n_252__18_,r_n_252__17_,r_n_252__16_,r_n_252__15_,r_n_252__14_,
  r_n_252__13_,r_n_252__12_,r_n_252__11_,r_n_252__10_,r_n_252__9_,r_n_252__8_,
  r_n_252__7_,r_n_252__6_,r_n_252__5_,r_n_252__4_,r_n_252__3_,r_n_252__2_,r_n_252__1_,
  r_n_252__0_,r_n_251__63_,r_n_251__62_,r_n_251__61_,r_n_251__60_,r_n_251__59_,
  r_n_251__58_,r_n_251__57_,r_n_251__56_,r_n_251__55_,r_n_251__54_,r_n_251__53_,
  r_n_251__52_,r_n_251__51_,r_n_251__50_,r_n_251__49_,r_n_251__48_,r_n_251__47_,
  r_n_251__46_,r_n_251__45_,r_n_251__44_,r_n_251__43_,r_n_251__42_,r_n_251__41_,
  r_n_251__40_,r_n_251__39_,r_n_251__38_,r_n_251__37_,r_n_251__36_,r_n_251__35_,
  r_n_251__34_,r_n_251__33_,r_n_251__32_,r_n_251__31_,r_n_251__30_,r_n_251__29_,r_n_251__28_,
  r_n_251__27_,r_n_251__26_,r_n_251__25_,r_n_251__24_,r_n_251__23_,r_n_251__22_,
  r_n_251__21_,r_n_251__20_,r_n_251__19_,r_n_251__18_,r_n_251__17_,r_n_251__16_,
  r_n_251__15_,r_n_251__14_,r_n_251__13_,r_n_251__12_,r_n_251__11_,r_n_251__10_,
  r_n_251__9_,r_n_251__8_,r_n_251__7_,r_n_251__6_,r_n_251__5_,r_n_251__4_,r_n_251__3_,
  r_n_251__2_,r_n_251__1_,r_n_251__0_,r_n_250__63_,r_n_250__62_,r_n_250__61_,
  r_n_250__60_,r_n_250__59_,r_n_250__58_,r_n_250__57_,r_n_250__56_,r_n_250__55_,
  r_n_250__54_,r_n_250__53_,r_n_250__52_,r_n_250__51_,r_n_250__50_,r_n_250__49_,
  r_n_250__48_,r_n_250__47_,r_n_250__46_,r_n_250__45_,r_n_250__44_,r_n_250__43_,r_n_250__42_,
  r_n_250__41_,r_n_250__40_,r_n_250__39_,r_n_250__38_,r_n_250__37_,r_n_250__36_,
  r_n_250__35_,r_n_250__34_,r_n_250__33_,r_n_250__32_,r_n_250__31_,r_n_250__30_,
  r_n_250__29_,r_n_250__28_,r_n_250__27_,r_n_250__26_,r_n_250__25_,r_n_250__24_,
  r_n_250__23_,r_n_250__22_,r_n_250__21_,r_n_250__20_,r_n_250__19_,r_n_250__18_,
  r_n_250__17_,r_n_250__16_,r_n_250__15_,r_n_250__14_,r_n_250__13_,r_n_250__12_,
  r_n_250__11_,r_n_250__10_,r_n_250__9_,r_n_250__8_,r_n_250__7_,r_n_250__6_,r_n_250__5_,
  r_n_250__4_,r_n_250__3_,r_n_250__2_,r_n_250__1_,r_n_250__0_,r_n_249__63_,
  r_n_249__62_,r_n_249__61_,r_n_249__60_,r_n_249__59_,r_n_249__58_,r_n_249__57_,r_n_249__56_,
  r_n_249__55_,r_n_249__54_,r_n_249__53_,r_n_249__52_,r_n_249__51_,r_n_249__50_,
  r_n_249__49_,r_n_249__48_,r_n_249__47_,r_n_249__46_,r_n_249__45_,r_n_249__44_,
  r_n_249__43_,r_n_249__42_,r_n_249__41_,r_n_249__40_,r_n_249__39_,r_n_249__38_,
  r_n_249__37_,r_n_249__36_,r_n_249__35_,r_n_249__34_,r_n_249__33_,r_n_249__32_,
  r_n_249__31_,r_n_249__30_,r_n_249__29_,r_n_249__28_,r_n_249__27_,r_n_249__26_,
  r_n_249__25_,r_n_249__24_,r_n_249__23_,r_n_249__22_,r_n_249__21_,r_n_249__20_,
  r_n_249__19_,r_n_249__18_,r_n_249__17_,r_n_249__16_,r_n_249__15_,r_n_249__14_,r_n_249__13_,
  r_n_249__12_,r_n_249__11_,r_n_249__10_,r_n_249__9_,r_n_249__8_,r_n_249__7_,
  r_n_249__6_,r_n_249__5_,r_n_249__4_,r_n_249__3_,r_n_249__2_,r_n_249__1_,r_n_249__0_,
  r_n_264__63_,r_n_264__62_,r_n_264__61_,r_n_264__60_,r_n_264__59_,r_n_264__58_,
  r_n_264__57_,r_n_264__56_,r_n_264__55_,r_n_264__54_,r_n_264__53_,r_n_264__52_,
  r_n_264__51_,r_n_264__50_,r_n_264__49_,r_n_264__48_,r_n_264__47_,r_n_264__46_,
  r_n_264__45_,r_n_264__44_,r_n_264__43_,r_n_264__42_,r_n_264__41_,r_n_264__40_,
  r_n_264__39_,r_n_264__38_,r_n_264__37_,r_n_264__36_,r_n_264__35_,r_n_264__34_,
  r_n_264__33_,r_n_264__32_,r_n_264__31_,r_n_264__30_,r_n_264__29_,r_n_264__28_,r_n_264__27_,
  r_n_264__26_,r_n_264__25_,r_n_264__24_,r_n_264__23_,r_n_264__22_,r_n_264__21_,
  r_n_264__20_,r_n_264__19_,r_n_264__18_,r_n_264__17_,r_n_264__16_,r_n_264__15_,
  r_n_264__14_,r_n_264__13_,r_n_264__12_,r_n_264__11_,r_n_264__10_,r_n_264__9_,
  r_n_264__8_,r_n_264__7_,r_n_264__6_,r_n_264__5_,r_n_264__4_,r_n_264__3_,r_n_264__2_,
  r_n_264__1_,r_n_264__0_,r_n_263__63_,r_n_263__62_,r_n_263__61_,r_n_263__60_,
  r_n_263__59_,r_n_263__58_,r_n_263__57_,r_n_263__56_,r_n_263__55_,r_n_263__54_,
  r_n_263__53_,r_n_263__52_,r_n_263__51_,r_n_263__50_,r_n_263__49_,r_n_263__48_,
  r_n_263__47_,r_n_263__46_,r_n_263__45_,r_n_263__44_,r_n_263__43_,r_n_263__42_,r_n_263__41_,
  r_n_263__40_,r_n_263__39_,r_n_263__38_,r_n_263__37_,r_n_263__36_,r_n_263__35_,
  r_n_263__34_,r_n_263__33_,r_n_263__32_,r_n_263__31_,r_n_263__30_,r_n_263__29_,
  r_n_263__28_,r_n_263__27_,r_n_263__26_,r_n_263__25_,r_n_263__24_,r_n_263__23_,
  r_n_263__22_,r_n_263__21_,r_n_263__20_,r_n_263__19_,r_n_263__18_,r_n_263__17_,
  r_n_263__16_,r_n_263__15_,r_n_263__14_,r_n_263__13_,r_n_263__12_,r_n_263__11_,
  r_n_263__10_,r_n_263__9_,r_n_263__8_,r_n_263__7_,r_n_263__6_,r_n_263__5_,r_n_263__4_,
  r_n_263__3_,r_n_263__2_,r_n_263__1_,r_n_263__0_,r_n_262__63_,r_n_262__62_,
  r_n_262__61_,r_n_262__60_,r_n_262__59_,r_n_262__58_,r_n_262__57_,r_n_262__56_,r_n_262__55_,
  r_n_262__54_,r_n_262__53_,r_n_262__52_,r_n_262__51_,r_n_262__50_,r_n_262__49_,
  r_n_262__48_,r_n_262__47_,r_n_262__46_,r_n_262__45_,r_n_262__44_,r_n_262__43_,
  r_n_262__42_,r_n_262__41_,r_n_262__40_,r_n_262__39_,r_n_262__38_,r_n_262__37_,
  r_n_262__36_,r_n_262__35_,r_n_262__34_,r_n_262__33_,r_n_262__32_,r_n_262__31_,
  r_n_262__30_,r_n_262__29_,r_n_262__28_,r_n_262__27_,r_n_262__26_,r_n_262__25_,
  r_n_262__24_,r_n_262__23_,r_n_262__22_,r_n_262__21_,r_n_262__20_,r_n_262__19_,r_n_262__18_,
  r_n_262__17_,r_n_262__16_,r_n_262__15_,r_n_262__14_,r_n_262__13_,r_n_262__12_,
  r_n_262__11_,r_n_262__10_,r_n_262__9_,r_n_262__8_,r_n_262__7_,r_n_262__6_,
  r_n_262__5_,r_n_262__4_,r_n_262__3_,r_n_262__2_,r_n_262__1_,r_n_262__0_,r_n_261__63_,
  r_n_261__62_,r_n_261__61_,r_n_261__60_,r_n_261__59_,r_n_261__58_,r_n_261__57_,
  r_n_261__56_,r_n_261__55_,r_n_261__54_,r_n_261__53_,r_n_261__52_,r_n_261__51_,
  r_n_261__50_,r_n_261__49_,r_n_261__48_,r_n_261__47_,r_n_261__46_,r_n_261__45_,
  r_n_261__44_,r_n_261__43_,r_n_261__42_,r_n_261__41_,r_n_261__40_,r_n_261__39_,
  r_n_261__38_,r_n_261__37_,r_n_261__36_,r_n_261__35_,r_n_261__34_,r_n_261__33_,r_n_261__32_,
  r_n_261__31_,r_n_261__30_,r_n_261__29_,r_n_261__28_,r_n_261__27_,r_n_261__26_,
  r_n_261__25_,r_n_261__24_,r_n_261__23_,r_n_261__22_,r_n_261__21_,r_n_261__20_,
  r_n_261__19_,r_n_261__18_,r_n_261__17_,r_n_261__16_,r_n_261__15_,r_n_261__14_,
  r_n_261__13_,r_n_261__12_,r_n_261__11_,r_n_261__10_,r_n_261__9_,r_n_261__8_,
  r_n_261__7_,r_n_261__6_,r_n_261__5_,r_n_261__4_,r_n_261__3_,r_n_261__2_,r_n_261__1_,
  r_n_261__0_,r_n_260__63_,r_n_260__62_,r_n_260__61_,r_n_260__60_,r_n_260__59_,
  r_n_260__58_,r_n_260__57_,r_n_260__56_,r_n_260__55_,r_n_260__54_,r_n_260__53_,
  r_n_260__52_,r_n_260__51_,r_n_260__50_,r_n_260__49_,r_n_260__48_,r_n_260__47_,r_n_260__46_,
  r_n_260__45_,r_n_260__44_,r_n_260__43_,r_n_260__42_,r_n_260__41_,r_n_260__40_,
  r_n_260__39_,r_n_260__38_,r_n_260__37_,r_n_260__36_,r_n_260__35_,r_n_260__34_,
  r_n_260__33_,r_n_260__32_,r_n_260__31_,r_n_260__30_,r_n_260__29_,r_n_260__28_,
  r_n_260__27_,r_n_260__26_,r_n_260__25_,r_n_260__24_,r_n_260__23_,r_n_260__22_,
  r_n_260__21_,r_n_260__20_,r_n_260__19_,r_n_260__18_,r_n_260__17_,r_n_260__16_,
  r_n_260__15_,r_n_260__14_,r_n_260__13_,r_n_260__12_,r_n_260__11_,r_n_260__10_,r_n_260__9_,
  r_n_260__8_,r_n_260__7_,r_n_260__6_,r_n_260__5_,r_n_260__4_,r_n_260__3_,
  r_n_260__2_,r_n_260__1_,r_n_260__0_,r_n_259__63_,r_n_259__62_,r_n_259__61_,r_n_259__60_,
  r_n_259__59_,r_n_259__58_,r_n_259__57_,r_n_259__56_,r_n_259__55_,r_n_259__54_,
  r_n_259__53_,r_n_259__52_,r_n_259__51_,r_n_259__50_,r_n_259__49_,r_n_259__48_,
  r_n_259__47_,r_n_259__46_,r_n_259__45_,r_n_259__44_,r_n_259__43_,r_n_259__42_,
  r_n_259__41_,r_n_259__40_,r_n_259__39_,r_n_259__38_,r_n_259__37_,r_n_259__36_,
  r_n_259__35_,r_n_259__34_,r_n_259__33_,r_n_259__32_,r_n_259__31_,r_n_259__30_,
  r_n_259__29_,r_n_259__28_,r_n_259__27_,r_n_259__26_,r_n_259__25_,r_n_259__24_,
  r_n_259__23_,r_n_259__22_,r_n_259__21_,r_n_259__20_,r_n_259__19_,r_n_259__18_,r_n_259__17_,
  r_n_259__16_,r_n_259__15_,r_n_259__14_,r_n_259__13_,r_n_259__12_,r_n_259__11_,
  r_n_259__10_,r_n_259__9_,r_n_259__8_,r_n_259__7_,r_n_259__6_,r_n_259__5_,
  r_n_259__4_,r_n_259__3_,r_n_259__2_,r_n_259__1_,r_n_259__0_,r_n_258__63_,r_n_258__62_,
  r_n_258__61_,r_n_258__60_,r_n_258__59_,r_n_258__58_,r_n_258__57_,r_n_258__56_,
  r_n_258__55_,r_n_258__54_,r_n_258__53_,r_n_258__52_,r_n_258__51_,r_n_258__50_,
  r_n_258__49_,r_n_258__48_,r_n_258__47_,r_n_258__46_,r_n_258__45_,r_n_258__44_,
  r_n_258__43_,r_n_258__42_,r_n_258__41_,r_n_258__40_,r_n_258__39_,r_n_258__38_,
  r_n_258__37_,r_n_258__36_,r_n_258__35_,r_n_258__34_,r_n_258__33_,r_n_258__32_,r_n_258__31_,
  r_n_258__30_,r_n_258__29_,r_n_258__28_,r_n_258__27_,r_n_258__26_,r_n_258__25_,
  r_n_258__24_,r_n_258__23_,r_n_258__22_,r_n_258__21_,r_n_258__20_,r_n_258__19_,
  r_n_258__18_,r_n_258__17_,r_n_258__16_,r_n_258__15_,r_n_258__14_,r_n_258__13_,
  r_n_258__12_,r_n_258__11_,r_n_258__10_,r_n_258__9_,r_n_258__8_,r_n_258__7_,r_n_258__6_,
  r_n_258__5_,r_n_258__4_,r_n_258__3_,r_n_258__2_,r_n_258__1_,r_n_258__0_,
  r_n_257__63_,r_n_257__62_,r_n_257__61_,r_n_257__60_,r_n_257__59_,r_n_257__58_,
  r_n_257__57_,r_n_257__56_,r_n_257__55_,r_n_257__54_,r_n_257__53_,r_n_257__52_,
  r_n_257__51_,r_n_257__50_,r_n_257__49_,r_n_257__48_,r_n_257__47_,r_n_257__46_,r_n_257__45_,
  r_n_257__44_,r_n_257__43_,r_n_257__42_,r_n_257__41_,r_n_257__40_,r_n_257__39_,
  r_n_257__38_,r_n_257__37_,r_n_257__36_,r_n_257__35_,r_n_257__34_,r_n_257__33_,
  r_n_257__32_,r_n_257__31_,r_n_257__30_,r_n_257__29_,r_n_257__28_,r_n_257__27_,
  r_n_257__26_,r_n_257__25_,r_n_257__24_,r_n_257__23_,r_n_257__22_,r_n_257__21_,
  r_n_257__20_,r_n_257__19_,r_n_257__18_,r_n_257__17_,r_n_257__16_,r_n_257__15_,
  r_n_257__14_,r_n_257__13_,r_n_257__12_,r_n_257__11_,r_n_257__10_,r_n_257__9_,r_n_257__8_,
  r_n_257__7_,r_n_257__6_,r_n_257__5_,r_n_257__4_,r_n_257__3_,r_n_257__2_,
  r_n_257__1_,r_n_257__0_,r_n_272__63_,r_n_272__62_,r_n_272__61_,r_n_272__60_,r_n_272__59_,
  r_n_272__58_,r_n_272__57_,r_n_272__56_,r_n_272__55_,r_n_272__54_,r_n_272__53_,
  r_n_272__52_,r_n_272__51_,r_n_272__50_,r_n_272__49_,r_n_272__48_,r_n_272__47_,
  r_n_272__46_,r_n_272__45_,r_n_272__44_,r_n_272__43_,r_n_272__42_,r_n_272__41_,
  r_n_272__40_,r_n_272__39_,r_n_272__38_,r_n_272__37_,r_n_272__36_,r_n_272__35_,
  r_n_272__34_,r_n_272__33_,r_n_272__32_,r_n_272__31_,r_n_272__30_,r_n_272__29_,
  r_n_272__28_,r_n_272__27_,r_n_272__26_,r_n_272__25_,r_n_272__24_,r_n_272__23_,r_n_272__22_,
  r_n_272__21_,r_n_272__20_,r_n_272__19_,r_n_272__18_,r_n_272__17_,r_n_272__16_,
  r_n_272__15_,r_n_272__14_,r_n_272__13_,r_n_272__12_,r_n_272__11_,r_n_272__10_,
  r_n_272__9_,r_n_272__8_,r_n_272__7_,r_n_272__6_,r_n_272__5_,r_n_272__4_,r_n_272__3_,
  r_n_272__2_,r_n_272__1_,r_n_272__0_,r_n_271__63_,r_n_271__62_,r_n_271__61_,
  r_n_271__60_,r_n_271__59_,r_n_271__58_,r_n_271__57_,r_n_271__56_,r_n_271__55_,
  r_n_271__54_,r_n_271__53_,r_n_271__52_,r_n_271__51_,r_n_271__50_,r_n_271__49_,
  r_n_271__48_,r_n_271__47_,r_n_271__46_,r_n_271__45_,r_n_271__44_,r_n_271__43_,
  r_n_271__42_,r_n_271__41_,r_n_271__40_,r_n_271__39_,r_n_271__38_,r_n_271__37_,r_n_271__36_,
  r_n_271__35_,r_n_271__34_,r_n_271__33_,r_n_271__32_,r_n_271__31_,r_n_271__30_,
  r_n_271__29_,r_n_271__28_,r_n_271__27_,r_n_271__26_,r_n_271__25_,r_n_271__24_,
  r_n_271__23_,r_n_271__22_,r_n_271__21_,r_n_271__20_,r_n_271__19_,r_n_271__18_,
  r_n_271__17_,r_n_271__16_,r_n_271__15_,r_n_271__14_,r_n_271__13_,r_n_271__12_,
  r_n_271__11_,r_n_271__10_,r_n_271__9_,r_n_271__8_,r_n_271__7_,r_n_271__6_,r_n_271__5_,
  r_n_271__4_,r_n_271__3_,r_n_271__2_,r_n_271__1_,r_n_271__0_,r_n_270__63_,
  r_n_270__62_,r_n_270__61_,r_n_270__60_,r_n_270__59_,r_n_270__58_,r_n_270__57_,
  r_n_270__56_,r_n_270__55_,r_n_270__54_,r_n_270__53_,r_n_270__52_,r_n_270__51_,r_n_270__50_,
  r_n_270__49_,r_n_270__48_,r_n_270__47_,r_n_270__46_,r_n_270__45_,r_n_270__44_,
  r_n_270__43_,r_n_270__42_,r_n_270__41_,r_n_270__40_,r_n_270__39_,r_n_270__38_,
  r_n_270__37_,r_n_270__36_,r_n_270__35_,r_n_270__34_,r_n_270__33_,r_n_270__32_,
  r_n_270__31_,r_n_270__30_,r_n_270__29_,r_n_270__28_,r_n_270__27_,r_n_270__26_,
  r_n_270__25_,r_n_270__24_,r_n_270__23_,r_n_270__22_,r_n_270__21_,r_n_270__20_,
  r_n_270__19_,r_n_270__18_,r_n_270__17_,r_n_270__16_,r_n_270__15_,r_n_270__14_,
  r_n_270__13_,r_n_270__12_,r_n_270__11_,r_n_270__10_,r_n_270__9_,r_n_270__8_,r_n_270__7_,
  r_n_270__6_,r_n_270__5_,r_n_270__4_,r_n_270__3_,r_n_270__2_,r_n_270__1_,r_n_270__0_,
  r_n_269__63_,r_n_269__62_,r_n_269__61_,r_n_269__60_,r_n_269__59_,r_n_269__58_,
  r_n_269__57_,r_n_269__56_,r_n_269__55_,r_n_269__54_,r_n_269__53_,r_n_269__52_,
  r_n_269__51_,r_n_269__50_,r_n_269__49_,r_n_269__48_,r_n_269__47_,r_n_269__46_,
  r_n_269__45_,r_n_269__44_,r_n_269__43_,r_n_269__42_,r_n_269__41_,r_n_269__40_,
  r_n_269__39_,r_n_269__38_,r_n_269__37_,r_n_269__36_,r_n_269__35_,r_n_269__34_,
  r_n_269__33_,r_n_269__32_,r_n_269__31_,r_n_269__30_,r_n_269__29_,r_n_269__28_,
  r_n_269__27_,r_n_269__26_,r_n_269__25_,r_n_269__24_,r_n_269__23_,r_n_269__22_,r_n_269__21_,
  r_n_269__20_,r_n_269__19_,r_n_269__18_,r_n_269__17_,r_n_269__16_,r_n_269__15_,
  r_n_269__14_,r_n_269__13_,r_n_269__12_,r_n_269__11_,r_n_269__10_,r_n_269__9_,
  r_n_269__8_,r_n_269__7_,r_n_269__6_,r_n_269__5_,r_n_269__4_,r_n_269__3_,r_n_269__2_,
  r_n_269__1_,r_n_269__0_,r_n_268__63_,r_n_268__62_,r_n_268__61_,r_n_268__60_,
  r_n_268__59_,r_n_268__58_,r_n_268__57_,r_n_268__56_,r_n_268__55_,r_n_268__54_,
  r_n_268__53_,r_n_268__52_,r_n_268__51_,r_n_268__50_,r_n_268__49_,r_n_268__48_,
  r_n_268__47_,r_n_268__46_,r_n_268__45_,r_n_268__44_,r_n_268__43_,r_n_268__42_,
  r_n_268__41_,r_n_268__40_,r_n_268__39_,r_n_268__38_,r_n_268__37_,r_n_268__36_,r_n_268__35_,
  r_n_268__34_,r_n_268__33_,r_n_268__32_,r_n_268__31_,r_n_268__30_,r_n_268__29_,
  r_n_268__28_,r_n_268__27_,r_n_268__26_,r_n_268__25_,r_n_268__24_,r_n_268__23_,
  r_n_268__22_,r_n_268__21_,r_n_268__20_,r_n_268__19_,r_n_268__18_,r_n_268__17_,
  r_n_268__16_,r_n_268__15_,r_n_268__14_,r_n_268__13_,r_n_268__12_,r_n_268__11_,
  r_n_268__10_,r_n_268__9_,r_n_268__8_,r_n_268__7_,r_n_268__6_,r_n_268__5_,r_n_268__4_,
  r_n_268__3_,r_n_268__2_,r_n_268__1_,r_n_268__0_,r_n_267__63_,r_n_267__62_,
  r_n_267__61_,r_n_267__60_,r_n_267__59_,r_n_267__58_,r_n_267__57_,r_n_267__56_,
  r_n_267__55_,r_n_267__54_,r_n_267__53_,r_n_267__52_,r_n_267__51_,r_n_267__50_,r_n_267__49_,
  r_n_267__48_,r_n_267__47_,r_n_267__46_,r_n_267__45_,r_n_267__44_,r_n_267__43_,
  r_n_267__42_,r_n_267__41_,r_n_267__40_,r_n_267__39_,r_n_267__38_,r_n_267__37_,
  r_n_267__36_,r_n_267__35_,r_n_267__34_,r_n_267__33_,r_n_267__32_,r_n_267__31_,
  r_n_267__30_,r_n_267__29_,r_n_267__28_,r_n_267__27_,r_n_267__26_,r_n_267__25_,
  r_n_267__24_,r_n_267__23_,r_n_267__22_,r_n_267__21_,r_n_267__20_,r_n_267__19_,
  r_n_267__18_,r_n_267__17_,r_n_267__16_,r_n_267__15_,r_n_267__14_,r_n_267__13_,r_n_267__12_,
  r_n_267__11_,r_n_267__10_,r_n_267__9_,r_n_267__8_,r_n_267__7_,r_n_267__6_,
  r_n_267__5_,r_n_267__4_,r_n_267__3_,r_n_267__2_,r_n_267__1_,r_n_267__0_,r_n_266__63_,
  r_n_266__62_,r_n_266__61_,r_n_266__60_,r_n_266__59_,r_n_266__58_,r_n_266__57_,
  r_n_266__56_,r_n_266__55_,r_n_266__54_,r_n_266__53_,r_n_266__52_,r_n_266__51_,
  r_n_266__50_,r_n_266__49_,r_n_266__48_,r_n_266__47_,r_n_266__46_,r_n_266__45_,
  r_n_266__44_,r_n_266__43_,r_n_266__42_,r_n_266__41_,r_n_266__40_,r_n_266__39_,
  r_n_266__38_,r_n_266__37_,r_n_266__36_,r_n_266__35_,r_n_266__34_,r_n_266__33_,
  r_n_266__32_,r_n_266__31_,r_n_266__30_,r_n_266__29_,r_n_266__28_,r_n_266__27_,r_n_266__26_,
  r_n_266__25_,r_n_266__24_,r_n_266__23_,r_n_266__22_,r_n_266__21_,r_n_266__20_,
  r_n_266__19_,r_n_266__18_,r_n_266__17_,r_n_266__16_,r_n_266__15_,r_n_266__14_,
  r_n_266__13_,r_n_266__12_,r_n_266__11_,r_n_266__10_,r_n_266__9_,r_n_266__8_,
  r_n_266__7_,r_n_266__6_,r_n_266__5_,r_n_266__4_,r_n_266__3_,r_n_266__2_,r_n_266__1_,
  r_n_266__0_,r_n_265__63_,r_n_265__62_,r_n_265__61_,r_n_265__60_,r_n_265__59_,
  r_n_265__58_,r_n_265__57_,r_n_265__56_,r_n_265__55_,r_n_265__54_,r_n_265__53_,
  r_n_265__52_,r_n_265__51_,r_n_265__50_,r_n_265__49_,r_n_265__48_,r_n_265__47_,
  r_n_265__46_,r_n_265__45_,r_n_265__44_,r_n_265__43_,r_n_265__42_,r_n_265__41_,r_n_265__40_,
  r_n_265__39_,r_n_265__38_,r_n_265__37_,r_n_265__36_,r_n_265__35_,r_n_265__34_,
  r_n_265__33_,r_n_265__32_,r_n_265__31_,r_n_265__30_,r_n_265__29_,r_n_265__28_,
  r_n_265__27_,r_n_265__26_,r_n_265__25_,r_n_265__24_,r_n_265__23_,r_n_265__22_,
  r_n_265__21_,r_n_265__20_,r_n_265__19_,r_n_265__18_,r_n_265__17_,r_n_265__16_,
  r_n_265__15_,r_n_265__14_,r_n_265__13_,r_n_265__12_,r_n_265__11_,r_n_265__10_,
  r_n_265__9_,r_n_265__8_,r_n_265__7_,r_n_265__6_,r_n_265__5_,r_n_265__4_,r_n_265__3_,
  r_n_265__2_,r_n_265__1_,r_n_265__0_,r_n_280__63_,r_n_280__62_,r_n_280__61_,
  r_n_280__60_,r_n_280__59_,r_n_280__58_,r_n_280__57_,r_n_280__56_,r_n_280__55_,r_n_280__54_,
  r_n_280__53_,r_n_280__52_,r_n_280__51_,r_n_280__50_,r_n_280__49_,r_n_280__48_,
  r_n_280__47_,r_n_280__46_,r_n_280__45_,r_n_280__44_,r_n_280__43_,r_n_280__42_,
  r_n_280__41_,r_n_280__40_,r_n_280__39_,r_n_280__38_,r_n_280__37_,r_n_280__36_,
  r_n_280__35_,r_n_280__34_,r_n_280__33_,r_n_280__32_,r_n_280__31_,r_n_280__30_,
  r_n_280__29_,r_n_280__28_,r_n_280__27_,r_n_280__26_,r_n_280__25_,r_n_280__24_,
  r_n_280__23_,r_n_280__22_,r_n_280__21_,r_n_280__20_,r_n_280__19_,r_n_280__18_,
  r_n_280__17_,r_n_280__16_,r_n_280__15_,r_n_280__14_,r_n_280__13_,r_n_280__12_,r_n_280__11_,
  r_n_280__10_,r_n_280__9_,r_n_280__8_,r_n_280__7_,r_n_280__6_,r_n_280__5_,
  r_n_280__4_,r_n_280__3_,r_n_280__2_,r_n_280__1_,r_n_280__0_,r_n_279__63_,r_n_279__62_,
  r_n_279__61_,r_n_279__60_,r_n_279__59_,r_n_279__58_,r_n_279__57_,r_n_279__56_,
  r_n_279__55_,r_n_279__54_,r_n_279__53_,r_n_279__52_,r_n_279__51_,r_n_279__50_,
  r_n_279__49_,r_n_279__48_,r_n_279__47_,r_n_279__46_,r_n_279__45_,r_n_279__44_,
  r_n_279__43_,r_n_279__42_,r_n_279__41_,r_n_279__40_,r_n_279__39_,r_n_279__38_,
  r_n_279__37_,r_n_279__36_,r_n_279__35_,r_n_279__34_,r_n_279__33_,r_n_279__32_,
  r_n_279__31_,r_n_279__30_,r_n_279__29_,r_n_279__28_,r_n_279__27_,r_n_279__26_,r_n_279__25_,
  r_n_279__24_,r_n_279__23_,r_n_279__22_,r_n_279__21_,r_n_279__20_,r_n_279__19_,
  r_n_279__18_,r_n_279__17_,r_n_279__16_,r_n_279__15_,r_n_279__14_,r_n_279__13_,
  r_n_279__12_,r_n_279__11_,r_n_279__10_,r_n_279__9_,r_n_279__8_,r_n_279__7_,
  r_n_279__6_,r_n_279__5_,r_n_279__4_,r_n_279__3_,r_n_279__2_,r_n_279__1_,r_n_279__0_,
  r_n_278__63_,r_n_278__62_,r_n_278__61_,r_n_278__60_,r_n_278__59_,r_n_278__58_,
  r_n_278__57_,r_n_278__56_,r_n_278__55_,r_n_278__54_,r_n_278__53_,r_n_278__52_,
  r_n_278__51_,r_n_278__50_,r_n_278__49_,r_n_278__48_,r_n_278__47_,r_n_278__46_,
  r_n_278__45_,r_n_278__44_,r_n_278__43_,r_n_278__42_,r_n_278__41_,r_n_278__40_,r_n_278__39_,
  r_n_278__38_,r_n_278__37_,r_n_278__36_,r_n_278__35_,r_n_278__34_,r_n_278__33_,
  r_n_278__32_,r_n_278__31_,r_n_278__30_,r_n_278__29_,r_n_278__28_,r_n_278__27_,
  r_n_278__26_,r_n_278__25_,r_n_278__24_,r_n_278__23_,r_n_278__22_,r_n_278__21_,
  r_n_278__20_,r_n_278__19_,r_n_278__18_,r_n_278__17_,r_n_278__16_,r_n_278__15_,
  r_n_278__14_,r_n_278__13_,r_n_278__12_,r_n_278__11_,r_n_278__10_,r_n_278__9_,r_n_278__8_,
  r_n_278__7_,r_n_278__6_,r_n_278__5_,r_n_278__4_,r_n_278__3_,r_n_278__2_,
  r_n_278__1_,r_n_278__0_,r_n_277__63_,r_n_277__62_,r_n_277__61_,r_n_277__60_,
  r_n_277__59_,r_n_277__58_,r_n_277__57_,r_n_277__56_,r_n_277__55_,r_n_277__54_,r_n_277__53_,
  r_n_277__52_,r_n_277__51_,r_n_277__50_,r_n_277__49_,r_n_277__48_,r_n_277__47_,
  r_n_277__46_,r_n_277__45_,r_n_277__44_,r_n_277__43_,r_n_277__42_,r_n_277__41_,
  r_n_277__40_,r_n_277__39_,r_n_277__38_,r_n_277__37_,r_n_277__36_,r_n_277__35_,
  r_n_277__34_,r_n_277__33_,r_n_277__32_,r_n_277__31_,r_n_277__30_,r_n_277__29_,
  r_n_277__28_,r_n_277__27_,r_n_277__26_,r_n_277__25_,r_n_277__24_,r_n_277__23_,
  r_n_277__22_,r_n_277__21_,r_n_277__20_,r_n_277__19_,r_n_277__18_,r_n_277__17_,r_n_277__16_,
  r_n_277__15_,r_n_277__14_,r_n_277__13_,r_n_277__12_,r_n_277__11_,r_n_277__10_,
  r_n_277__9_,r_n_277__8_,r_n_277__7_,r_n_277__6_,r_n_277__5_,r_n_277__4_,
  r_n_277__3_,r_n_277__2_,r_n_277__1_,r_n_277__0_,r_n_276__63_,r_n_276__62_,r_n_276__61_,
  r_n_276__60_,r_n_276__59_,r_n_276__58_,r_n_276__57_,r_n_276__56_,r_n_276__55_,
  r_n_276__54_,r_n_276__53_,r_n_276__52_,r_n_276__51_,r_n_276__50_,r_n_276__49_,
  r_n_276__48_,r_n_276__47_,r_n_276__46_,r_n_276__45_,r_n_276__44_,r_n_276__43_,
  r_n_276__42_,r_n_276__41_,r_n_276__40_,r_n_276__39_,r_n_276__38_,r_n_276__37_,
  r_n_276__36_,r_n_276__35_,r_n_276__34_,r_n_276__33_,r_n_276__32_,r_n_276__31_,r_n_276__30_,
  r_n_276__29_,r_n_276__28_,r_n_276__27_,r_n_276__26_,r_n_276__25_,r_n_276__24_,
  r_n_276__23_,r_n_276__22_,r_n_276__21_,r_n_276__20_,r_n_276__19_,r_n_276__18_,
  r_n_276__17_,r_n_276__16_,r_n_276__15_,r_n_276__14_,r_n_276__13_,r_n_276__12_,
  r_n_276__11_,r_n_276__10_,r_n_276__9_,r_n_276__8_,r_n_276__7_,r_n_276__6_,r_n_276__5_,
  r_n_276__4_,r_n_276__3_,r_n_276__2_,r_n_276__1_,r_n_276__0_,r_n_275__63_,
  r_n_275__62_,r_n_275__61_,r_n_275__60_,r_n_275__59_,r_n_275__58_,r_n_275__57_,
  r_n_275__56_,r_n_275__55_,r_n_275__54_,r_n_275__53_,r_n_275__52_,r_n_275__51_,
  r_n_275__50_,r_n_275__49_,r_n_275__48_,r_n_275__47_,r_n_275__46_,r_n_275__45_,r_n_275__44_,
  r_n_275__43_,r_n_275__42_,r_n_275__41_,r_n_275__40_,r_n_275__39_,r_n_275__38_,
  r_n_275__37_,r_n_275__36_,r_n_275__35_,r_n_275__34_,r_n_275__33_,r_n_275__32_,
  r_n_275__31_,r_n_275__30_,r_n_275__29_,r_n_275__28_,r_n_275__27_,r_n_275__26_,
  r_n_275__25_,r_n_275__24_,r_n_275__23_,r_n_275__22_,r_n_275__21_,r_n_275__20_,
  r_n_275__19_,r_n_275__18_,r_n_275__17_,r_n_275__16_,r_n_275__15_,r_n_275__14_,
  r_n_275__13_,r_n_275__12_,r_n_275__11_,r_n_275__10_,r_n_275__9_,r_n_275__8_,r_n_275__7_,
  r_n_275__6_,r_n_275__5_,r_n_275__4_,r_n_275__3_,r_n_275__2_,r_n_275__1_,
  r_n_275__0_,r_n_274__63_,r_n_274__62_,r_n_274__61_,r_n_274__60_,r_n_274__59_,r_n_274__58_,
  r_n_274__57_,r_n_274__56_,r_n_274__55_,r_n_274__54_,r_n_274__53_,r_n_274__52_,
  r_n_274__51_,r_n_274__50_,r_n_274__49_,r_n_274__48_,r_n_274__47_,r_n_274__46_,
  r_n_274__45_,r_n_274__44_,r_n_274__43_,r_n_274__42_,r_n_274__41_,r_n_274__40_,
  r_n_274__39_,r_n_274__38_,r_n_274__37_,r_n_274__36_,r_n_274__35_,r_n_274__34_,
  r_n_274__33_,r_n_274__32_,r_n_274__31_,r_n_274__30_,r_n_274__29_,r_n_274__28_,
  r_n_274__27_,r_n_274__26_,r_n_274__25_,r_n_274__24_,r_n_274__23_,r_n_274__22_,
  r_n_274__21_,r_n_274__20_,r_n_274__19_,r_n_274__18_,r_n_274__17_,r_n_274__16_,r_n_274__15_,
  r_n_274__14_,r_n_274__13_,r_n_274__12_,r_n_274__11_,r_n_274__10_,r_n_274__9_,
  r_n_274__8_,r_n_274__7_,r_n_274__6_,r_n_274__5_,r_n_274__4_,r_n_274__3_,r_n_274__2_,
  r_n_274__1_,r_n_274__0_,r_n_273__63_,r_n_273__62_,r_n_273__61_,r_n_273__60_,
  r_n_273__59_,r_n_273__58_,r_n_273__57_,r_n_273__56_,r_n_273__55_,r_n_273__54_,
  r_n_273__53_,r_n_273__52_,r_n_273__51_,r_n_273__50_,r_n_273__49_,r_n_273__48_,
  r_n_273__47_,r_n_273__46_,r_n_273__45_,r_n_273__44_,r_n_273__43_,r_n_273__42_,
  r_n_273__41_,r_n_273__40_,r_n_273__39_,r_n_273__38_,r_n_273__37_,r_n_273__36_,
  r_n_273__35_,r_n_273__34_,r_n_273__33_,r_n_273__32_,r_n_273__31_,r_n_273__30_,r_n_273__29_,
  r_n_273__28_,r_n_273__27_,r_n_273__26_,r_n_273__25_,r_n_273__24_,r_n_273__23_,
  r_n_273__22_,r_n_273__21_,r_n_273__20_,r_n_273__19_,r_n_273__18_,r_n_273__17_,
  r_n_273__16_,r_n_273__15_,r_n_273__14_,r_n_273__13_,r_n_273__12_,r_n_273__11_,
  r_n_273__10_,r_n_273__9_,r_n_273__8_,r_n_273__7_,r_n_273__6_,r_n_273__5_,r_n_273__4_,
  r_n_273__3_,r_n_273__2_,r_n_273__1_,r_n_273__0_,r_n_288__63_,r_n_288__62_,
  r_n_288__61_,r_n_288__60_,r_n_288__59_,r_n_288__58_,r_n_288__57_,r_n_288__56_,
  r_n_288__55_,r_n_288__54_,r_n_288__53_,r_n_288__52_,r_n_288__51_,r_n_288__50_,
  r_n_288__49_,r_n_288__48_,r_n_288__47_,r_n_288__46_,r_n_288__45_,r_n_288__44_,r_n_288__43_,
  r_n_288__42_,r_n_288__41_,r_n_288__40_,r_n_288__39_,r_n_288__38_,r_n_288__37_,
  r_n_288__36_,r_n_288__35_,r_n_288__34_,r_n_288__33_,r_n_288__32_,r_n_288__31_,
  r_n_288__30_,r_n_288__29_,r_n_288__28_,r_n_288__27_,r_n_288__26_,r_n_288__25_,
  r_n_288__24_,r_n_288__23_,r_n_288__22_,r_n_288__21_,r_n_288__20_,r_n_288__19_,
  r_n_288__18_,r_n_288__17_,r_n_288__16_,r_n_288__15_,r_n_288__14_,r_n_288__13_,
  r_n_288__12_,r_n_288__11_,r_n_288__10_,r_n_288__9_,r_n_288__8_,r_n_288__7_,r_n_288__6_,
  r_n_288__5_,r_n_288__4_,r_n_288__3_,r_n_288__2_,r_n_288__1_,r_n_288__0_,
  r_n_287__63_,r_n_287__62_,r_n_287__61_,r_n_287__60_,r_n_287__59_,r_n_287__58_,r_n_287__57_,
  r_n_287__56_,r_n_287__55_,r_n_287__54_,r_n_287__53_,r_n_287__52_,r_n_287__51_,
  r_n_287__50_,r_n_287__49_,r_n_287__48_,r_n_287__47_,r_n_287__46_,r_n_287__45_,
  r_n_287__44_,r_n_287__43_,r_n_287__42_,r_n_287__41_,r_n_287__40_,r_n_287__39_,
  r_n_287__38_,r_n_287__37_,r_n_287__36_,r_n_287__35_,r_n_287__34_,r_n_287__33_,
  r_n_287__32_,r_n_287__31_,r_n_287__30_,r_n_287__29_,r_n_287__28_,r_n_287__27_,
  r_n_287__26_,r_n_287__25_,r_n_287__24_,r_n_287__23_,r_n_287__22_,r_n_287__21_,r_n_287__20_,
  r_n_287__19_,r_n_287__18_,r_n_287__17_,r_n_287__16_,r_n_287__15_,r_n_287__14_,
  r_n_287__13_,r_n_287__12_,r_n_287__11_,r_n_287__10_,r_n_287__9_,r_n_287__8_,
  r_n_287__7_,r_n_287__6_,r_n_287__5_,r_n_287__4_,r_n_287__3_,r_n_287__2_,r_n_287__1_,
  r_n_287__0_,r_n_286__63_,r_n_286__62_,r_n_286__61_,r_n_286__60_,r_n_286__59_,
  r_n_286__58_,r_n_286__57_,r_n_286__56_,r_n_286__55_,r_n_286__54_,r_n_286__53_,
  r_n_286__52_,r_n_286__51_,r_n_286__50_,r_n_286__49_,r_n_286__48_,r_n_286__47_,
  r_n_286__46_,r_n_286__45_,r_n_286__44_,r_n_286__43_,r_n_286__42_,r_n_286__41_,
  r_n_286__40_,r_n_286__39_,r_n_286__38_,r_n_286__37_,r_n_286__36_,r_n_286__35_,r_n_286__34_,
  r_n_286__33_,r_n_286__32_,r_n_286__31_,r_n_286__30_,r_n_286__29_,r_n_286__28_,
  r_n_286__27_,r_n_286__26_,r_n_286__25_,r_n_286__24_,r_n_286__23_,r_n_286__22_,
  r_n_286__21_,r_n_286__20_,r_n_286__19_,r_n_286__18_,r_n_286__17_,r_n_286__16_,
  r_n_286__15_,r_n_286__14_,r_n_286__13_,r_n_286__12_,r_n_286__11_,r_n_286__10_,
  r_n_286__9_,r_n_286__8_,r_n_286__7_,r_n_286__6_,r_n_286__5_,r_n_286__4_,r_n_286__3_,
  r_n_286__2_,r_n_286__1_,r_n_286__0_,r_n_285__63_,r_n_285__62_,r_n_285__61_,
  r_n_285__60_,r_n_285__59_,r_n_285__58_,r_n_285__57_,r_n_285__56_,r_n_285__55_,
  r_n_285__54_,r_n_285__53_,r_n_285__52_,r_n_285__51_,r_n_285__50_,r_n_285__49_,r_n_285__48_,
  r_n_285__47_,r_n_285__46_,r_n_285__45_,r_n_285__44_,r_n_285__43_,r_n_285__42_,
  r_n_285__41_,r_n_285__40_,r_n_285__39_,r_n_285__38_,r_n_285__37_,r_n_285__36_,
  r_n_285__35_,r_n_285__34_,r_n_285__33_,r_n_285__32_,r_n_285__31_,r_n_285__30_,
  r_n_285__29_,r_n_285__28_,r_n_285__27_,r_n_285__26_,r_n_285__25_,r_n_285__24_,
  r_n_285__23_,r_n_285__22_,r_n_285__21_,r_n_285__20_,r_n_285__19_,r_n_285__18_,
  r_n_285__17_,r_n_285__16_,r_n_285__15_,r_n_285__14_,r_n_285__13_,r_n_285__12_,
  r_n_285__11_,r_n_285__10_,r_n_285__9_,r_n_285__8_,r_n_285__7_,r_n_285__6_,r_n_285__5_,
  r_n_285__4_,r_n_285__3_,r_n_285__2_,r_n_285__1_,r_n_285__0_,r_n_284__63_,r_n_284__62_,
  r_n_284__61_,r_n_284__60_,r_n_284__59_,r_n_284__58_,r_n_284__57_,r_n_284__56_,
  r_n_284__55_,r_n_284__54_,r_n_284__53_,r_n_284__52_,r_n_284__51_,r_n_284__50_,
  r_n_284__49_,r_n_284__48_,r_n_284__47_,r_n_284__46_,r_n_284__45_,r_n_284__44_,
  r_n_284__43_,r_n_284__42_,r_n_284__41_,r_n_284__40_,r_n_284__39_,r_n_284__38_,
  r_n_284__37_,r_n_284__36_,r_n_284__35_,r_n_284__34_,r_n_284__33_,r_n_284__32_,
  r_n_284__31_,r_n_284__30_,r_n_284__29_,r_n_284__28_,r_n_284__27_,r_n_284__26_,
  r_n_284__25_,r_n_284__24_,r_n_284__23_,r_n_284__22_,r_n_284__21_,r_n_284__20_,r_n_284__19_,
  r_n_284__18_,r_n_284__17_,r_n_284__16_,r_n_284__15_,r_n_284__14_,r_n_284__13_,
  r_n_284__12_,r_n_284__11_,r_n_284__10_,r_n_284__9_,r_n_284__8_,r_n_284__7_,
  r_n_284__6_,r_n_284__5_,r_n_284__4_,r_n_284__3_,r_n_284__2_,r_n_284__1_,r_n_284__0_,
  r_n_283__63_,r_n_283__62_,r_n_283__61_,r_n_283__60_,r_n_283__59_,r_n_283__58_,
  r_n_283__57_,r_n_283__56_,r_n_283__55_,r_n_283__54_,r_n_283__53_,r_n_283__52_,
  r_n_283__51_,r_n_283__50_,r_n_283__49_,r_n_283__48_,r_n_283__47_,r_n_283__46_,
  r_n_283__45_,r_n_283__44_,r_n_283__43_,r_n_283__42_,r_n_283__41_,r_n_283__40_,
  r_n_283__39_,r_n_283__38_,r_n_283__37_,r_n_283__36_,r_n_283__35_,r_n_283__34_,r_n_283__33_,
  r_n_283__32_,r_n_283__31_,r_n_283__30_,r_n_283__29_,r_n_283__28_,r_n_283__27_,
  r_n_283__26_,r_n_283__25_,r_n_283__24_,r_n_283__23_,r_n_283__22_,r_n_283__21_,
  r_n_283__20_,r_n_283__19_,r_n_283__18_,r_n_283__17_,r_n_283__16_,r_n_283__15_,
  r_n_283__14_,r_n_283__13_,r_n_283__12_,r_n_283__11_,r_n_283__10_,r_n_283__9_,
  r_n_283__8_,r_n_283__7_,r_n_283__6_,r_n_283__5_,r_n_283__4_,r_n_283__3_,r_n_283__2_,
  r_n_283__1_,r_n_283__0_,r_n_282__63_,r_n_282__62_,r_n_282__61_,r_n_282__60_,
  r_n_282__59_,r_n_282__58_,r_n_282__57_,r_n_282__56_,r_n_282__55_,r_n_282__54_,
  r_n_282__53_,r_n_282__52_,r_n_282__51_,r_n_282__50_,r_n_282__49_,r_n_282__48_,r_n_282__47_,
  r_n_282__46_,r_n_282__45_,r_n_282__44_,r_n_282__43_,r_n_282__42_,r_n_282__41_,
  r_n_282__40_,r_n_282__39_,r_n_282__38_,r_n_282__37_,r_n_282__36_,r_n_282__35_,
  r_n_282__34_,r_n_282__33_,r_n_282__32_,r_n_282__31_,r_n_282__30_,r_n_282__29_,
  r_n_282__28_,r_n_282__27_,r_n_282__26_,r_n_282__25_,r_n_282__24_,r_n_282__23_,
  r_n_282__22_,r_n_282__21_,r_n_282__20_,r_n_282__19_,r_n_282__18_,r_n_282__17_,
  r_n_282__16_,r_n_282__15_,r_n_282__14_,r_n_282__13_,r_n_282__12_,r_n_282__11_,r_n_282__10_,
  r_n_282__9_,r_n_282__8_,r_n_282__7_,r_n_282__6_,r_n_282__5_,r_n_282__4_,
  r_n_282__3_,r_n_282__2_,r_n_282__1_,r_n_282__0_,r_n_281__63_,r_n_281__62_,r_n_281__61_,
  r_n_281__60_,r_n_281__59_,r_n_281__58_,r_n_281__57_,r_n_281__56_,r_n_281__55_,
  r_n_281__54_,r_n_281__53_,r_n_281__52_,r_n_281__51_,r_n_281__50_,r_n_281__49_,
  r_n_281__48_,r_n_281__47_,r_n_281__46_,r_n_281__45_,r_n_281__44_,r_n_281__43_,
  r_n_281__42_,r_n_281__41_,r_n_281__40_,r_n_281__39_,r_n_281__38_,r_n_281__37_,
  r_n_281__36_,r_n_281__35_,r_n_281__34_,r_n_281__33_,r_n_281__32_,r_n_281__31_,
  r_n_281__30_,r_n_281__29_,r_n_281__28_,r_n_281__27_,r_n_281__26_,r_n_281__25_,r_n_281__24_,
  r_n_281__23_,r_n_281__22_,r_n_281__21_,r_n_281__20_,r_n_281__19_,r_n_281__18_,
  r_n_281__17_,r_n_281__16_,r_n_281__15_,r_n_281__14_,r_n_281__13_,r_n_281__12_,
  r_n_281__11_,r_n_281__10_,r_n_281__9_,r_n_281__8_,r_n_281__7_,r_n_281__6_,
  r_n_281__5_,r_n_281__4_,r_n_281__3_,r_n_281__2_,r_n_281__1_,r_n_281__0_,r_n_296__63_,
  r_n_296__62_,r_n_296__61_,r_n_296__60_,r_n_296__59_,r_n_296__58_,r_n_296__57_,
  r_n_296__56_,r_n_296__55_,r_n_296__54_,r_n_296__53_,r_n_296__52_,r_n_296__51_,
  r_n_296__50_,r_n_296__49_,r_n_296__48_,r_n_296__47_,r_n_296__46_,r_n_296__45_,
  r_n_296__44_,r_n_296__43_,r_n_296__42_,r_n_296__41_,r_n_296__40_,r_n_296__39_,r_n_296__38_,
  r_n_296__37_,r_n_296__36_,r_n_296__35_,r_n_296__34_,r_n_296__33_,r_n_296__32_,
  r_n_296__31_,r_n_296__30_,r_n_296__29_,r_n_296__28_,r_n_296__27_,r_n_296__26_,
  r_n_296__25_,r_n_296__24_,r_n_296__23_,r_n_296__22_,r_n_296__21_,r_n_296__20_,
  r_n_296__19_,r_n_296__18_,r_n_296__17_,r_n_296__16_,r_n_296__15_,r_n_296__14_,
  r_n_296__13_,r_n_296__12_,r_n_296__11_,r_n_296__10_,r_n_296__9_,r_n_296__8_,r_n_296__7_,
  r_n_296__6_,r_n_296__5_,r_n_296__4_,r_n_296__3_,r_n_296__2_,r_n_296__1_,
  r_n_296__0_,r_n_295__63_,r_n_295__62_,r_n_295__61_,r_n_295__60_,r_n_295__59_,
  r_n_295__58_,r_n_295__57_,r_n_295__56_,r_n_295__55_,r_n_295__54_,r_n_295__53_,r_n_295__52_,
  r_n_295__51_,r_n_295__50_,r_n_295__49_,r_n_295__48_,r_n_295__47_,r_n_295__46_,
  r_n_295__45_,r_n_295__44_,r_n_295__43_,r_n_295__42_,r_n_295__41_,r_n_295__40_,
  r_n_295__39_,r_n_295__38_,r_n_295__37_,r_n_295__36_,r_n_295__35_,r_n_295__34_,
  r_n_295__33_,r_n_295__32_,r_n_295__31_,r_n_295__30_,r_n_295__29_,r_n_295__28_,
  r_n_295__27_,r_n_295__26_,r_n_295__25_,r_n_295__24_,r_n_295__23_,r_n_295__22_,
  r_n_295__21_,r_n_295__20_,r_n_295__19_,r_n_295__18_,r_n_295__17_,r_n_295__16_,
  r_n_295__15_,r_n_295__14_,r_n_295__13_,r_n_295__12_,r_n_295__11_,r_n_295__10_,r_n_295__9_,
  r_n_295__8_,r_n_295__7_,r_n_295__6_,r_n_295__5_,r_n_295__4_,r_n_295__3_,
  r_n_295__2_,r_n_295__1_,r_n_295__0_,r_n_294__63_,r_n_294__62_,r_n_294__61_,r_n_294__60_,
  r_n_294__59_,r_n_294__58_,r_n_294__57_,r_n_294__56_,r_n_294__55_,r_n_294__54_,
  r_n_294__53_,r_n_294__52_,r_n_294__51_,r_n_294__50_,r_n_294__49_,r_n_294__48_,
  r_n_294__47_,r_n_294__46_,r_n_294__45_,r_n_294__44_,r_n_294__43_,r_n_294__42_,
  r_n_294__41_,r_n_294__40_,r_n_294__39_,r_n_294__38_,r_n_294__37_,r_n_294__36_,
  r_n_294__35_,r_n_294__34_,r_n_294__33_,r_n_294__32_,r_n_294__31_,r_n_294__30_,
  r_n_294__29_,r_n_294__28_,r_n_294__27_,r_n_294__26_,r_n_294__25_,r_n_294__24_,r_n_294__23_,
  r_n_294__22_,r_n_294__21_,r_n_294__20_,r_n_294__19_,r_n_294__18_,r_n_294__17_,
  r_n_294__16_,r_n_294__15_,r_n_294__14_,r_n_294__13_,r_n_294__12_,r_n_294__11_,
  r_n_294__10_,r_n_294__9_,r_n_294__8_,r_n_294__7_,r_n_294__6_,r_n_294__5_,r_n_294__4_,
  r_n_294__3_,r_n_294__2_,r_n_294__1_,r_n_294__0_,r_n_293__63_,r_n_293__62_,
  r_n_293__61_,r_n_293__60_,r_n_293__59_,r_n_293__58_,r_n_293__57_,r_n_293__56_,
  r_n_293__55_,r_n_293__54_,r_n_293__53_,r_n_293__52_,r_n_293__51_,r_n_293__50_,
  r_n_293__49_,r_n_293__48_,r_n_293__47_,r_n_293__46_,r_n_293__45_,r_n_293__44_,
  r_n_293__43_,r_n_293__42_,r_n_293__41_,r_n_293__40_,r_n_293__39_,r_n_293__38_,r_n_293__37_,
  r_n_293__36_,r_n_293__35_,r_n_293__34_,r_n_293__33_,r_n_293__32_,r_n_293__31_,
  r_n_293__30_,r_n_293__29_,r_n_293__28_,r_n_293__27_,r_n_293__26_,r_n_293__25_,
  r_n_293__24_,r_n_293__23_,r_n_293__22_,r_n_293__21_,r_n_293__20_,r_n_293__19_,
  r_n_293__18_,r_n_293__17_,r_n_293__16_,r_n_293__15_,r_n_293__14_,r_n_293__13_,
  r_n_293__12_,r_n_293__11_,r_n_293__10_,r_n_293__9_,r_n_293__8_,r_n_293__7_,r_n_293__6_,
  r_n_293__5_,r_n_293__4_,r_n_293__3_,r_n_293__2_,r_n_293__1_,r_n_293__0_,
  r_n_292__63_,r_n_292__62_,r_n_292__61_,r_n_292__60_,r_n_292__59_,r_n_292__58_,
  r_n_292__57_,r_n_292__56_,r_n_292__55_,r_n_292__54_,r_n_292__53_,r_n_292__52_,r_n_292__51_,
  r_n_292__50_,r_n_292__49_,r_n_292__48_,r_n_292__47_,r_n_292__46_,r_n_292__45_,
  r_n_292__44_,r_n_292__43_,r_n_292__42_,r_n_292__41_,r_n_292__40_,r_n_292__39_,
  r_n_292__38_,r_n_292__37_,r_n_292__36_,r_n_292__35_,r_n_292__34_,r_n_292__33_,
  r_n_292__32_,r_n_292__31_,r_n_292__30_,r_n_292__29_,r_n_292__28_,r_n_292__27_,
  r_n_292__26_,r_n_292__25_,r_n_292__24_,r_n_292__23_,r_n_292__22_,r_n_292__21_,
  r_n_292__20_,r_n_292__19_,r_n_292__18_,r_n_292__17_,r_n_292__16_,r_n_292__15_,r_n_292__14_,
  r_n_292__13_,r_n_292__12_,r_n_292__11_,r_n_292__10_,r_n_292__9_,r_n_292__8_,
  r_n_292__7_,r_n_292__6_,r_n_292__5_,r_n_292__4_,r_n_292__3_,r_n_292__2_,r_n_292__1_,
  r_n_292__0_,r_n_291__63_,r_n_291__62_,r_n_291__61_,r_n_291__60_,r_n_291__59_,
  r_n_291__58_,r_n_291__57_,r_n_291__56_,r_n_291__55_,r_n_291__54_,r_n_291__53_,
  r_n_291__52_,r_n_291__51_,r_n_291__50_,r_n_291__49_,r_n_291__48_,r_n_291__47_,
  r_n_291__46_,r_n_291__45_,r_n_291__44_,r_n_291__43_,r_n_291__42_,r_n_291__41_,
  r_n_291__40_,r_n_291__39_,r_n_291__38_,r_n_291__37_,r_n_291__36_,r_n_291__35_,
  r_n_291__34_,r_n_291__33_,r_n_291__32_,r_n_291__31_,r_n_291__30_,r_n_291__29_,r_n_291__28_,
  r_n_291__27_,r_n_291__26_,r_n_291__25_,r_n_291__24_,r_n_291__23_,r_n_291__22_,
  r_n_291__21_,r_n_291__20_,r_n_291__19_,r_n_291__18_,r_n_291__17_,r_n_291__16_,
  r_n_291__15_,r_n_291__14_,r_n_291__13_,r_n_291__12_,r_n_291__11_,r_n_291__10_,
  r_n_291__9_,r_n_291__8_,r_n_291__7_,r_n_291__6_,r_n_291__5_,r_n_291__4_,r_n_291__3_,
  r_n_291__2_,r_n_291__1_,r_n_291__0_,r_n_290__63_,r_n_290__62_,r_n_290__61_,
  r_n_290__60_,r_n_290__59_,r_n_290__58_,r_n_290__57_,r_n_290__56_,r_n_290__55_,
  r_n_290__54_,r_n_290__53_,r_n_290__52_,r_n_290__51_,r_n_290__50_,r_n_290__49_,
  r_n_290__48_,r_n_290__47_,r_n_290__46_,r_n_290__45_,r_n_290__44_,r_n_290__43_,r_n_290__42_,
  r_n_290__41_,r_n_290__40_,r_n_290__39_,r_n_290__38_,r_n_290__37_,r_n_290__36_,
  r_n_290__35_,r_n_290__34_,r_n_290__33_,r_n_290__32_,r_n_290__31_,r_n_290__30_,
  r_n_290__29_,r_n_290__28_,r_n_290__27_,r_n_290__26_,r_n_290__25_,r_n_290__24_,
  r_n_290__23_,r_n_290__22_,r_n_290__21_,r_n_290__20_,r_n_290__19_,r_n_290__18_,
  r_n_290__17_,r_n_290__16_,r_n_290__15_,r_n_290__14_,r_n_290__13_,r_n_290__12_,
  r_n_290__11_,r_n_290__10_,r_n_290__9_,r_n_290__8_,r_n_290__7_,r_n_290__6_,r_n_290__5_,
  r_n_290__4_,r_n_290__3_,r_n_290__2_,r_n_290__1_,r_n_290__0_,r_n_289__63_,
  r_n_289__62_,r_n_289__61_,r_n_289__60_,r_n_289__59_,r_n_289__58_,r_n_289__57_,r_n_289__56_,
  r_n_289__55_,r_n_289__54_,r_n_289__53_,r_n_289__52_,r_n_289__51_,r_n_289__50_,
  r_n_289__49_,r_n_289__48_,r_n_289__47_,r_n_289__46_,r_n_289__45_,r_n_289__44_,
  r_n_289__43_,r_n_289__42_,r_n_289__41_,r_n_289__40_,r_n_289__39_,r_n_289__38_,
  r_n_289__37_,r_n_289__36_,r_n_289__35_,r_n_289__34_,r_n_289__33_,r_n_289__32_,
  r_n_289__31_,r_n_289__30_,r_n_289__29_,r_n_289__28_,r_n_289__27_,r_n_289__26_,
  r_n_289__25_,r_n_289__24_,r_n_289__23_,r_n_289__22_,r_n_289__21_,r_n_289__20_,
  r_n_289__19_,r_n_289__18_,r_n_289__17_,r_n_289__16_,r_n_289__15_,r_n_289__14_,r_n_289__13_,
  r_n_289__12_,r_n_289__11_,r_n_289__10_,r_n_289__9_,r_n_289__8_,r_n_289__7_,
  r_n_289__6_,r_n_289__5_,r_n_289__4_,r_n_289__3_,r_n_289__2_,r_n_289__1_,r_n_289__0_,
  r_n_304__63_,r_n_304__62_,r_n_304__61_,r_n_304__60_,r_n_304__59_,r_n_304__58_,
  r_n_304__57_,r_n_304__56_,r_n_304__55_,r_n_304__54_,r_n_304__53_,r_n_304__52_,
  r_n_304__51_,r_n_304__50_,r_n_304__49_,r_n_304__48_,r_n_304__47_,r_n_304__46_,
  r_n_304__45_,r_n_304__44_,r_n_304__43_,r_n_304__42_,r_n_304__41_,r_n_304__40_,
  r_n_304__39_,r_n_304__38_,r_n_304__37_,r_n_304__36_,r_n_304__35_,r_n_304__34_,
  r_n_304__33_,r_n_304__32_,r_n_304__31_,r_n_304__30_,r_n_304__29_,r_n_304__28_,r_n_304__27_,
  r_n_304__26_,r_n_304__25_,r_n_304__24_,r_n_304__23_,r_n_304__22_,r_n_304__21_,
  r_n_304__20_,r_n_304__19_,r_n_304__18_,r_n_304__17_,r_n_304__16_,r_n_304__15_,
  r_n_304__14_,r_n_304__13_,r_n_304__12_,r_n_304__11_,r_n_304__10_,r_n_304__9_,
  r_n_304__8_,r_n_304__7_,r_n_304__6_,r_n_304__5_,r_n_304__4_,r_n_304__3_,r_n_304__2_,
  r_n_304__1_,r_n_304__0_,r_n_303__63_,r_n_303__62_,r_n_303__61_,r_n_303__60_,
  r_n_303__59_,r_n_303__58_,r_n_303__57_,r_n_303__56_,r_n_303__55_,r_n_303__54_,
  r_n_303__53_,r_n_303__52_,r_n_303__51_,r_n_303__50_,r_n_303__49_,r_n_303__48_,
  r_n_303__47_,r_n_303__46_,r_n_303__45_,r_n_303__44_,r_n_303__43_,r_n_303__42_,r_n_303__41_,
  r_n_303__40_,r_n_303__39_,r_n_303__38_,r_n_303__37_,r_n_303__36_,r_n_303__35_,
  r_n_303__34_,r_n_303__33_,r_n_303__32_,r_n_303__31_,r_n_303__30_,r_n_303__29_,
  r_n_303__28_,r_n_303__27_,r_n_303__26_,r_n_303__25_,r_n_303__24_,r_n_303__23_,
  r_n_303__22_,r_n_303__21_,r_n_303__20_,r_n_303__19_,r_n_303__18_,r_n_303__17_,
  r_n_303__16_,r_n_303__15_,r_n_303__14_,r_n_303__13_,r_n_303__12_,r_n_303__11_,
  r_n_303__10_,r_n_303__9_,r_n_303__8_,r_n_303__7_,r_n_303__6_,r_n_303__5_,r_n_303__4_,
  r_n_303__3_,r_n_303__2_,r_n_303__1_,r_n_303__0_,r_n_302__63_,r_n_302__62_,
  r_n_302__61_,r_n_302__60_,r_n_302__59_,r_n_302__58_,r_n_302__57_,r_n_302__56_,r_n_302__55_,
  r_n_302__54_,r_n_302__53_,r_n_302__52_,r_n_302__51_,r_n_302__50_,r_n_302__49_,
  r_n_302__48_,r_n_302__47_,r_n_302__46_,r_n_302__45_,r_n_302__44_,r_n_302__43_,
  r_n_302__42_,r_n_302__41_,r_n_302__40_,r_n_302__39_,r_n_302__38_,r_n_302__37_,
  r_n_302__36_,r_n_302__35_,r_n_302__34_,r_n_302__33_,r_n_302__32_,r_n_302__31_,
  r_n_302__30_,r_n_302__29_,r_n_302__28_,r_n_302__27_,r_n_302__26_,r_n_302__25_,
  r_n_302__24_,r_n_302__23_,r_n_302__22_,r_n_302__21_,r_n_302__20_,r_n_302__19_,r_n_302__18_,
  r_n_302__17_,r_n_302__16_,r_n_302__15_,r_n_302__14_,r_n_302__13_,r_n_302__12_,
  r_n_302__11_,r_n_302__10_,r_n_302__9_,r_n_302__8_,r_n_302__7_,r_n_302__6_,
  r_n_302__5_,r_n_302__4_,r_n_302__3_,r_n_302__2_,r_n_302__1_,r_n_302__0_,r_n_301__63_,
  r_n_301__62_,r_n_301__61_,r_n_301__60_,r_n_301__59_,r_n_301__58_,r_n_301__57_,
  r_n_301__56_,r_n_301__55_,r_n_301__54_,r_n_301__53_,r_n_301__52_,r_n_301__51_,
  r_n_301__50_,r_n_301__49_,r_n_301__48_,r_n_301__47_,r_n_301__46_,r_n_301__45_,
  r_n_301__44_,r_n_301__43_,r_n_301__42_,r_n_301__41_,r_n_301__40_,r_n_301__39_,
  r_n_301__38_,r_n_301__37_,r_n_301__36_,r_n_301__35_,r_n_301__34_,r_n_301__33_,r_n_301__32_,
  r_n_301__31_,r_n_301__30_,r_n_301__29_,r_n_301__28_,r_n_301__27_,r_n_301__26_,
  r_n_301__25_,r_n_301__24_,r_n_301__23_,r_n_301__22_,r_n_301__21_,r_n_301__20_,
  r_n_301__19_,r_n_301__18_,r_n_301__17_,r_n_301__16_,r_n_301__15_,r_n_301__14_,
  r_n_301__13_,r_n_301__12_,r_n_301__11_,r_n_301__10_,r_n_301__9_,r_n_301__8_,
  r_n_301__7_,r_n_301__6_,r_n_301__5_,r_n_301__4_,r_n_301__3_,r_n_301__2_,r_n_301__1_,
  r_n_301__0_,r_n_300__63_,r_n_300__62_,r_n_300__61_,r_n_300__60_,r_n_300__59_,
  r_n_300__58_,r_n_300__57_,r_n_300__56_,r_n_300__55_,r_n_300__54_,r_n_300__53_,
  r_n_300__52_,r_n_300__51_,r_n_300__50_,r_n_300__49_,r_n_300__48_,r_n_300__47_,r_n_300__46_,
  r_n_300__45_,r_n_300__44_,r_n_300__43_,r_n_300__42_,r_n_300__41_,r_n_300__40_,
  r_n_300__39_,r_n_300__38_,r_n_300__37_,r_n_300__36_,r_n_300__35_,r_n_300__34_,
  r_n_300__33_,r_n_300__32_,r_n_300__31_,r_n_300__30_,r_n_300__29_,r_n_300__28_,
  r_n_300__27_,r_n_300__26_,r_n_300__25_,r_n_300__24_,r_n_300__23_,r_n_300__22_,
  r_n_300__21_,r_n_300__20_,r_n_300__19_,r_n_300__18_,r_n_300__17_,r_n_300__16_,
  r_n_300__15_,r_n_300__14_,r_n_300__13_,r_n_300__12_,r_n_300__11_,r_n_300__10_,r_n_300__9_,
  r_n_300__8_,r_n_300__7_,r_n_300__6_,r_n_300__5_,r_n_300__4_,r_n_300__3_,
  r_n_300__2_,r_n_300__1_,r_n_300__0_,r_n_299__63_,r_n_299__62_,r_n_299__61_,r_n_299__60_,
  r_n_299__59_,r_n_299__58_,r_n_299__57_,r_n_299__56_,r_n_299__55_,r_n_299__54_,
  r_n_299__53_,r_n_299__52_,r_n_299__51_,r_n_299__50_,r_n_299__49_,r_n_299__48_,
  r_n_299__47_,r_n_299__46_,r_n_299__45_,r_n_299__44_,r_n_299__43_,r_n_299__42_,
  r_n_299__41_,r_n_299__40_,r_n_299__39_,r_n_299__38_,r_n_299__37_,r_n_299__36_,
  r_n_299__35_,r_n_299__34_,r_n_299__33_,r_n_299__32_,r_n_299__31_,r_n_299__30_,
  r_n_299__29_,r_n_299__28_,r_n_299__27_,r_n_299__26_,r_n_299__25_,r_n_299__24_,
  r_n_299__23_,r_n_299__22_,r_n_299__21_,r_n_299__20_,r_n_299__19_,r_n_299__18_,r_n_299__17_,
  r_n_299__16_,r_n_299__15_,r_n_299__14_,r_n_299__13_,r_n_299__12_,r_n_299__11_,
  r_n_299__10_,r_n_299__9_,r_n_299__8_,r_n_299__7_,r_n_299__6_,r_n_299__5_,
  r_n_299__4_,r_n_299__3_,r_n_299__2_,r_n_299__1_,r_n_299__0_,r_n_298__63_,r_n_298__62_,
  r_n_298__61_,r_n_298__60_,r_n_298__59_,r_n_298__58_,r_n_298__57_,r_n_298__56_,
  r_n_298__55_,r_n_298__54_,r_n_298__53_,r_n_298__52_,r_n_298__51_,r_n_298__50_,
  r_n_298__49_,r_n_298__48_,r_n_298__47_,r_n_298__46_,r_n_298__45_,r_n_298__44_,
  r_n_298__43_,r_n_298__42_,r_n_298__41_,r_n_298__40_,r_n_298__39_,r_n_298__38_,
  r_n_298__37_,r_n_298__36_,r_n_298__35_,r_n_298__34_,r_n_298__33_,r_n_298__32_,r_n_298__31_,
  r_n_298__30_,r_n_298__29_,r_n_298__28_,r_n_298__27_,r_n_298__26_,r_n_298__25_,
  r_n_298__24_,r_n_298__23_,r_n_298__22_,r_n_298__21_,r_n_298__20_,r_n_298__19_,
  r_n_298__18_,r_n_298__17_,r_n_298__16_,r_n_298__15_,r_n_298__14_,r_n_298__13_,
  r_n_298__12_,r_n_298__11_,r_n_298__10_,r_n_298__9_,r_n_298__8_,r_n_298__7_,r_n_298__6_,
  r_n_298__5_,r_n_298__4_,r_n_298__3_,r_n_298__2_,r_n_298__1_,r_n_298__0_,
  r_n_297__63_,r_n_297__62_,r_n_297__61_,r_n_297__60_,r_n_297__59_,r_n_297__58_,
  r_n_297__57_,r_n_297__56_,r_n_297__55_,r_n_297__54_,r_n_297__53_,r_n_297__52_,
  r_n_297__51_,r_n_297__50_,r_n_297__49_,r_n_297__48_,r_n_297__47_,r_n_297__46_,r_n_297__45_,
  r_n_297__44_,r_n_297__43_,r_n_297__42_,r_n_297__41_,r_n_297__40_,r_n_297__39_,
  r_n_297__38_,r_n_297__37_,r_n_297__36_,r_n_297__35_,r_n_297__34_,r_n_297__33_,
  r_n_297__32_,r_n_297__31_,r_n_297__30_,r_n_297__29_,r_n_297__28_,r_n_297__27_,
  r_n_297__26_,r_n_297__25_,r_n_297__24_,r_n_297__23_,r_n_297__22_,r_n_297__21_,
  r_n_297__20_,r_n_297__19_,r_n_297__18_,r_n_297__17_,r_n_297__16_,r_n_297__15_,
  r_n_297__14_,r_n_297__13_,r_n_297__12_,r_n_297__11_,r_n_297__10_,r_n_297__9_,r_n_297__8_,
  r_n_297__7_,r_n_297__6_,r_n_297__5_,r_n_297__4_,r_n_297__3_,r_n_297__2_,
  r_n_297__1_,r_n_297__0_,r_n_312__63_,r_n_312__62_,r_n_312__61_,r_n_312__60_,r_n_312__59_,
  r_n_312__58_,r_n_312__57_,r_n_312__56_,r_n_312__55_,r_n_312__54_,r_n_312__53_,
  r_n_312__52_,r_n_312__51_,r_n_312__50_,r_n_312__49_,r_n_312__48_,r_n_312__47_,
  r_n_312__46_,r_n_312__45_,r_n_312__44_,r_n_312__43_,r_n_312__42_,r_n_312__41_,
  r_n_312__40_,r_n_312__39_,r_n_312__38_,r_n_312__37_,r_n_312__36_,r_n_312__35_,
  r_n_312__34_,r_n_312__33_,r_n_312__32_,r_n_312__31_,r_n_312__30_,r_n_312__29_,
  r_n_312__28_,r_n_312__27_,r_n_312__26_,r_n_312__25_,r_n_312__24_,r_n_312__23_,r_n_312__22_,
  r_n_312__21_,r_n_312__20_,r_n_312__19_,r_n_312__18_,r_n_312__17_,r_n_312__16_,
  r_n_312__15_,r_n_312__14_,r_n_312__13_,r_n_312__12_,r_n_312__11_,r_n_312__10_,
  r_n_312__9_,r_n_312__8_,r_n_312__7_,r_n_312__6_,r_n_312__5_,r_n_312__4_,r_n_312__3_,
  r_n_312__2_,r_n_312__1_,r_n_312__0_,r_n_311__63_,r_n_311__62_,r_n_311__61_,
  r_n_311__60_,r_n_311__59_,r_n_311__58_,r_n_311__57_,r_n_311__56_,r_n_311__55_,
  r_n_311__54_,r_n_311__53_,r_n_311__52_,r_n_311__51_,r_n_311__50_,r_n_311__49_,
  r_n_311__48_,r_n_311__47_,r_n_311__46_,r_n_311__45_,r_n_311__44_,r_n_311__43_,
  r_n_311__42_,r_n_311__41_,r_n_311__40_,r_n_311__39_,r_n_311__38_,r_n_311__37_,r_n_311__36_,
  r_n_311__35_,r_n_311__34_,r_n_311__33_,r_n_311__32_,r_n_311__31_,r_n_311__30_,
  r_n_311__29_,r_n_311__28_,r_n_311__27_,r_n_311__26_,r_n_311__25_,r_n_311__24_,
  r_n_311__23_,r_n_311__22_,r_n_311__21_,r_n_311__20_,r_n_311__19_,r_n_311__18_,
  r_n_311__17_,r_n_311__16_,r_n_311__15_,r_n_311__14_,r_n_311__13_,r_n_311__12_,
  r_n_311__11_,r_n_311__10_,r_n_311__9_,r_n_311__8_,r_n_311__7_,r_n_311__6_,r_n_311__5_,
  r_n_311__4_,r_n_311__3_,r_n_311__2_,r_n_311__1_,r_n_311__0_,r_n_310__63_,
  r_n_310__62_,r_n_310__61_,r_n_310__60_,r_n_310__59_,r_n_310__58_,r_n_310__57_,
  r_n_310__56_,r_n_310__55_,r_n_310__54_,r_n_310__53_,r_n_310__52_,r_n_310__51_,r_n_310__50_,
  r_n_310__49_,r_n_310__48_,r_n_310__47_,r_n_310__46_,r_n_310__45_,r_n_310__44_,
  r_n_310__43_,r_n_310__42_,r_n_310__41_,r_n_310__40_,r_n_310__39_,r_n_310__38_,
  r_n_310__37_,r_n_310__36_,r_n_310__35_,r_n_310__34_,r_n_310__33_,r_n_310__32_,
  r_n_310__31_,r_n_310__30_,r_n_310__29_,r_n_310__28_,r_n_310__27_,r_n_310__26_,
  r_n_310__25_,r_n_310__24_,r_n_310__23_,r_n_310__22_,r_n_310__21_,r_n_310__20_,
  r_n_310__19_,r_n_310__18_,r_n_310__17_,r_n_310__16_,r_n_310__15_,r_n_310__14_,
  r_n_310__13_,r_n_310__12_,r_n_310__11_,r_n_310__10_,r_n_310__9_,r_n_310__8_,r_n_310__7_,
  r_n_310__6_,r_n_310__5_,r_n_310__4_,r_n_310__3_,r_n_310__2_,r_n_310__1_,r_n_310__0_,
  r_n_309__63_,r_n_309__62_,r_n_309__61_,r_n_309__60_,r_n_309__59_,r_n_309__58_,
  r_n_309__57_,r_n_309__56_,r_n_309__55_,r_n_309__54_,r_n_309__53_,r_n_309__52_,
  r_n_309__51_,r_n_309__50_,r_n_309__49_,r_n_309__48_,r_n_309__47_,r_n_309__46_,
  r_n_309__45_,r_n_309__44_,r_n_309__43_,r_n_309__42_,r_n_309__41_,r_n_309__40_,
  r_n_309__39_,r_n_309__38_,r_n_309__37_,r_n_309__36_,r_n_309__35_,r_n_309__34_,
  r_n_309__33_,r_n_309__32_,r_n_309__31_,r_n_309__30_,r_n_309__29_,r_n_309__28_,
  r_n_309__27_,r_n_309__26_,r_n_309__25_,r_n_309__24_,r_n_309__23_,r_n_309__22_,r_n_309__21_,
  r_n_309__20_,r_n_309__19_,r_n_309__18_,r_n_309__17_,r_n_309__16_,r_n_309__15_,
  r_n_309__14_,r_n_309__13_,r_n_309__12_,r_n_309__11_,r_n_309__10_,r_n_309__9_,
  r_n_309__8_,r_n_309__7_,r_n_309__6_,r_n_309__5_,r_n_309__4_,r_n_309__3_,r_n_309__2_,
  r_n_309__1_,r_n_309__0_,r_n_308__63_,r_n_308__62_,r_n_308__61_,r_n_308__60_,
  r_n_308__59_,r_n_308__58_,r_n_308__57_,r_n_308__56_,r_n_308__55_,r_n_308__54_,
  r_n_308__53_,r_n_308__52_,r_n_308__51_,r_n_308__50_,r_n_308__49_,r_n_308__48_,
  r_n_308__47_,r_n_308__46_,r_n_308__45_,r_n_308__44_,r_n_308__43_,r_n_308__42_,
  r_n_308__41_,r_n_308__40_,r_n_308__39_,r_n_308__38_,r_n_308__37_,r_n_308__36_,r_n_308__35_,
  r_n_308__34_,r_n_308__33_,r_n_308__32_,r_n_308__31_,r_n_308__30_,r_n_308__29_,
  r_n_308__28_,r_n_308__27_,r_n_308__26_,r_n_308__25_,r_n_308__24_,r_n_308__23_,
  r_n_308__22_,r_n_308__21_,r_n_308__20_,r_n_308__19_,r_n_308__18_,r_n_308__17_,
  r_n_308__16_,r_n_308__15_,r_n_308__14_,r_n_308__13_,r_n_308__12_,r_n_308__11_,
  r_n_308__10_,r_n_308__9_,r_n_308__8_,r_n_308__7_,r_n_308__6_,r_n_308__5_,r_n_308__4_,
  r_n_308__3_,r_n_308__2_,r_n_308__1_,r_n_308__0_,r_n_307__63_,r_n_307__62_,
  r_n_307__61_,r_n_307__60_,r_n_307__59_,r_n_307__58_,r_n_307__57_,r_n_307__56_,
  r_n_307__55_,r_n_307__54_,r_n_307__53_,r_n_307__52_,r_n_307__51_,r_n_307__50_,r_n_307__49_,
  r_n_307__48_,r_n_307__47_,r_n_307__46_,r_n_307__45_,r_n_307__44_,r_n_307__43_,
  r_n_307__42_,r_n_307__41_,r_n_307__40_,r_n_307__39_,r_n_307__38_,r_n_307__37_,
  r_n_307__36_,r_n_307__35_,r_n_307__34_,r_n_307__33_,r_n_307__32_,r_n_307__31_,
  r_n_307__30_,r_n_307__29_,r_n_307__28_,r_n_307__27_,r_n_307__26_,r_n_307__25_,
  r_n_307__24_,r_n_307__23_,r_n_307__22_,r_n_307__21_,r_n_307__20_,r_n_307__19_,
  r_n_307__18_,r_n_307__17_,r_n_307__16_,r_n_307__15_,r_n_307__14_,r_n_307__13_,r_n_307__12_,
  r_n_307__11_,r_n_307__10_,r_n_307__9_,r_n_307__8_,r_n_307__7_,r_n_307__6_,
  r_n_307__5_,r_n_307__4_,r_n_307__3_,r_n_307__2_,r_n_307__1_,r_n_307__0_,r_n_306__63_,
  r_n_306__62_,r_n_306__61_,r_n_306__60_,r_n_306__59_,r_n_306__58_,r_n_306__57_,
  r_n_306__56_,r_n_306__55_,r_n_306__54_,r_n_306__53_,r_n_306__52_,r_n_306__51_,
  r_n_306__50_,r_n_306__49_,r_n_306__48_,r_n_306__47_,r_n_306__46_,r_n_306__45_,
  r_n_306__44_,r_n_306__43_,r_n_306__42_,r_n_306__41_,r_n_306__40_,r_n_306__39_,
  r_n_306__38_,r_n_306__37_,r_n_306__36_,r_n_306__35_,r_n_306__34_,r_n_306__33_,
  r_n_306__32_,r_n_306__31_,r_n_306__30_,r_n_306__29_,r_n_306__28_,r_n_306__27_,r_n_306__26_,
  r_n_306__25_,r_n_306__24_,r_n_306__23_,r_n_306__22_,r_n_306__21_,r_n_306__20_,
  r_n_306__19_,r_n_306__18_,r_n_306__17_,r_n_306__16_,r_n_306__15_,r_n_306__14_,
  r_n_306__13_,r_n_306__12_,r_n_306__11_,r_n_306__10_,r_n_306__9_,r_n_306__8_,
  r_n_306__7_,r_n_306__6_,r_n_306__5_,r_n_306__4_,r_n_306__3_,r_n_306__2_,r_n_306__1_,
  r_n_306__0_,r_n_305__63_,r_n_305__62_,r_n_305__61_,r_n_305__60_,r_n_305__59_,
  r_n_305__58_,r_n_305__57_,r_n_305__56_,r_n_305__55_,r_n_305__54_,r_n_305__53_,
  r_n_305__52_,r_n_305__51_,r_n_305__50_,r_n_305__49_,r_n_305__48_,r_n_305__47_,
  r_n_305__46_,r_n_305__45_,r_n_305__44_,r_n_305__43_,r_n_305__42_,r_n_305__41_,r_n_305__40_,
  r_n_305__39_,r_n_305__38_,r_n_305__37_,r_n_305__36_,r_n_305__35_,r_n_305__34_,
  r_n_305__33_,r_n_305__32_,r_n_305__31_,r_n_305__30_,r_n_305__29_,r_n_305__28_,
  r_n_305__27_,r_n_305__26_,r_n_305__25_,r_n_305__24_,r_n_305__23_,r_n_305__22_,
  r_n_305__21_,r_n_305__20_,r_n_305__19_,r_n_305__18_,r_n_305__17_,r_n_305__16_,
  r_n_305__15_,r_n_305__14_,r_n_305__13_,r_n_305__12_,r_n_305__11_,r_n_305__10_,
  r_n_305__9_,r_n_305__8_,r_n_305__7_,r_n_305__6_,r_n_305__5_,r_n_305__4_,r_n_305__3_,
  r_n_305__2_,r_n_305__1_,r_n_305__0_,r_n_320__63_,r_n_320__62_,r_n_320__61_,
  r_n_320__60_,r_n_320__59_,r_n_320__58_,r_n_320__57_,r_n_320__56_,r_n_320__55_,r_n_320__54_,
  r_n_320__53_,r_n_320__52_,r_n_320__51_,r_n_320__50_,r_n_320__49_,r_n_320__48_,
  r_n_320__47_,r_n_320__46_,r_n_320__45_,r_n_320__44_,r_n_320__43_,r_n_320__42_,
  r_n_320__41_,r_n_320__40_,r_n_320__39_,r_n_320__38_,r_n_320__37_,r_n_320__36_,
  r_n_320__35_,r_n_320__34_,r_n_320__33_,r_n_320__32_,r_n_320__31_,r_n_320__30_,
  r_n_320__29_,r_n_320__28_,r_n_320__27_,r_n_320__26_,r_n_320__25_,r_n_320__24_,
  r_n_320__23_,r_n_320__22_,r_n_320__21_,r_n_320__20_,r_n_320__19_,r_n_320__18_,
  r_n_320__17_,r_n_320__16_,r_n_320__15_,r_n_320__14_,r_n_320__13_,r_n_320__12_,r_n_320__11_,
  r_n_320__10_,r_n_320__9_,r_n_320__8_,r_n_320__7_,r_n_320__6_,r_n_320__5_,
  r_n_320__4_,r_n_320__3_,r_n_320__2_,r_n_320__1_,r_n_320__0_,r_n_319__63_,r_n_319__62_,
  r_n_319__61_,r_n_319__60_,r_n_319__59_,r_n_319__58_,r_n_319__57_,r_n_319__56_,
  r_n_319__55_,r_n_319__54_,r_n_319__53_,r_n_319__52_,r_n_319__51_,r_n_319__50_,
  r_n_319__49_,r_n_319__48_,r_n_319__47_,r_n_319__46_,r_n_319__45_,r_n_319__44_,
  r_n_319__43_,r_n_319__42_,r_n_319__41_,r_n_319__40_,r_n_319__39_,r_n_319__38_,
  r_n_319__37_,r_n_319__36_,r_n_319__35_,r_n_319__34_,r_n_319__33_,r_n_319__32_,
  r_n_319__31_,r_n_319__30_,r_n_319__29_,r_n_319__28_,r_n_319__27_,r_n_319__26_,r_n_319__25_,
  r_n_319__24_,r_n_319__23_,r_n_319__22_,r_n_319__21_,r_n_319__20_,r_n_319__19_,
  r_n_319__18_,r_n_319__17_,r_n_319__16_,r_n_319__15_,r_n_319__14_,r_n_319__13_,
  r_n_319__12_,r_n_319__11_,r_n_319__10_,r_n_319__9_,r_n_319__8_,r_n_319__7_,
  r_n_319__6_,r_n_319__5_,r_n_319__4_,r_n_319__3_,r_n_319__2_,r_n_319__1_,r_n_319__0_,
  r_n_318__63_,r_n_318__62_,r_n_318__61_,r_n_318__60_,r_n_318__59_,r_n_318__58_,
  r_n_318__57_,r_n_318__56_,r_n_318__55_,r_n_318__54_,r_n_318__53_,r_n_318__52_,
  r_n_318__51_,r_n_318__50_,r_n_318__49_,r_n_318__48_,r_n_318__47_,r_n_318__46_,
  r_n_318__45_,r_n_318__44_,r_n_318__43_,r_n_318__42_,r_n_318__41_,r_n_318__40_,r_n_318__39_,
  r_n_318__38_,r_n_318__37_,r_n_318__36_,r_n_318__35_,r_n_318__34_,r_n_318__33_,
  r_n_318__32_,r_n_318__31_,r_n_318__30_,r_n_318__29_,r_n_318__28_,r_n_318__27_,
  r_n_318__26_,r_n_318__25_,r_n_318__24_,r_n_318__23_,r_n_318__22_,r_n_318__21_,
  r_n_318__20_,r_n_318__19_,r_n_318__18_,r_n_318__17_,r_n_318__16_,r_n_318__15_,
  r_n_318__14_,r_n_318__13_,r_n_318__12_,r_n_318__11_,r_n_318__10_,r_n_318__9_,r_n_318__8_,
  r_n_318__7_,r_n_318__6_,r_n_318__5_,r_n_318__4_,r_n_318__3_,r_n_318__2_,
  r_n_318__1_,r_n_318__0_,r_n_317__63_,r_n_317__62_,r_n_317__61_,r_n_317__60_,
  r_n_317__59_,r_n_317__58_,r_n_317__57_,r_n_317__56_,r_n_317__55_,r_n_317__54_,r_n_317__53_,
  r_n_317__52_,r_n_317__51_,r_n_317__50_,r_n_317__49_,r_n_317__48_,r_n_317__47_,
  r_n_317__46_,r_n_317__45_,r_n_317__44_,r_n_317__43_,r_n_317__42_,r_n_317__41_,
  r_n_317__40_,r_n_317__39_,r_n_317__38_,r_n_317__37_,r_n_317__36_,r_n_317__35_,
  r_n_317__34_,r_n_317__33_,r_n_317__32_,r_n_317__31_,r_n_317__30_,r_n_317__29_,
  r_n_317__28_,r_n_317__27_,r_n_317__26_,r_n_317__25_,r_n_317__24_,r_n_317__23_,
  r_n_317__22_,r_n_317__21_,r_n_317__20_,r_n_317__19_,r_n_317__18_,r_n_317__17_,r_n_317__16_,
  r_n_317__15_,r_n_317__14_,r_n_317__13_,r_n_317__12_,r_n_317__11_,r_n_317__10_,
  r_n_317__9_,r_n_317__8_,r_n_317__7_,r_n_317__6_,r_n_317__5_,r_n_317__4_,
  r_n_317__3_,r_n_317__2_,r_n_317__1_,r_n_317__0_,r_n_316__63_,r_n_316__62_,r_n_316__61_,
  r_n_316__60_,r_n_316__59_,r_n_316__58_,r_n_316__57_,r_n_316__56_,r_n_316__55_,
  r_n_316__54_,r_n_316__53_,r_n_316__52_,r_n_316__51_,r_n_316__50_,r_n_316__49_,
  r_n_316__48_,r_n_316__47_,r_n_316__46_,r_n_316__45_,r_n_316__44_,r_n_316__43_,
  r_n_316__42_,r_n_316__41_,r_n_316__40_,r_n_316__39_,r_n_316__38_,r_n_316__37_,
  r_n_316__36_,r_n_316__35_,r_n_316__34_,r_n_316__33_,r_n_316__32_,r_n_316__31_,r_n_316__30_,
  r_n_316__29_,r_n_316__28_,r_n_316__27_,r_n_316__26_,r_n_316__25_,r_n_316__24_,
  r_n_316__23_,r_n_316__22_,r_n_316__21_,r_n_316__20_,r_n_316__19_,r_n_316__18_,
  r_n_316__17_,r_n_316__16_,r_n_316__15_,r_n_316__14_,r_n_316__13_,r_n_316__12_,
  r_n_316__11_,r_n_316__10_,r_n_316__9_,r_n_316__8_,r_n_316__7_,r_n_316__6_,r_n_316__5_,
  r_n_316__4_,r_n_316__3_,r_n_316__2_,r_n_316__1_,r_n_316__0_,r_n_315__63_,
  r_n_315__62_,r_n_315__61_,r_n_315__60_,r_n_315__59_,r_n_315__58_,r_n_315__57_,
  r_n_315__56_,r_n_315__55_,r_n_315__54_,r_n_315__53_,r_n_315__52_,r_n_315__51_,
  r_n_315__50_,r_n_315__49_,r_n_315__48_,r_n_315__47_,r_n_315__46_,r_n_315__45_,r_n_315__44_,
  r_n_315__43_,r_n_315__42_,r_n_315__41_,r_n_315__40_,r_n_315__39_,r_n_315__38_,
  r_n_315__37_,r_n_315__36_,r_n_315__35_,r_n_315__34_,r_n_315__33_,r_n_315__32_,
  r_n_315__31_,r_n_315__30_,r_n_315__29_,r_n_315__28_,r_n_315__27_,r_n_315__26_,
  r_n_315__25_,r_n_315__24_,r_n_315__23_,r_n_315__22_,r_n_315__21_,r_n_315__20_,
  r_n_315__19_,r_n_315__18_,r_n_315__17_,r_n_315__16_,r_n_315__15_,r_n_315__14_,
  r_n_315__13_,r_n_315__12_,r_n_315__11_,r_n_315__10_,r_n_315__9_,r_n_315__8_,r_n_315__7_,
  r_n_315__6_,r_n_315__5_,r_n_315__4_,r_n_315__3_,r_n_315__2_,r_n_315__1_,
  r_n_315__0_,r_n_314__63_,r_n_314__62_,r_n_314__61_,r_n_314__60_,r_n_314__59_,r_n_314__58_,
  r_n_314__57_,r_n_314__56_,r_n_314__55_,r_n_314__54_,r_n_314__53_,r_n_314__52_,
  r_n_314__51_,r_n_314__50_,r_n_314__49_,r_n_314__48_,r_n_314__47_,r_n_314__46_,
  r_n_314__45_,r_n_314__44_,r_n_314__43_,r_n_314__42_,r_n_314__41_,r_n_314__40_,
  r_n_314__39_,r_n_314__38_,r_n_314__37_,r_n_314__36_,r_n_314__35_,r_n_314__34_,
  r_n_314__33_,r_n_314__32_,r_n_314__31_,r_n_314__30_,r_n_314__29_,r_n_314__28_,
  r_n_314__27_,r_n_314__26_,r_n_314__25_,r_n_314__24_,r_n_314__23_,r_n_314__22_,
  r_n_314__21_,r_n_314__20_,r_n_314__19_,r_n_314__18_,r_n_314__17_,r_n_314__16_,r_n_314__15_,
  r_n_314__14_,r_n_314__13_,r_n_314__12_,r_n_314__11_,r_n_314__10_,r_n_314__9_,
  r_n_314__8_,r_n_314__7_,r_n_314__6_,r_n_314__5_,r_n_314__4_,r_n_314__3_,r_n_314__2_,
  r_n_314__1_,r_n_314__0_,r_n_313__63_,r_n_313__62_,r_n_313__61_,r_n_313__60_,
  r_n_313__59_,r_n_313__58_,r_n_313__57_,r_n_313__56_,r_n_313__55_,r_n_313__54_,
  r_n_313__53_,r_n_313__52_,r_n_313__51_,r_n_313__50_,r_n_313__49_,r_n_313__48_,
  r_n_313__47_,r_n_313__46_,r_n_313__45_,r_n_313__44_,r_n_313__43_,r_n_313__42_,
  r_n_313__41_,r_n_313__40_,r_n_313__39_,r_n_313__38_,r_n_313__37_,r_n_313__36_,
  r_n_313__35_,r_n_313__34_,r_n_313__33_,r_n_313__32_,r_n_313__31_,r_n_313__30_,r_n_313__29_,
  r_n_313__28_,r_n_313__27_,r_n_313__26_,r_n_313__25_,r_n_313__24_,r_n_313__23_,
  r_n_313__22_,r_n_313__21_,r_n_313__20_,r_n_313__19_,r_n_313__18_,r_n_313__17_,
  r_n_313__16_,r_n_313__15_,r_n_313__14_,r_n_313__13_,r_n_313__12_,r_n_313__11_,
  r_n_313__10_,r_n_313__9_,r_n_313__8_,r_n_313__7_,r_n_313__6_,r_n_313__5_,r_n_313__4_,
  r_n_313__3_,r_n_313__2_,r_n_313__1_,r_n_313__0_,r_n_328__63_,r_n_328__62_,
  r_n_328__61_,r_n_328__60_,r_n_328__59_,r_n_328__58_,r_n_328__57_,r_n_328__56_,
  r_n_328__55_,r_n_328__54_,r_n_328__53_,r_n_328__52_,r_n_328__51_,r_n_328__50_,
  r_n_328__49_,r_n_328__48_,r_n_328__47_,r_n_328__46_,r_n_328__45_,r_n_328__44_,r_n_328__43_,
  r_n_328__42_,r_n_328__41_,r_n_328__40_,r_n_328__39_,r_n_328__38_,r_n_328__37_,
  r_n_328__36_,r_n_328__35_,r_n_328__34_,r_n_328__33_,r_n_328__32_,r_n_328__31_,
  r_n_328__30_,r_n_328__29_,r_n_328__28_,r_n_328__27_,r_n_328__26_,r_n_328__25_,
  r_n_328__24_,r_n_328__23_,r_n_328__22_,r_n_328__21_,r_n_328__20_,r_n_328__19_,
  r_n_328__18_,r_n_328__17_,r_n_328__16_,r_n_328__15_,r_n_328__14_,r_n_328__13_,
  r_n_328__12_,r_n_328__11_,r_n_328__10_,r_n_328__9_,r_n_328__8_,r_n_328__7_,r_n_328__6_,
  r_n_328__5_,r_n_328__4_,r_n_328__3_,r_n_328__2_,r_n_328__1_,r_n_328__0_,
  r_n_327__63_,r_n_327__62_,r_n_327__61_,r_n_327__60_,r_n_327__59_,r_n_327__58_,r_n_327__57_,
  r_n_327__56_,r_n_327__55_,r_n_327__54_,r_n_327__53_,r_n_327__52_,r_n_327__51_,
  r_n_327__50_,r_n_327__49_,r_n_327__48_,r_n_327__47_,r_n_327__46_,r_n_327__45_,
  r_n_327__44_,r_n_327__43_,r_n_327__42_,r_n_327__41_,r_n_327__40_,r_n_327__39_,
  r_n_327__38_,r_n_327__37_,r_n_327__36_,r_n_327__35_,r_n_327__34_,r_n_327__33_,
  r_n_327__32_,r_n_327__31_,r_n_327__30_,r_n_327__29_,r_n_327__28_,r_n_327__27_,
  r_n_327__26_,r_n_327__25_,r_n_327__24_,r_n_327__23_,r_n_327__22_,r_n_327__21_,r_n_327__20_,
  r_n_327__19_,r_n_327__18_,r_n_327__17_,r_n_327__16_,r_n_327__15_,r_n_327__14_,
  r_n_327__13_,r_n_327__12_,r_n_327__11_,r_n_327__10_,r_n_327__9_,r_n_327__8_,
  r_n_327__7_,r_n_327__6_,r_n_327__5_,r_n_327__4_,r_n_327__3_,r_n_327__2_,r_n_327__1_,
  r_n_327__0_,r_n_326__63_,r_n_326__62_,r_n_326__61_,r_n_326__60_,r_n_326__59_,
  r_n_326__58_,r_n_326__57_,r_n_326__56_,r_n_326__55_,r_n_326__54_,r_n_326__53_,
  r_n_326__52_,r_n_326__51_,r_n_326__50_,r_n_326__49_,r_n_326__48_,r_n_326__47_,
  r_n_326__46_,r_n_326__45_,r_n_326__44_,r_n_326__43_,r_n_326__42_,r_n_326__41_,
  r_n_326__40_,r_n_326__39_,r_n_326__38_,r_n_326__37_,r_n_326__36_,r_n_326__35_,r_n_326__34_,
  r_n_326__33_,r_n_326__32_,r_n_326__31_,r_n_326__30_,r_n_326__29_,r_n_326__28_,
  r_n_326__27_,r_n_326__26_,r_n_326__25_,r_n_326__24_,r_n_326__23_,r_n_326__22_,
  r_n_326__21_,r_n_326__20_,r_n_326__19_,r_n_326__18_,r_n_326__17_,r_n_326__16_,
  r_n_326__15_,r_n_326__14_,r_n_326__13_,r_n_326__12_,r_n_326__11_,r_n_326__10_,
  r_n_326__9_,r_n_326__8_,r_n_326__7_,r_n_326__6_,r_n_326__5_,r_n_326__4_,r_n_326__3_,
  r_n_326__2_,r_n_326__1_,r_n_326__0_,r_n_325__63_,r_n_325__62_,r_n_325__61_,
  r_n_325__60_,r_n_325__59_,r_n_325__58_,r_n_325__57_,r_n_325__56_,r_n_325__55_,
  r_n_325__54_,r_n_325__53_,r_n_325__52_,r_n_325__51_,r_n_325__50_,r_n_325__49_,r_n_325__48_,
  r_n_325__47_,r_n_325__46_,r_n_325__45_,r_n_325__44_,r_n_325__43_,r_n_325__42_,
  r_n_325__41_,r_n_325__40_,r_n_325__39_,r_n_325__38_,r_n_325__37_,r_n_325__36_,
  r_n_325__35_,r_n_325__34_,r_n_325__33_,r_n_325__32_,r_n_325__31_,r_n_325__30_,
  r_n_325__29_,r_n_325__28_,r_n_325__27_,r_n_325__26_,r_n_325__25_,r_n_325__24_,
  r_n_325__23_,r_n_325__22_,r_n_325__21_,r_n_325__20_,r_n_325__19_,r_n_325__18_,
  r_n_325__17_,r_n_325__16_,r_n_325__15_,r_n_325__14_,r_n_325__13_,r_n_325__12_,
  r_n_325__11_,r_n_325__10_,r_n_325__9_,r_n_325__8_,r_n_325__7_,r_n_325__6_,r_n_325__5_,
  r_n_325__4_,r_n_325__3_,r_n_325__2_,r_n_325__1_,r_n_325__0_,r_n_324__63_,r_n_324__62_,
  r_n_324__61_,r_n_324__60_,r_n_324__59_,r_n_324__58_,r_n_324__57_,r_n_324__56_,
  r_n_324__55_,r_n_324__54_,r_n_324__53_,r_n_324__52_,r_n_324__51_,r_n_324__50_,
  r_n_324__49_,r_n_324__48_,r_n_324__47_,r_n_324__46_,r_n_324__45_,r_n_324__44_,
  r_n_324__43_,r_n_324__42_,r_n_324__41_,r_n_324__40_,r_n_324__39_,r_n_324__38_,
  r_n_324__37_,r_n_324__36_,r_n_324__35_,r_n_324__34_,r_n_324__33_,r_n_324__32_,
  r_n_324__31_,r_n_324__30_,r_n_324__29_,r_n_324__28_,r_n_324__27_,r_n_324__26_,
  r_n_324__25_,r_n_324__24_,r_n_324__23_,r_n_324__22_,r_n_324__21_,r_n_324__20_,r_n_324__19_,
  r_n_324__18_,r_n_324__17_,r_n_324__16_,r_n_324__15_,r_n_324__14_,r_n_324__13_,
  r_n_324__12_,r_n_324__11_,r_n_324__10_,r_n_324__9_,r_n_324__8_,r_n_324__7_,
  r_n_324__6_,r_n_324__5_,r_n_324__4_,r_n_324__3_,r_n_324__2_,r_n_324__1_,r_n_324__0_,
  r_n_323__63_,r_n_323__62_,r_n_323__61_,r_n_323__60_,r_n_323__59_,r_n_323__58_,
  r_n_323__57_,r_n_323__56_,r_n_323__55_,r_n_323__54_,r_n_323__53_,r_n_323__52_,
  r_n_323__51_,r_n_323__50_,r_n_323__49_,r_n_323__48_,r_n_323__47_,r_n_323__46_,
  r_n_323__45_,r_n_323__44_,r_n_323__43_,r_n_323__42_,r_n_323__41_,r_n_323__40_,
  r_n_323__39_,r_n_323__38_,r_n_323__37_,r_n_323__36_,r_n_323__35_,r_n_323__34_,r_n_323__33_,
  r_n_323__32_,r_n_323__31_,r_n_323__30_,r_n_323__29_,r_n_323__28_,r_n_323__27_,
  r_n_323__26_,r_n_323__25_,r_n_323__24_,r_n_323__23_,r_n_323__22_,r_n_323__21_,
  r_n_323__20_,r_n_323__19_,r_n_323__18_,r_n_323__17_,r_n_323__16_,r_n_323__15_,
  r_n_323__14_,r_n_323__13_,r_n_323__12_,r_n_323__11_,r_n_323__10_,r_n_323__9_,
  r_n_323__8_,r_n_323__7_,r_n_323__6_,r_n_323__5_,r_n_323__4_,r_n_323__3_,r_n_323__2_,
  r_n_323__1_,r_n_323__0_,r_n_322__63_,r_n_322__62_,r_n_322__61_,r_n_322__60_,
  r_n_322__59_,r_n_322__58_,r_n_322__57_,r_n_322__56_,r_n_322__55_,r_n_322__54_,
  r_n_322__53_,r_n_322__52_,r_n_322__51_,r_n_322__50_,r_n_322__49_,r_n_322__48_,r_n_322__47_,
  r_n_322__46_,r_n_322__45_,r_n_322__44_,r_n_322__43_,r_n_322__42_,r_n_322__41_,
  r_n_322__40_,r_n_322__39_,r_n_322__38_,r_n_322__37_,r_n_322__36_,r_n_322__35_,
  r_n_322__34_,r_n_322__33_,r_n_322__32_,r_n_322__31_,r_n_322__30_,r_n_322__29_,
  r_n_322__28_,r_n_322__27_,r_n_322__26_,r_n_322__25_,r_n_322__24_,r_n_322__23_,
  r_n_322__22_,r_n_322__21_,r_n_322__20_,r_n_322__19_,r_n_322__18_,r_n_322__17_,
  r_n_322__16_,r_n_322__15_,r_n_322__14_,r_n_322__13_,r_n_322__12_,r_n_322__11_,r_n_322__10_,
  r_n_322__9_,r_n_322__8_,r_n_322__7_,r_n_322__6_,r_n_322__5_,r_n_322__4_,
  r_n_322__3_,r_n_322__2_,r_n_322__1_,r_n_322__0_,r_n_321__63_,r_n_321__62_,r_n_321__61_,
  r_n_321__60_,r_n_321__59_,r_n_321__58_,r_n_321__57_,r_n_321__56_,r_n_321__55_,
  r_n_321__54_,r_n_321__53_,r_n_321__52_,r_n_321__51_,r_n_321__50_,r_n_321__49_,
  r_n_321__48_,r_n_321__47_,r_n_321__46_,r_n_321__45_,r_n_321__44_,r_n_321__43_,
  r_n_321__42_,r_n_321__41_,r_n_321__40_,r_n_321__39_,r_n_321__38_,r_n_321__37_,
  r_n_321__36_,r_n_321__35_,r_n_321__34_,r_n_321__33_,r_n_321__32_,r_n_321__31_,
  r_n_321__30_,r_n_321__29_,r_n_321__28_,r_n_321__27_,r_n_321__26_,r_n_321__25_,r_n_321__24_,
  r_n_321__23_,r_n_321__22_,r_n_321__21_,r_n_321__20_,r_n_321__19_,r_n_321__18_,
  r_n_321__17_,r_n_321__16_,r_n_321__15_,r_n_321__14_,r_n_321__13_,r_n_321__12_,
  r_n_321__11_,r_n_321__10_,r_n_321__9_,r_n_321__8_,r_n_321__7_,r_n_321__6_,
  r_n_321__5_,r_n_321__4_,r_n_321__3_,r_n_321__2_,r_n_321__1_,r_n_321__0_,r_n_336__63_,
  r_n_336__62_,r_n_336__61_,r_n_336__60_,r_n_336__59_,r_n_336__58_,r_n_336__57_,
  r_n_336__56_,r_n_336__55_,r_n_336__54_,r_n_336__53_,r_n_336__52_,r_n_336__51_,
  r_n_336__50_,r_n_336__49_,r_n_336__48_,r_n_336__47_,r_n_336__46_,r_n_336__45_,
  r_n_336__44_,r_n_336__43_,r_n_336__42_,r_n_336__41_,r_n_336__40_,r_n_336__39_,r_n_336__38_,
  r_n_336__37_,r_n_336__36_,r_n_336__35_,r_n_336__34_,r_n_336__33_,r_n_336__32_,
  r_n_336__31_,r_n_336__30_,r_n_336__29_,r_n_336__28_,r_n_336__27_,r_n_336__26_,
  r_n_336__25_,r_n_336__24_,r_n_336__23_,r_n_336__22_,r_n_336__21_,r_n_336__20_,
  r_n_336__19_,r_n_336__18_,r_n_336__17_,r_n_336__16_,r_n_336__15_,r_n_336__14_,
  r_n_336__13_,r_n_336__12_,r_n_336__11_,r_n_336__10_,r_n_336__9_,r_n_336__8_,r_n_336__7_,
  r_n_336__6_,r_n_336__5_,r_n_336__4_,r_n_336__3_,r_n_336__2_,r_n_336__1_,
  r_n_336__0_,r_n_335__63_,r_n_335__62_,r_n_335__61_,r_n_335__60_,r_n_335__59_,
  r_n_335__58_,r_n_335__57_,r_n_335__56_,r_n_335__55_,r_n_335__54_,r_n_335__53_,r_n_335__52_,
  r_n_335__51_,r_n_335__50_,r_n_335__49_,r_n_335__48_,r_n_335__47_,r_n_335__46_,
  r_n_335__45_,r_n_335__44_,r_n_335__43_,r_n_335__42_,r_n_335__41_,r_n_335__40_,
  r_n_335__39_,r_n_335__38_,r_n_335__37_,r_n_335__36_,r_n_335__35_,r_n_335__34_,
  r_n_335__33_,r_n_335__32_,r_n_335__31_,r_n_335__30_,r_n_335__29_,r_n_335__28_,
  r_n_335__27_,r_n_335__26_,r_n_335__25_,r_n_335__24_,r_n_335__23_,r_n_335__22_,
  r_n_335__21_,r_n_335__20_,r_n_335__19_,r_n_335__18_,r_n_335__17_,r_n_335__16_,
  r_n_335__15_,r_n_335__14_,r_n_335__13_,r_n_335__12_,r_n_335__11_,r_n_335__10_,r_n_335__9_,
  r_n_335__8_,r_n_335__7_,r_n_335__6_,r_n_335__5_,r_n_335__4_,r_n_335__3_,
  r_n_335__2_,r_n_335__1_,r_n_335__0_,r_n_334__63_,r_n_334__62_,r_n_334__61_,r_n_334__60_,
  r_n_334__59_,r_n_334__58_,r_n_334__57_,r_n_334__56_,r_n_334__55_,r_n_334__54_,
  r_n_334__53_,r_n_334__52_,r_n_334__51_,r_n_334__50_,r_n_334__49_,r_n_334__48_,
  r_n_334__47_,r_n_334__46_,r_n_334__45_,r_n_334__44_,r_n_334__43_,r_n_334__42_,
  r_n_334__41_,r_n_334__40_,r_n_334__39_,r_n_334__38_,r_n_334__37_,r_n_334__36_,
  r_n_334__35_,r_n_334__34_,r_n_334__33_,r_n_334__32_,r_n_334__31_,r_n_334__30_,
  r_n_334__29_,r_n_334__28_,r_n_334__27_,r_n_334__26_,r_n_334__25_,r_n_334__24_,r_n_334__23_,
  r_n_334__22_,r_n_334__21_,r_n_334__20_,r_n_334__19_,r_n_334__18_,r_n_334__17_,
  r_n_334__16_,r_n_334__15_,r_n_334__14_,r_n_334__13_,r_n_334__12_,r_n_334__11_,
  r_n_334__10_,r_n_334__9_,r_n_334__8_,r_n_334__7_,r_n_334__6_,r_n_334__5_,r_n_334__4_,
  r_n_334__3_,r_n_334__2_,r_n_334__1_,r_n_334__0_,r_n_333__63_,r_n_333__62_,
  r_n_333__61_,r_n_333__60_,r_n_333__59_,r_n_333__58_,r_n_333__57_,r_n_333__56_,
  r_n_333__55_,r_n_333__54_,r_n_333__53_,r_n_333__52_,r_n_333__51_,r_n_333__50_,
  r_n_333__49_,r_n_333__48_,r_n_333__47_,r_n_333__46_,r_n_333__45_,r_n_333__44_,
  r_n_333__43_,r_n_333__42_,r_n_333__41_,r_n_333__40_,r_n_333__39_,r_n_333__38_,r_n_333__37_,
  r_n_333__36_,r_n_333__35_,r_n_333__34_,r_n_333__33_,r_n_333__32_,r_n_333__31_,
  r_n_333__30_,r_n_333__29_,r_n_333__28_,r_n_333__27_,r_n_333__26_,r_n_333__25_,
  r_n_333__24_,r_n_333__23_,r_n_333__22_,r_n_333__21_,r_n_333__20_,r_n_333__19_,
  r_n_333__18_,r_n_333__17_,r_n_333__16_,r_n_333__15_,r_n_333__14_,r_n_333__13_,
  r_n_333__12_,r_n_333__11_,r_n_333__10_,r_n_333__9_,r_n_333__8_,r_n_333__7_,r_n_333__6_,
  r_n_333__5_,r_n_333__4_,r_n_333__3_,r_n_333__2_,r_n_333__1_,r_n_333__0_,
  r_n_332__63_,r_n_332__62_,r_n_332__61_,r_n_332__60_,r_n_332__59_,r_n_332__58_,
  r_n_332__57_,r_n_332__56_,r_n_332__55_,r_n_332__54_,r_n_332__53_,r_n_332__52_,r_n_332__51_,
  r_n_332__50_,r_n_332__49_,r_n_332__48_,r_n_332__47_,r_n_332__46_,r_n_332__45_,
  r_n_332__44_,r_n_332__43_,r_n_332__42_,r_n_332__41_,r_n_332__40_,r_n_332__39_,
  r_n_332__38_,r_n_332__37_,r_n_332__36_,r_n_332__35_,r_n_332__34_,r_n_332__33_,
  r_n_332__32_,r_n_332__31_,r_n_332__30_,r_n_332__29_,r_n_332__28_,r_n_332__27_,
  r_n_332__26_,r_n_332__25_,r_n_332__24_,r_n_332__23_,r_n_332__22_,r_n_332__21_,
  r_n_332__20_,r_n_332__19_,r_n_332__18_,r_n_332__17_,r_n_332__16_,r_n_332__15_,r_n_332__14_,
  r_n_332__13_,r_n_332__12_,r_n_332__11_,r_n_332__10_,r_n_332__9_,r_n_332__8_,
  r_n_332__7_,r_n_332__6_,r_n_332__5_,r_n_332__4_,r_n_332__3_,r_n_332__2_,r_n_332__1_,
  r_n_332__0_,r_n_331__63_,r_n_331__62_,r_n_331__61_,r_n_331__60_,r_n_331__59_,
  r_n_331__58_,r_n_331__57_,r_n_331__56_,r_n_331__55_,r_n_331__54_,r_n_331__53_,
  r_n_331__52_,r_n_331__51_,r_n_331__50_,r_n_331__49_,r_n_331__48_,r_n_331__47_,
  r_n_331__46_,r_n_331__45_,r_n_331__44_,r_n_331__43_,r_n_331__42_,r_n_331__41_,
  r_n_331__40_,r_n_331__39_,r_n_331__38_,r_n_331__37_,r_n_331__36_,r_n_331__35_,
  r_n_331__34_,r_n_331__33_,r_n_331__32_,r_n_331__31_,r_n_331__30_,r_n_331__29_,r_n_331__28_,
  r_n_331__27_,r_n_331__26_,r_n_331__25_,r_n_331__24_,r_n_331__23_,r_n_331__22_,
  r_n_331__21_,r_n_331__20_,r_n_331__19_,r_n_331__18_,r_n_331__17_,r_n_331__16_,
  r_n_331__15_,r_n_331__14_,r_n_331__13_,r_n_331__12_,r_n_331__11_,r_n_331__10_,
  r_n_331__9_,r_n_331__8_,r_n_331__7_,r_n_331__6_,r_n_331__5_,r_n_331__4_,r_n_331__3_,
  r_n_331__2_,r_n_331__1_,r_n_331__0_,r_n_330__63_,r_n_330__62_,r_n_330__61_,
  r_n_330__60_,r_n_330__59_,r_n_330__58_,r_n_330__57_,r_n_330__56_,r_n_330__55_,
  r_n_330__54_,r_n_330__53_,r_n_330__52_,r_n_330__51_,r_n_330__50_,r_n_330__49_,
  r_n_330__48_,r_n_330__47_,r_n_330__46_,r_n_330__45_,r_n_330__44_,r_n_330__43_,r_n_330__42_,
  r_n_330__41_,r_n_330__40_,r_n_330__39_,r_n_330__38_,r_n_330__37_,r_n_330__36_,
  r_n_330__35_,r_n_330__34_,r_n_330__33_,r_n_330__32_,r_n_330__31_,r_n_330__30_,
  r_n_330__29_,r_n_330__28_,r_n_330__27_,r_n_330__26_,r_n_330__25_,r_n_330__24_,
  r_n_330__23_,r_n_330__22_,r_n_330__21_,r_n_330__20_,r_n_330__19_,r_n_330__18_,
  r_n_330__17_,r_n_330__16_,r_n_330__15_,r_n_330__14_,r_n_330__13_,r_n_330__12_,
  r_n_330__11_,r_n_330__10_,r_n_330__9_,r_n_330__8_,r_n_330__7_,r_n_330__6_,r_n_330__5_,
  r_n_330__4_,r_n_330__3_,r_n_330__2_,r_n_330__1_,r_n_330__0_,r_n_329__63_,
  r_n_329__62_,r_n_329__61_,r_n_329__60_,r_n_329__59_,r_n_329__58_,r_n_329__57_,r_n_329__56_,
  r_n_329__55_,r_n_329__54_,r_n_329__53_,r_n_329__52_,r_n_329__51_,r_n_329__50_,
  r_n_329__49_,r_n_329__48_,r_n_329__47_,r_n_329__46_,r_n_329__45_,r_n_329__44_,
  r_n_329__43_,r_n_329__42_,r_n_329__41_,r_n_329__40_,r_n_329__39_,r_n_329__38_,
  r_n_329__37_,r_n_329__36_,r_n_329__35_,r_n_329__34_,r_n_329__33_,r_n_329__32_,
  r_n_329__31_,r_n_329__30_,r_n_329__29_,r_n_329__28_,r_n_329__27_,r_n_329__26_,
  r_n_329__25_,r_n_329__24_,r_n_329__23_,r_n_329__22_,r_n_329__21_,r_n_329__20_,
  r_n_329__19_,r_n_329__18_,r_n_329__17_,r_n_329__16_,r_n_329__15_,r_n_329__14_,r_n_329__13_,
  r_n_329__12_,r_n_329__11_,r_n_329__10_,r_n_329__9_,r_n_329__8_,r_n_329__7_,
  r_n_329__6_,r_n_329__5_,r_n_329__4_,r_n_329__3_,r_n_329__2_,r_n_329__1_,r_n_329__0_,
  r_n_344__63_,r_n_344__62_,r_n_344__61_,r_n_344__60_,r_n_344__59_,r_n_344__58_,
  r_n_344__57_,r_n_344__56_,r_n_344__55_,r_n_344__54_,r_n_344__53_,r_n_344__52_,
  r_n_344__51_,r_n_344__50_,r_n_344__49_,r_n_344__48_,r_n_344__47_,r_n_344__46_,
  r_n_344__45_,r_n_344__44_,r_n_344__43_,r_n_344__42_,r_n_344__41_,r_n_344__40_,
  r_n_344__39_,r_n_344__38_,r_n_344__37_,r_n_344__36_,r_n_344__35_,r_n_344__34_,
  r_n_344__33_,r_n_344__32_,r_n_344__31_,r_n_344__30_,r_n_344__29_,r_n_344__28_,r_n_344__27_,
  r_n_344__26_,r_n_344__25_,r_n_344__24_,r_n_344__23_,r_n_344__22_,r_n_344__21_,
  r_n_344__20_,r_n_344__19_,r_n_344__18_,r_n_344__17_,r_n_344__16_,r_n_344__15_,
  r_n_344__14_,r_n_344__13_,r_n_344__12_,r_n_344__11_,r_n_344__10_,r_n_344__9_,
  r_n_344__8_,r_n_344__7_,r_n_344__6_,r_n_344__5_,r_n_344__4_,r_n_344__3_,r_n_344__2_,
  r_n_344__1_,r_n_344__0_,r_n_343__63_,r_n_343__62_,r_n_343__61_,r_n_343__60_,
  r_n_343__59_,r_n_343__58_,r_n_343__57_,r_n_343__56_,r_n_343__55_,r_n_343__54_,
  r_n_343__53_,r_n_343__52_,r_n_343__51_,r_n_343__50_,r_n_343__49_,r_n_343__48_,
  r_n_343__47_,r_n_343__46_,r_n_343__45_,r_n_343__44_,r_n_343__43_,r_n_343__42_,r_n_343__41_,
  r_n_343__40_,r_n_343__39_,r_n_343__38_,r_n_343__37_,r_n_343__36_,r_n_343__35_,
  r_n_343__34_,r_n_343__33_,r_n_343__32_,r_n_343__31_,r_n_343__30_,r_n_343__29_,
  r_n_343__28_,r_n_343__27_,r_n_343__26_,r_n_343__25_,r_n_343__24_,r_n_343__23_,
  r_n_343__22_,r_n_343__21_,r_n_343__20_,r_n_343__19_,r_n_343__18_,r_n_343__17_,
  r_n_343__16_,r_n_343__15_,r_n_343__14_,r_n_343__13_,r_n_343__12_,r_n_343__11_,
  r_n_343__10_,r_n_343__9_,r_n_343__8_,r_n_343__7_,r_n_343__6_,r_n_343__5_,r_n_343__4_,
  r_n_343__3_,r_n_343__2_,r_n_343__1_,r_n_343__0_,r_n_342__63_,r_n_342__62_,
  r_n_342__61_,r_n_342__60_,r_n_342__59_,r_n_342__58_,r_n_342__57_,r_n_342__56_,r_n_342__55_,
  r_n_342__54_,r_n_342__53_,r_n_342__52_,r_n_342__51_,r_n_342__50_,r_n_342__49_,
  r_n_342__48_,r_n_342__47_,r_n_342__46_,r_n_342__45_,r_n_342__44_,r_n_342__43_,
  r_n_342__42_,r_n_342__41_,r_n_342__40_,r_n_342__39_,r_n_342__38_,r_n_342__37_,
  r_n_342__36_,r_n_342__35_,r_n_342__34_,r_n_342__33_,r_n_342__32_,r_n_342__31_,
  r_n_342__30_,r_n_342__29_,r_n_342__28_,r_n_342__27_,r_n_342__26_,r_n_342__25_,
  r_n_342__24_,r_n_342__23_,r_n_342__22_,r_n_342__21_,r_n_342__20_,r_n_342__19_,r_n_342__18_,
  r_n_342__17_,r_n_342__16_,r_n_342__15_,r_n_342__14_,r_n_342__13_,r_n_342__12_,
  r_n_342__11_,r_n_342__10_,r_n_342__9_,r_n_342__8_,r_n_342__7_,r_n_342__6_,
  r_n_342__5_,r_n_342__4_,r_n_342__3_,r_n_342__2_,r_n_342__1_,r_n_342__0_,r_n_341__63_,
  r_n_341__62_,r_n_341__61_,r_n_341__60_,r_n_341__59_,r_n_341__58_,r_n_341__57_,
  r_n_341__56_,r_n_341__55_,r_n_341__54_,r_n_341__53_,r_n_341__52_,r_n_341__51_,
  r_n_341__50_,r_n_341__49_,r_n_341__48_,r_n_341__47_,r_n_341__46_,r_n_341__45_,
  r_n_341__44_,r_n_341__43_,r_n_341__42_,r_n_341__41_,r_n_341__40_,r_n_341__39_,
  r_n_341__38_,r_n_341__37_,r_n_341__36_,r_n_341__35_,r_n_341__34_,r_n_341__33_,r_n_341__32_,
  r_n_341__31_,r_n_341__30_,r_n_341__29_,r_n_341__28_,r_n_341__27_,r_n_341__26_,
  r_n_341__25_,r_n_341__24_,r_n_341__23_,r_n_341__22_,r_n_341__21_,r_n_341__20_,
  r_n_341__19_,r_n_341__18_,r_n_341__17_,r_n_341__16_,r_n_341__15_,r_n_341__14_,
  r_n_341__13_,r_n_341__12_,r_n_341__11_,r_n_341__10_,r_n_341__9_,r_n_341__8_,
  r_n_341__7_,r_n_341__6_,r_n_341__5_,r_n_341__4_,r_n_341__3_,r_n_341__2_,r_n_341__1_,
  r_n_341__0_,r_n_340__63_,r_n_340__62_,r_n_340__61_,r_n_340__60_,r_n_340__59_,
  r_n_340__58_,r_n_340__57_,r_n_340__56_,r_n_340__55_,r_n_340__54_,r_n_340__53_,
  r_n_340__52_,r_n_340__51_,r_n_340__50_,r_n_340__49_,r_n_340__48_,r_n_340__47_,r_n_340__46_,
  r_n_340__45_,r_n_340__44_,r_n_340__43_,r_n_340__42_,r_n_340__41_,r_n_340__40_,
  r_n_340__39_,r_n_340__38_,r_n_340__37_,r_n_340__36_,r_n_340__35_,r_n_340__34_,
  r_n_340__33_,r_n_340__32_,r_n_340__31_,r_n_340__30_,r_n_340__29_,r_n_340__28_,
  r_n_340__27_,r_n_340__26_,r_n_340__25_,r_n_340__24_,r_n_340__23_,r_n_340__22_,
  r_n_340__21_,r_n_340__20_,r_n_340__19_,r_n_340__18_,r_n_340__17_,r_n_340__16_,
  r_n_340__15_,r_n_340__14_,r_n_340__13_,r_n_340__12_,r_n_340__11_,r_n_340__10_,r_n_340__9_,
  r_n_340__8_,r_n_340__7_,r_n_340__6_,r_n_340__5_,r_n_340__4_,r_n_340__3_,
  r_n_340__2_,r_n_340__1_,r_n_340__0_,r_n_339__63_,r_n_339__62_,r_n_339__61_,r_n_339__60_,
  r_n_339__59_,r_n_339__58_,r_n_339__57_,r_n_339__56_,r_n_339__55_,r_n_339__54_,
  r_n_339__53_,r_n_339__52_,r_n_339__51_,r_n_339__50_,r_n_339__49_,r_n_339__48_,
  r_n_339__47_,r_n_339__46_,r_n_339__45_,r_n_339__44_,r_n_339__43_,r_n_339__42_,
  r_n_339__41_,r_n_339__40_,r_n_339__39_,r_n_339__38_,r_n_339__37_,r_n_339__36_,
  r_n_339__35_,r_n_339__34_,r_n_339__33_,r_n_339__32_,r_n_339__31_,r_n_339__30_,
  r_n_339__29_,r_n_339__28_,r_n_339__27_,r_n_339__26_,r_n_339__25_,r_n_339__24_,
  r_n_339__23_,r_n_339__22_,r_n_339__21_,r_n_339__20_,r_n_339__19_,r_n_339__18_,r_n_339__17_,
  r_n_339__16_,r_n_339__15_,r_n_339__14_,r_n_339__13_,r_n_339__12_,r_n_339__11_,
  r_n_339__10_,r_n_339__9_,r_n_339__8_,r_n_339__7_,r_n_339__6_,r_n_339__5_,
  r_n_339__4_,r_n_339__3_,r_n_339__2_,r_n_339__1_,r_n_339__0_,r_n_338__63_,r_n_338__62_,
  r_n_338__61_,r_n_338__60_,r_n_338__59_,r_n_338__58_,r_n_338__57_,r_n_338__56_,
  r_n_338__55_,r_n_338__54_,r_n_338__53_,r_n_338__52_,r_n_338__51_,r_n_338__50_,
  r_n_338__49_,r_n_338__48_,r_n_338__47_,r_n_338__46_,r_n_338__45_,r_n_338__44_,
  r_n_338__43_,r_n_338__42_,r_n_338__41_,r_n_338__40_,r_n_338__39_,r_n_338__38_,
  r_n_338__37_,r_n_338__36_,r_n_338__35_,r_n_338__34_,r_n_338__33_,r_n_338__32_,r_n_338__31_,
  r_n_338__30_,r_n_338__29_,r_n_338__28_,r_n_338__27_,r_n_338__26_,r_n_338__25_,
  r_n_338__24_,r_n_338__23_,r_n_338__22_,r_n_338__21_,r_n_338__20_,r_n_338__19_,
  r_n_338__18_,r_n_338__17_,r_n_338__16_,r_n_338__15_,r_n_338__14_,r_n_338__13_,
  r_n_338__12_,r_n_338__11_,r_n_338__10_,r_n_338__9_,r_n_338__8_,r_n_338__7_,r_n_338__6_,
  r_n_338__5_,r_n_338__4_,r_n_338__3_,r_n_338__2_,r_n_338__1_,r_n_338__0_,
  r_n_337__63_,r_n_337__62_,r_n_337__61_,r_n_337__60_,r_n_337__59_,r_n_337__58_,
  r_n_337__57_,r_n_337__56_,r_n_337__55_,r_n_337__54_,r_n_337__53_,r_n_337__52_,
  r_n_337__51_,r_n_337__50_,r_n_337__49_,r_n_337__48_,r_n_337__47_,r_n_337__46_,r_n_337__45_,
  r_n_337__44_,r_n_337__43_,r_n_337__42_,r_n_337__41_,r_n_337__40_,r_n_337__39_,
  r_n_337__38_,r_n_337__37_,r_n_337__36_,r_n_337__35_,r_n_337__34_,r_n_337__33_,
  r_n_337__32_,r_n_337__31_,r_n_337__30_,r_n_337__29_,r_n_337__28_,r_n_337__27_,
  r_n_337__26_,r_n_337__25_,r_n_337__24_,r_n_337__23_,r_n_337__22_,r_n_337__21_,
  r_n_337__20_,r_n_337__19_,r_n_337__18_,r_n_337__17_,r_n_337__16_,r_n_337__15_,
  r_n_337__14_,r_n_337__13_,r_n_337__12_,r_n_337__11_,r_n_337__10_,r_n_337__9_,r_n_337__8_,
  r_n_337__7_,r_n_337__6_,r_n_337__5_,r_n_337__4_,r_n_337__3_,r_n_337__2_,
  r_n_337__1_,r_n_337__0_,r_n_352__63_,r_n_352__62_,r_n_352__61_,r_n_352__60_,r_n_352__59_,
  r_n_352__58_,r_n_352__57_,r_n_352__56_,r_n_352__55_,r_n_352__54_,r_n_352__53_,
  r_n_352__52_,r_n_352__51_,r_n_352__50_,r_n_352__49_,r_n_352__48_,r_n_352__47_,
  r_n_352__46_,r_n_352__45_,r_n_352__44_,r_n_352__43_,r_n_352__42_,r_n_352__41_,
  r_n_352__40_,r_n_352__39_,r_n_352__38_,r_n_352__37_,r_n_352__36_,r_n_352__35_,
  r_n_352__34_,r_n_352__33_,r_n_352__32_,r_n_352__31_,r_n_352__30_,r_n_352__29_,
  r_n_352__28_,r_n_352__27_,r_n_352__26_,r_n_352__25_,r_n_352__24_,r_n_352__23_,r_n_352__22_,
  r_n_352__21_,r_n_352__20_,r_n_352__19_,r_n_352__18_,r_n_352__17_,r_n_352__16_,
  r_n_352__15_,r_n_352__14_,r_n_352__13_,r_n_352__12_,r_n_352__11_,r_n_352__10_,
  r_n_352__9_,r_n_352__8_,r_n_352__7_,r_n_352__6_,r_n_352__5_,r_n_352__4_,r_n_352__3_,
  r_n_352__2_,r_n_352__1_,r_n_352__0_,r_n_351__63_,r_n_351__62_,r_n_351__61_,
  r_n_351__60_,r_n_351__59_,r_n_351__58_,r_n_351__57_,r_n_351__56_,r_n_351__55_,
  r_n_351__54_,r_n_351__53_,r_n_351__52_,r_n_351__51_,r_n_351__50_,r_n_351__49_,
  r_n_351__48_,r_n_351__47_,r_n_351__46_,r_n_351__45_,r_n_351__44_,r_n_351__43_,
  r_n_351__42_,r_n_351__41_,r_n_351__40_,r_n_351__39_,r_n_351__38_,r_n_351__37_,r_n_351__36_,
  r_n_351__35_,r_n_351__34_,r_n_351__33_,r_n_351__32_,r_n_351__31_,r_n_351__30_,
  r_n_351__29_,r_n_351__28_,r_n_351__27_,r_n_351__26_,r_n_351__25_,r_n_351__24_,
  r_n_351__23_,r_n_351__22_,r_n_351__21_,r_n_351__20_,r_n_351__19_,r_n_351__18_,
  r_n_351__17_,r_n_351__16_,r_n_351__15_,r_n_351__14_,r_n_351__13_,r_n_351__12_,
  r_n_351__11_,r_n_351__10_,r_n_351__9_,r_n_351__8_,r_n_351__7_,r_n_351__6_,r_n_351__5_,
  r_n_351__4_,r_n_351__3_,r_n_351__2_,r_n_351__1_,r_n_351__0_,r_n_350__63_,
  r_n_350__62_,r_n_350__61_,r_n_350__60_,r_n_350__59_,r_n_350__58_,r_n_350__57_,
  r_n_350__56_,r_n_350__55_,r_n_350__54_,r_n_350__53_,r_n_350__52_,r_n_350__51_,r_n_350__50_,
  r_n_350__49_,r_n_350__48_,r_n_350__47_,r_n_350__46_,r_n_350__45_,r_n_350__44_,
  r_n_350__43_,r_n_350__42_,r_n_350__41_,r_n_350__40_,r_n_350__39_,r_n_350__38_,
  r_n_350__37_,r_n_350__36_,r_n_350__35_,r_n_350__34_,r_n_350__33_,r_n_350__32_,
  r_n_350__31_,r_n_350__30_,r_n_350__29_,r_n_350__28_,r_n_350__27_,r_n_350__26_,
  r_n_350__25_,r_n_350__24_,r_n_350__23_,r_n_350__22_,r_n_350__21_,r_n_350__20_,
  r_n_350__19_,r_n_350__18_,r_n_350__17_,r_n_350__16_,r_n_350__15_,r_n_350__14_,
  r_n_350__13_,r_n_350__12_,r_n_350__11_,r_n_350__10_,r_n_350__9_,r_n_350__8_,r_n_350__7_,
  r_n_350__6_,r_n_350__5_,r_n_350__4_,r_n_350__3_,r_n_350__2_,r_n_350__1_,r_n_350__0_,
  r_n_349__63_,r_n_349__62_,r_n_349__61_,r_n_349__60_,r_n_349__59_,r_n_349__58_,
  r_n_349__57_,r_n_349__56_,r_n_349__55_,r_n_349__54_,r_n_349__53_,r_n_349__52_,
  r_n_349__51_,r_n_349__50_,r_n_349__49_,r_n_349__48_,r_n_349__47_,r_n_349__46_,
  r_n_349__45_,r_n_349__44_,r_n_349__43_,r_n_349__42_,r_n_349__41_,r_n_349__40_,
  r_n_349__39_,r_n_349__38_,r_n_349__37_,r_n_349__36_,r_n_349__35_,r_n_349__34_,
  r_n_349__33_,r_n_349__32_,r_n_349__31_,r_n_349__30_,r_n_349__29_,r_n_349__28_,
  r_n_349__27_,r_n_349__26_,r_n_349__25_,r_n_349__24_,r_n_349__23_,r_n_349__22_,r_n_349__21_,
  r_n_349__20_,r_n_349__19_,r_n_349__18_,r_n_349__17_,r_n_349__16_,r_n_349__15_,
  r_n_349__14_,r_n_349__13_,r_n_349__12_,r_n_349__11_,r_n_349__10_,r_n_349__9_,
  r_n_349__8_,r_n_349__7_,r_n_349__6_,r_n_349__5_,r_n_349__4_,r_n_349__3_,r_n_349__2_,
  r_n_349__1_,r_n_349__0_,r_n_348__63_,r_n_348__62_,r_n_348__61_,r_n_348__60_,
  r_n_348__59_,r_n_348__58_,r_n_348__57_,r_n_348__56_,r_n_348__55_,r_n_348__54_,
  r_n_348__53_,r_n_348__52_,r_n_348__51_,r_n_348__50_,r_n_348__49_,r_n_348__48_,
  r_n_348__47_,r_n_348__46_,r_n_348__45_,r_n_348__44_,r_n_348__43_,r_n_348__42_,
  r_n_348__41_,r_n_348__40_,r_n_348__39_,r_n_348__38_,r_n_348__37_,r_n_348__36_,r_n_348__35_,
  r_n_348__34_,r_n_348__33_,r_n_348__32_,r_n_348__31_,r_n_348__30_,r_n_348__29_,
  r_n_348__28_,r_n_348__27_,r_n_348__26_,r_n_348__25_,r_n_348__24_,r_n_348__23_,
  r_n_348__22_,r_n_348__21_,r_n_348__20_,r_n_348__19_,r_n_348__18_,r_n_348__17_,
  r_n_348__16_,r_n_348__15_,r_n_348__14_,r_n_348__13_,r_n_348__12_,r_n_348__11_,
  r_n_348__10_,r_n_348__9_,r_n_348__8_,r_n_348__7_,r_n_348__6_,r_n_348__5_,r_n_348__4_,
  r_n_348__3_,r_n_348__2_,r_n_348__1_,r_n_348__0_,r_n_347__63_,r_n_347__62_,
  r_n_347__61_,r_n_347__60_,r_n_347__59_,r_n_347__58_,r_n_347__57_,r_n_347__56_,
  r_n_347__55_,r_n_347__54_,r_n_347__53_,r_n_347__52_,r_n_347__51_,r_n_347__50_,r_n_347__49_,
  r_n_347__48_,r_n_347__47_,r_n_347__46_,r_n_347__45_,r_n_347__44_,r_n_347__43_,
  r_n_347__42_,r_n_347__41_,r_n_347__40_,r_n_347__39_,r_n_347__38_,r_n_347__37_,
  r_n_347__36_,r_n_347__35_,r_n_347__34_,r_n_347__33_,r_n_347__32_,r_n_347__31_,
  r_n_347__30_,r_n_347__29_,r_n_347__28_,r_n_347__27_,r_n_347__26_,r_n_347__25_,
  r_n_347__24_,r_n_347__23_,r_n_347__22_,r_n_347__21_,r_n_347__20_,r_n_347__19_,
  r_n_347__18_,r_n_347__17_,r_n_347__16_,r_n_347__15_,r_n_347__14_,r_n_347__13_,r_n_347__12_,
  r_n_347__11_,r_n_347__10_,r_n_347__9_,r_n_347__8_,r_n_347__7_,r_n_347__6_,
  r_n_347__5_,r_n_347__4_,r_n_347__3_,r_n_347__2_,r_n_347__1_,r_n_347__0_,r_n_346__63_,
  r_n_346__62_,r_n_346__61_,r_n_346__60_,r_n_346__59_,r_n_346__58_,r_n_346__57_,
  r_n_346__56_,r_n_346__55_,r_n_346__54_,r_n_346__53_,r_n_346__52_,r_n_346__51_,
  r_n_346__50_,r_n_346__49_,r_n_346__48_,r_n_346__47_,r_n_346__46_,r_n_346__45_,
  r_n_346__44_,r_n_346__43_,r_n_346__42_,r_n_346__41_,r_n_346__40_,r_n_346__39_,
  r_n_346__38_,r_n_346__37_,r_n_346__36_,r_n_346__35_,r_n_346__34_,r_n_346__33_,
  r_n_346__32_,r_n_346__31_,r_n_346__30_,r_n_346__29_,r_n_346__28_,r_n_346__27_,r_n_346__26_,
  r_n_346__25_,r_n_346__24_,r_n_346__23_,r_n_346__22_,r_n_346__21_,r_n_346__20_,
  r_n_346__19_,r_n_346__18_,r_n_346__17_,r_n_346__16_,r_n_346__15_,r_n_346__14_,
  r_n_346__13_,r_n_346__12_,r_n_346__11_,r_n_346__10_,r_n_346__9_,r_n_346__8_,
  r_n_346__7_,r_n_346__6_,r_n_346__5_,r_n_346__4_,r_n_346__3_,r_n_346__2_,r_n_346__1_,
  r_n_346__0_,r_n_345__63_,r_n_345__62_,r_n_345__61_,r_n_345__60_,r_n_345__59_,
  r_n_345__58_,r_n_345__57_,r_n_345__56_,r_n_345__55_,r_n_345__54_,r_n_345__53_,
  r_n_345__52_,r_n_345__51_,r_n_345__50_,r_n_345__49_,r_n_345__48_,r_n_345__47_,
  r_n_345__46_,r_n_345__45_,r_n_345__44_,r_n_345__43_,r_n_345__42_,r_n_345__41_,r_n_345__40_,
  r_n_345__39_,r_n_345__38_,r_n_345__37_,r_n_345__36_,r_n_345__35_,r_n_345__34_,
  r_n_345__33_,r_n_345__32_,r_n_345__31_,r_n_345__30_,r_n_345__29_,r_n_345__28_,
  r_n_345__27_,r_n_345__26_,r_n_345__25_,r_n_345__24_,r_n_345__23_,r_n_345__22_,
  r_n_345__21_,r_n_345__20_,r_n_345__19_,r_n_345__18_,r_n_345__17_,r_n_345__16_,
  r_n_345__15_,r_n_345__14_,r_n_345__13_,r_n_345__12_,r_n_345__11_,r_n_345__10_,
  r_n_345__9_,r_n_345__8_,r_n_345__7_,r_n_345__6_,r_n_345__5_,r_n_345__4_,r_n_345__3_,
  r_n_345__2_,r_n_345__1_,r_n_345__0_,r_n_360__63_,r_n_360__62_,r_n_360__61_,
  r_n_360__60_,r_n_360__59_,r_n_360__58_,r_n_360__57_,r_n_360__56_,r_n_360__55_,r_n_360__54_,
  r_n_360__53_,r_n_360__52_,r_n_360__51_,r_n_360__50_,r_n_360__49_,r_n_360__48_,
  r_n_360__47_,r_n_360__46_,r_n_360__45_,r_n_360__44_,r_n_360__43_,r_n_360__42_,
  r_n_360__41_,r_n_360__40_,r_n_360__39_,r_n_360__38_,r_n_360__37_,r_n_360__36_,
  r_n_360__35_,r_n_360__34_,r_n_360__33_,r_n_360__32_,r_n_360__31_,r_n_360__30_,
  r_n_360__29_,r_n_360__28_,r_n_360__27_,r_n_360__26_,r_n_360__25_,r_n_360__24_,
  r_n_360__23_,r_n_360__22_,r_n_360__21_,r_n_360__20_,r_n_360__19_,r_n_360__18_,
  r_n_360__17_,r_n_360__16_,r_n_360__15_,r_n_360__14_,r_n_360__13_,r_n_360__12_,r_n_360__11_,
  r_n_360__10_,r_n_360__9_,r_n_360__8_,r_n_360__7_,r_n_360__6_,r_n_360__5_,
  r_n_360__4_,r_n_360__3_,r_n_360__2_,r_n_360__1_,r_n_360__0_,r_n_359__63_,r_n_359__62_,
  r_n_359__61_,r_n_359__60_,r_n_359__59_,r_n_359__58_,r_n_359__57_,r_n_359__56_,
  r_n_359__55_,r_n_359__54_,r_n_359__53_,r_n_359__52_,r_n_359__51_,r_n_359__50_,
  r_n_359__49_,r_n_359__48_,r_n_359__47_,r_n_359__46_,r_n_359__45_,r_n_359__44_,
  r_n_359__43_,r_n_359__42_,r_n_359__41_,r_n_359__40_,r_n_359__39_,r_n_359__38_,
  r_n_359__37_,r_n_359__36_,r_n_359__35_,r_n_359__34_,r_n_359__33_,r_n_359__32_,
  r_n_359__31_,r_n_359__30_,r_n_359__29_,r_n_359__28_,r_n_359__27_,r_n_359__26_,r_n_359__25_,
  r_n_359__24_,r_n_359__23_,r_n_359__22_,r_n_359__21_,r_n_359__20_,r_n_359__19_,
  r_n_359__18_,r_n_359__17_,r_n_359__16_,r_n_359__15_,r_n_359__14_,r_n_359__13_,
  r_n_359__12_,r_n_359__11_,r_n_359__10_,r_n_359__9_,r_n_359__8_,r_n_359__7_,
  r_n_359__6_,r_n_359__5_,r_n_359__4_,r_n_359__3_,r_n_359__2_,r_n_359__1_,r_n_359__0_,
  r_n_358__63_,r_n_358__62_,r_n_358__61_,r_n_358__60_,r_n_358__59_,r_n_358__58_,
  r_n_358__57_,r_n_358__56_,r_n_358__55_,r_n_358__54_,r_n_358__53_,r_n_358__52_,
  r_n_358__51_,r_n_358__50_,r_n_358__49_,r_n_358__48_,r_n_358__47_,r_n_358__46_,
  r_n_358__45_,r_n_358__44_,r_n_358__43_,r_n_358__42_,r_n_358__41_,r_n_358__40_,r_n_358__39_,
  r_n_358__38_,r_n_358__37_,r_n_358__36_,r_n_358__35_,r_n_358__34_,r_n_358__33_,
  r_n_358__32_,r_n_358__31_,r_n_358__30_,r_n_358__29_,r_n_358__28_,r_n_358__27_,
  r_n_358__26_,r_n_358__25_,r_n_358__24_,r_n_358__23_,r_n_358__22_,r_n_358__21_,
  r_n_358__20_,r_n_358__19_,r_n_358__18_,r_n_358__17_,r_n_358__16_,r_n_358__15_,
  r_n_358__14_,r_n_358__13_,r_n_358__12_,r_n_358__11_,r_n_358__10_,r_n_358__9_,r_n_358__8_,
  r_n_358__7_,r_n_358__6_,r_n_358__5_,r_n_358__4_,r_n_358__3_,r_n_358__2_,
  r_n_358__1_,r_n_358__0_,r_n_357__63_,r_n_357__62_,r_n_357__61_,r_n_357__60_,
  r_n_357__59_,r_n_357__58_,r_n_357__57_,r_n_357__56_,r_n_357__55_,r_n_357__54_,r_n_357__53_,
  r_n_357__52_,r_n_357__51_,r_n_357__50_,r_n_357__49_,r_n_357__48_,r_n_357__47_,
  r_n_357__46_,r_n_357__45_,r_n_357__44_,r_n_357__43_,r_n_357__42_,r_n_357__41_,
  r_n_357__40_,r_n_357__39_,r_n_357__38_,r_n_357__37_,r_n_357__36_,r_n_357__35_,
  r_n_357__34_,r_n_357__33_,r_n_357__32_,r_n_357__31_,r_n_357__30_,r_n_357__29_,
  r_n_357__28_,r_n_357__27_,r_n_357__26_,r_n_357__25_,r_n_357__24_,r_n_357__23_,
  r_n_357__22_,r_n_357__21_,r_n_357__20_,r_n_357__19_,r_n_357__18_,r_n_357__17_,r_n_357__16_,
  r_n_357__15_,r_n_357__14_,r_n_357__13_,r_n_357__12_,r_n_357__11_,r_n_357__10_,
  r_n_357__9_,r_n_357__8_,r_n_357__7_,r_n_357__6_,r_n_357__5_,r_n_357__4_,
  r_n_357__3_,r_n_357__2_,r_n_357__1_,r_n_357__0_,r_n_356__63_,r_n_356__62_,r_n_356__61_,
  r_n_356__60_,r_n_356__59_,r_n_356__58_,r_n_356__57_,r_n_356__56_,r_n_356__55_,
  r_n_356__54_,r_n_356__53_,r_n_356__52_,r_n_356__51_,r_n_356__50_,r_n_356__49_,
  r_n_356__48_,r_n_356__47_,r_n_356__46_,r_n_356__45_,r_n_356__44_,r_n_356__43_,
  r_n_356__42_,r_n_356__41_,r_n_356__40_,r_n_356__39_,r_n_356__38_,r_n_356__37_,
  r_n_356__36_,r_n_356__35_,r_n_356__34_,r_n_356__33_,r_n_356__32_,r_n_356__31_,r_n_356__30_,
  r_n_356__29_,r_n_356__28_,r_n_356__27_,r_n_356__26_,r_n_356__25_,r_n_356__24_,
  r_n_356__23_,r_n_356__22_,r_n_356__21_,r_n_356__20_,r_n_356__19_,r_n_356__18_,
  r_n_356__17_,r_n_356__16_,r_n_356__15_,r_n_356__14_,r_n_356__13_,r_n_356__12_,
  r_n_356__11_,r_n_356__10_,r_n_356__9_,r_n_356__8_,r_n_356__7_,r_n_356__6_,r_n_356__5_,
  r_n_356__4_,r_n_356__3_,r_n_356__2_,r_n_356__1_,r_n_356__0_,r_n_355__63_,
  r_n_355__62_,r_n_355__61_,r_n_355__60_,r_n_355__59_,r_n_355__58_,r_n_355__57_,
  r_n_355__56_,r_n_355__55_,r_n_355__54_,r_n_355__53_,r_n_355__52_,r_n_355__51_,
  r_n_355__50_,r_n_355__49_,r_n_355__48_,r_n_355__47_,r_n_355__46_,r_n_355__45_,r_n_355__44_,
  r_n_355__43_,r_n_355__42_,r_n_355__41_,r_n_355__40_,r_n_355__39_,r_n_355__38_,
  r_n_355__37_,r_n_355__36_,r_n_355__35_,r_n_355__34_,r_n_355__33_,r_n_355__32_,
  r_n_355__31_,r_n_355__30_,r_n_355__29_,r_n_355__28_,r_n_355__27_,r_n_355__26_,
  r_n_355__25_,r_n_355__24_,r_n_355__23_,r_n_355__22_,r_n_355__21_,r_n_355__20_,
  r_n_355__19_,r_n_355__18_,r_n_355__17_,r_n_355__16_,r_n_355__15_,r_n_355__14_,
  r_n_355__13_,r_n_355__12_,r_n_355__11_,r_n_355__10_,r_n_355__9_,r_n_355__8_,r_n_355__7_,
  r_n_355__6_,r_n_355__5_,r_n_355__4_,r_n_355__3_,r_n_355__2_,r_n_355__1_,
  r_n_355__0_,r_n_354__63_,r_n_354__62_,r_n_354__61_,r_n_354__60_,r_n_354__59_,r_n_354__58_,
  r_n_354__57_,r_n_354__56_,r_n_354__55_,r_n_354__54_,r_n_354__53_,r_n_354__52_,
  r_n_354__51_,r_n_354__50_,r_n_354__49_,r_n_354__48_,r_n_354__47_,r_n_354__46_,
  r_n_354__45_,r_n_354__44_,r_n_354__43_,r_n_354__42_,r_n_354__41_,r_n_354__40_,
  r_n_354__39_,r_n_354__38_,r_n_354__37_,r_n_354__36_,r_n_354__35_,r_n_354__34_,
  r_n_354__33_,r_n_354__32_,r_n_354__31_,r_n_354__30_,r_n_354__29_,r_n_354__28_,
  r_n_354__27_,r_n_354__26_,r_n_354__25_,r_n_354__24_,r_n_354__23_,r_n_354__22_,
  r_n_354__21_,r_n_354__20_,r_n_354__19_,r_n_354__18_,r_n_354__17_,r_n_354__16_,r_n_354__15_,
  r_n_354__14_,r_n_354__13_,r_n_354__12_,r_n_354__11_,r_n_354__10_,r_n_354__9_,
  r_n_354__8_,r_n_354__7_,r_n_354__6_,r_n_354__5_,r_n_354__4_,r_n_354__3_,r_n_354__2_,
  r_n_354__1_,r_n_354__0_,r_n_353__63_,r_n_353__62_,r_n_353__61_,r_n_353__60_,
  r_n_353__59_,r_n_353__58_,r_n_353__57_,r_n_353__56_,r_n_353__55_,r_n_353__54_,
  r_n_353__53_,r_n_353__52_,r_n_353__51_,r_n_353__50_,r_n_353__49_,r_n_353__48_,
  r_n_353__47_,r_n_353__46_,r_n_353__45_,r_n_353__44_,r_n_353__43_,r_n_353__42_,
  r_n_353__41_,r_n_353__40_,r_n_353__39_,r_n_353__38_,r_n_353__37_,r_n_353__36_,
  r_n_353__35_,r_n_353__34_,r_n_353__33_,r_n_353__32_,r_n_353__31_,r_n_353__30_,r_n_353__29_,
  r_n_353__28_,r_n_353__27_,r_n_353__26_,r_n_353__25_,r_n_353__24_,r_n_353__23_,
  r_n_353__22_,r_n_353__21_,r_n_353__20_,r_n_353__19_,r_n_353__18_,r_n_353__17_,
  r_n_353__16_,r_n_353__15_,r_n_353__14_,r_n_353__13_,r_n_353__12_,r_n_353__11_,
  r_n_353__10_,r_n_353__9_,r_n_353__8_,r_n_353__7_,r_n_353__6_,r_n_353__5_,r_n_353__4_,
  r_n_353__3_,r_n_353__2_,r_n_353__1_,r_n_353__0_,r_n_368__63_,r_n_368__62_,
  r_n_368__61_,r_n_368__60_,r_n_368__59_,r_n_368__58_,r_n_368__57_,r_n_368__56_,
  r_n_368__55_,r_n_368__54_,r_n_368__53_,r_n_368__52_,r_n_368__51_,r_n_368__50_,
  r_n_368__49_,r_n_368__48_,r_n_368__47_,r_n_368__46_,r_n_368__45_,r_n_368__44_,r_n_368__43_,
  r_n_368__42_,r_n_368__41_,r_n_368__40_,r_n_368__39_,r_n_368__38_,r_n_368__37_,
  r_n_368__36_,r_n_368__35_,r_n_368__34_,r_n_368__33_,r_n_368__32_,r_n_368__31_,
  r_n_368__30_,r_n_368__29_,r_n_368__28_,r_n_368__27_,r_n_368__26_,r_n_368__25_,
  r_n_368__24_,r_n_368__23_,r_n_368__22_,r_n_368__21_,r_n_368__20_,r_n_368__19_,
  r_n_368__18_,r_n_368__17_,r_n_368__16_,r_n_368__15_,r_n_368__14_,r_n_368__13_,
  r_n_368__12_,r_n_368__11_,r_n_368__10_,r_n_368__9_,r_n_368__8_,r_n_368__7_,r_n_368__6_,
  r_n_368__5_,r_n_368__4_,r_n_368__3_,r_n_368__2_,r_n_368__1_,r_n_368__0_,
  r_n_367__63_,r_n_367__62_,r_n_367__61_,r_n_367__60_,r_n_367__59_,r_n_367__58_,r_n_367__57_,
  r_n_367__56_,r_n_367__55_,r_n_367__54_,r_n_367__53_,r_n_367__52_,r_n_367__51_,
  r_n_367__50_,r_n_367__49_,r_n_367__48_,r_n_367__47_,r_n_367__46_,r_n_367__45_,
  r_n_367__44_,r_n_367__43_,r_n_367__42_,r_n_367__41_,r_n_367__40_,r_n_367__39_,
  r_n_367__38_,r_n_367__37_,r_n_367__36_,r_n_367__35_,r_n_367__34_,r_n_367__33_,
  r_n_367__32_,r_n_367__31_,r_n_367__30_,r_n_367__29_,r_n_367__28_,r_n_367__27_,
  r_n_367__26_,r_n_367__25_,r_n_367__24_,r_n_367__23_,r_n_367__22_,r_n_367__21_,r_n_367__20_,
  r_n_367__19_,r_n_367__18_,r_n_367__17_,r_n_367__16_,r_n_367__15_,r_n_367__14_,
  r_n_367__13_,r_n_367__12_,r_n_367__11_,r_n_367__10_,r_n_367__9_,r_n_367__8_,
  r_n_367__7_,r_n_367__6_,r_n_367__5_,r_n_367__4_,r_n_367__3_,r_n_367__2_,r_n_367__1_,
  r_n_367__0_,r_n_366__63_,r_n_366__62_,r_n_366__61_,r_n_366__60_,r_n_366__59_,
  r_n_366__58_,r_n_366__57_,r_n_366__56_,r_n_366__55_,r_n_366__54_,r_n_366__53_,
  r_n_366__52_,r_n_366__51_,r_n_366__50_,r_n_366__49_,r_n_366__48_,r_n_366__47_,
  r_n_366__46_,r_n_366__45_,r_n_366__44_,r_n_366__43_,r_n_366__42_,r_n_366__41_,
  r_n_366__40_,r_n_366__39_,r_n_366__38_,r_n_366__37_,r_n_366__36_,r_n_366__35_,r_n_366__34_,
  r_n_366__33_,r_n_366__32_,r_n_366__31_,r_n_366__30_,r_n_366__29_,r_n_366__28_,
  r_n_366__27_,r_n_366__26_,r_n_366__25_,r_n_366__24_,r_n_366__23_,r_n_366__22_,
  r_n_366__21_,r_n_366__20_,r_n_366__19_,r_n_366__18_,r_n_366__17_,r_n_366__16_,
  r_n_366__15_,r_n_366__14_,r_n_366__13_,r_n_366__12_,r_n_366__11_,r_n_366__10_,
  r_n_366__9_,r_n_366__8_,r_n_366__7_,r_n_366__6_,r_n_366__5_,r_n_366__4_,r_n_366__3_,
  r_n_366__2_,r_n_366__1_,r_n_366__0_,r_n_365__63_,r_n_365__62_,r_n_365__61_,
  r_n_365__60_,r_n_365__59_,r_n_365__58_,r_n_365__57_,r_n_365__56_,r_n_365__55_,
  r_n_365__54_,r_n_365__53_,r_n_365__52_,r_n_365__51_,r_n_365__50_,r_n_365__49_,r_n_365__48_,
  r_n_365__47_,r_n_365__46_,r_n_365__45_,r_n_365__44_,r_n_365__43_,r_n_365__42_,
  r_n_365__41_,r_n_365__40_,r_n_365__39_,r_n_365__38_,r_n_365__37_,r_n_365__36_,
  r_n_365__35_,r_n_365__34_,r_n_365__33_,r_n_365__32_,r_n_365__31_,r_n_365__30_,
  r_n_365__29_,r_n_365__28_,r_n_365__27_,r_n_365__26_,r_n_365__25_,r_n_365__24_,
  r_n_365__23_,r_n_365__22_,r_n_365__21_,r_n_365__20_,r_n_365__19_,r_n_365__18_,
  r_n_365__17_,r_n_365__16_,r_n_365__15_,r_n_365__14_,r_n_365__13_,r_n_365__12_,
  r_n_365__11_,r_n_365__10_,r_n_365__9_,r_n_365__8_,r_n_365__7_,r_n_365__6_,r_n_365__5_,
  r_n_365__4_,r_n_365__3_,r_n_365__2_,r_n_365__1_,r_n_365__0_,r_n_364__63_,r_n_364__62_,
  r_n_364__61_,r_n_364__60_,r_n_364__59_,r_n_364__58_,r_n_364__57_,r_n_364__56_,
  r_n_364__55_,r_n_364__54_,r_n_364__53_,r_n_364__52_,r_n_364__51_,r_n_364__50_,
  r_n_364__49_,r_n_364__48_,r_n_364__47_,r_n_364__46_,r_n_364__45_,r_n_364__44_,
  r_n_364__43_,r_n_364__42_,r_n_364__41_,r_n_364__40_,r_n_364__39_,r_n_364__38_,
  r_n_364__37_,r_n_364__36_,r_n_364__35_,r_n_364__34_,r_n_364__33_,r_n_364__32_,
  r_n_364__31_,r_n_364__30_,r_n_364__29_,r_n_364__28_,r_n_364__27_,r_n_364__26_,
  r_n_364__25_,r_n_364__24_,r_n_364__23_,r_n_364__22_,r_n_364__21_,r_n_364__20_,r_n_364__19_,
  r_n_364__18_,r_n_364__17_,r_n_364__16_,r_n_364__15_,r_n_364__14_,r_n_364__13_,
  r_n_364__12_,r_n_364__11_,r_n_364__10_,r_n_364__9_,r_n_364__8_,r_n_364__7_,
  r_n_364__6_,r_n_364__5_,r_n_364__4_,r_n_364__3_,r_n_364__2_,r_n_364__1_,r_n_364__0_,
  r_n_363__63_,r_n_363__62_,r_n_363__61_,r_n_363__60_,r_n_363__59_,r_n_363__58_,
  r_n_363__57_,r_n_363__56_,r_n_363__55_,r_n_363__54_,r_n_363__53_,r_n_363__52_,
  r_n_363__51_,r_n_363__50_,r_n_363__49_,r_n_363__48_,r_n_363__47_,r_n_363__46_,
  r_n_363__45_,r_n_363__44_,r_n_363__43_,r_n_363__42_,r_n_363__41_,r_n_363__40_,
  r_n_363__39_,r_n_363__38_,r_n_363__37_,r_n_363__36_,r_n_363__35_,r_n_363__34_,r_n_363__33_,
  r_n_363__32_,r_n_363__31_,r_n_363__30_,r_n_363__29_,r_n_363__28_,r_n_363__27_,
  r_n_363__26_,r_n_363__25_,r_n_363__24_,r_n_363__23_,r_n_363__22_,r_n_363__21_,
  r_n_363__20_,r_n_363__19_,r_n_363__18_,r_n_363__17_,r_n_363__16_,r_n_363__15_,
  r_n_363__14_,r_n_363__13_,r_n_363__12_,r_n_363__11_,r_n_363__10_,r_n_363__9_,
  r_n_363__8_,r_n_363__7_,r_n_363__6_,r_n_363__5_,r_n_363__4_,r_n_363__3_,r_n_363__2_,
  r_n_363__1_,r_n_363__0_,r_n_362__63_,r_n_362__62_,r_n_362__61_,r_n_362__60_,
  r_n_362__59_,r_n_362__58_,r_n_362__57_,r_n_362__56_,r_n_362__55_,r_n_362__54_,
  r_n_362__53_,r_n_362__52_,r_n_362__51_,r_n_362__50_,r_n_362__49_,r_n_362__48_,r_n_362__47_,
  r_n_362__46_,r_n_362__45_,r_n_362__44_,r_n_362__43_,r_n_362__42_,r_n_362__41_,
  r_n_362__40_,r_n_362__39_,r_n_362__38_,r_n_362__37_,r_n_362__36_,r_n_362__35_,
  r_n_362__34_,r_n_362__33_,r_n_362__32_,r_n_362__31_,r_n_362__30_,r_n_362__29_,
  r_n_362__28_,r_n_362__27_,r_n_362__26_,r_n_362__25_,r_n_362__24_,r_n_362__23_,
  r_n_362__22_,r_n_362__21_,r_n_362__20_,r_n_362__19_,r_n_362__18_,r_n_362__17_,
  r_n_362__16_,r_n_362__15_,r_n_362__14_,r_n_362__13_,r_n_362__12_,r_n_362__11_,r_n_362__10_,
  r_n_362__9_,r_n_362__8_,r_n_362__7_,r_n_362__6_,r_n_362__5_,r_n_362__4_,
  r_n_362__3_,r_n_362__2_,r_n_362__1_,r_n_362__0_,r_n_361__63_,r_n_361__62_,r_n_361__61_,
  r_n_361__60_,r_n_361__59_,r_n_361__58_,r_n_361__57_,r_n_361__56_,r_n_361__55_,
  r_n_361__54_,r_n_361__53_,r_n_361__52_,r_n_361__51_,r_n_361__50_,r_n_361__49_,
  r_n_361__48_,r_n_361__47_,r_n_361__46_,r_n_361__45_,r_n_361__44_,r_n_361__43_,
  r_n_361__42_,r_n_361__41_,r_n_361__40_,r_n_361__39_,r_n_361__38_,r_n_361__37_,
  r_n_361__36_,r_n_361__35_,r_n_361__34_,r_n_361__33_,r_n_361__32_,r_n_361__31_,
  r_n_361__30_,r_n_361__29_,r_n_361__28_,r_n_361__27_,r_n_361__26_,r_n_361__25_,r_n_361__24_,
  r_n_361__23_,r_n_361__22_,r_n_361__21_,r_n_361__20_,r_n_361__19_,r_n_361__18_,
  r_n_361__17_,r_n_361__16_,r_n_361__15_,r_n_361__14_,r_n_361__13_,r_n_361__12_,
  r_n_361__11_,r_n_361__10_,r_n_361__9_,r_n_361__8_,r_n_361__7_,r_n_361__6_,
  r_n_361__5_,r_n_361__4_,r_n_361__3_,r_n_361__2_,r_n_361__1_,r_n_361__0_,r_n_376__63_,
  r_n_376__62_,r_n_376__61_,r_n_376__60_,r_n_376__59_,r_n_376__58_,r_n_376__57_,
  r_n_376__56_,r_n_376__55_,r_n_376__54_,r_n_376__53_,r_n_376__52_,r_n_376__51_,
  r_n_376__50_,r_n_376__49_,r_n_376__48_,r_n_376__47_,r_n_376__46_,r_n_376__45_,
  r_n_376__44_,r_n_376__43_,r_n_376__42_,r_n_376__41_,r_n_376__40_,r_n_376__39_,r_n_376__38_,
  r_n_376__37_,r_n_376__36_,r_n_376__35_,r_n_376__34_,r_n_376__33_,r_n_376__32_,
  r_n_376__31_,r_n_376__30_,r_n_376__29_,r_n_376__28_,r_n_376__27_,r_n_376__26_,
  r_n_376__25_,r_n_376__24_,r_n_376__23_,r_n_376__22_,r_n_376__21_,r_n_376__20_,
  r_n_376__19_,r_n_376__18_,r_n_376__17_,r_n_376__16_,r_n_376__15_,r_n_376__14_,
  r_n_376__13_,r_n_376__12_,r_n_376__11_,r_n_376__10_,r_n_376__9_,r_n_376__8_,r_n_376__7_,
  r_n_376__6_,r_n_376__5_,r_n_376__4_,r_n_376__3_,r_n_376__2_,r_n_376__1_,
  r_n_376__0_,r_n_375__63_,r_n_375__62_,r_n_375__61_,r_n_375__60_,r_n_375__59_,
  r_n_375__58_,r_n_375__57_,r_n_375__56_,r_n_375__55_,r_n_375__54_,r_n_375__53_,r_n_375__52_,
  r_n_375__51_,r_n_375__50_,r_n_375__49_,r_n_375__48_,r_n_375__47_,r_n_375__46_,
  r_n_375__45_,r_n_375__44_,r_n_375__43_,r_n_375__42_,r_n_375__41_,r_n_375__40_,
  r_n_375__39_,r_n_375__38_,r_n_375__37_,r_n_375__36_,r_n_375__35_,r_n_375__34_,
  r_n_375__33_,r_n_375__32_,r_n_375__31_,r_n_375__30_,r_n_375__29_,r_n_375__28_,
  r_n_375__27_,r_n_375__26_,r_n_375__25_,r_n_375__24_,r_n_375__23_,r_n_375__22_,
  r_n_375__21_,r_n_375__20_,r_n_375__19_,r_n_375__18_,r_n_375__17_,r_n_375__16_,
  r_n_375__15_,r_n_375__14_,r_n_375__13_,r_n_375__12_,r_n_375__11_,r_n_375__10_,r_n_375__9_,
  r_n_375__8_,r_n_375__7_,r_n_375__6_,r_n_375__5_,r_n_375__4_,r_n_375__3_,
  r_n_375__2_,r_n_375__1_,r_n_375__0_,r_n_374__63_,r_n_374__62_,r_n_374__61_,r_n_374__60_,
  r_n_374__59_,r_n_374__58_,r_n_374__57_,r_n_374__56_,r_n_374__55_,r_n_374__54_,
  r_n_374__53_,r_n_374__52_,r_n_374__51_,r_n_374__50_,r_n_374__49_,r_n_374__48_,
  r_n_374__47_,r_n_374__46_,r_n_374__45_,r_n_374__44_,r_n_374__43_,r_n_374__42_,
  r_n_374__41_,r_n_374__40_,r_n_374__39_,r_n_374__38_,r_n_374__37_,r_n_374__36_,
  r_n_374__35_,r_n_374__34_,r_n_374__33_,r_n_374__32_,r_n_374__31_,r_n_374__30_,
  r_n_374__29_,r_n_374__28_,r_n_374__27_,r_n_374__26_,r_n_374__25_,r_n_374__24_,r_n_374__23_,
  r_n_374__22_,r_n_374__21_,r_n_374__20_,r_n_374__19_,r_n_374__18_,r_n_374__17_,
  r_n_374__16_,r_n_374__15_,r_n_374__14_,r_n_374__13_,r_n_374__12_,r_n_374__11_,
  r_n_374__10_,r_n_374__9_,r_n_374__8_,r_n_374__7_,r_n_374__6_,r_n_374__5_,r_n_374__4_,
  r_n_374__3_,r_n_374__2_,r_n_374__1_,r_n_374__0_,r_n_373__63_,r_n_373__62_,
  r_n_373__61_,r_n_373__60_,r_n_373__59_,r_n_373__58_,r_n_373__57_,r_n_373__56_,
  r_n_373__55_,r_n_373__54_,r_n_373__53_,r_n_373__52_,r_n_373__51_,r_n_373__50_,
  r_n_373__49_,r_n_373__48_,r_n_373__47_,r_n_373__46_,r_n_373__45_,r_n_373__44_,
  r_n_373__43_,r_n_373__42_,r_n_373__41_,r_n_373__40_,r_n_373__39_,r_n_373__38_,r_n_373__37_,
  r_n_373__36_,r_n_373__35_,r_n_373__34_,r_n_373__33_,r_n_373__32_,r_n_373__31_,
  r_n_373__30_,r_n_373__29_,r_n_373__28_,r_n_373__27_,r_n_373__26_,r_n_373__25_,
  r_n_373__24_,r_n_373__23_,r_n_373__22_,r_n_373__21_,r_n_373__20_,r_n_373__19_,
  r_n_373__18_,r_n_373__17_,r_n_373__16_,r_n_373__15_,r_n_373__14_,r_n_373__13_,
  r_n_373__12_,r_n_373__11_,r_n_373__10_,r_n_373__9_,r_n_373__8_,r_n_373__7_,r_n_373__6_,
  r_n_373__5_,r_n_373__4_,r_n_373__3_,r_n_373__2_,r_n_373__1_,r_n_373__0_,
  r_n_372__63_,r_n_372__62_,r_n_372__61_,r_n_372__60_,r_n_372__59_,r_n_372__58_,
  r_n_372__57_,r_n_372__56_,r_n_372__55_,r_n_372__54_,r_n_372__53_,r_n_372__52_,r_n_372__51_,
  r_n_372__50_,r_n_372__49_,r_n_372__48_,r_n_372__47_,r_n_372__46_,r_n_372__45_,
  r_n_372__44_,r_n_372__43_,r_n_372__42_,r_n_372__41_,r_n_372__40_,r_n_372__39_,
  r_n_372__38_,r_n_372__37_,r_n_372__36_,r_n_372__35_,r_n_372__34_,r_n_372__33_,
  r_n_372__32_,r_n_372__31_,r_n_372__30_,r_n_372__29_,r_n_372__28_,r_n_372__27_,
  r_n_372__26_,r_n_372__25_,r_n_372__24_,r_n_372__23_,r_n_372__22_,r_n_372__21_,
  r_n_372__20_,r_n_372__19_,r_n_372__18_,r_n_372__17_,r_n_372__16_,r_n_372__15_,r_n_372__14_,
  r_n_372__13_,r_n_372__12_,r_n_372__11_,r_n_372__10_,r_n_372__9_,r_n_372__8_,
  r_n_372__7_,r_n_372__6_,r_n_372__5_,r_n_372__4_,r_n_372__3_,r_n_372__2_,r_n_372__1_,
  r_n_372__0_,r_n_371__63_,r_n_371__62_,r_n_371__61_,r_n_371__60_,r_n_371__59_,
  r_n_371__58_,r_n_371__57_,r_n_371__56_,r_n_371__55_,r_n_371__54_,r_n_371__53_,
  r_n_371__52_,r_n_371__51_,r_n_371__50_,r_n_371__49_,r_n_371__48_,r_n_371__47_,
  r_n_371__46_,r_n_371__45_,r_n_371__44_,r_n_371__43_,r_n_371__42_,r_n_371__41_,
  r_n_371__40_,r_n_371__39_,r_n_371__38_,r_n_371__37_,r_n_371__36_,r_n_371__35_,
  r_n_371__34_,r_n_371__33_,r_n_371__32_,r_n_371__31_,r_n_371__30_,r_n_371__29_,r_n_371__28_,
  r_n_371__27_,r_n_371__26_,r_n_371__25_,r_n_371__24_,r_n_371__23_,r_n_371__22_,
  r_n_371__21_,r_n_371__20_,r_n_371__19_,r_n_371__18_,r_n_371__17_,r_n_371__16_,
  r_n_371__15_,r_n_371__14_,r_n_371__13_,r_n_371__12_,r_n_371__11_,r_n_371__10_,
  r_n_371__9_,r_n_371__8_,r_n_371__7_,r_n_371__6_,r_n_371__5_,r_n_371__4_,r_n_371__3_,
  r_n_371__2_,r_n_371__1_,r_n_371__0_,r_n_370__63_,r_n_370__62_,r_n_370__61_,
  r_n_370__60_,r_n_370__59_,r_n_370__58_,r_n_370__57_,r_n_370__56_,r_n_370__55_,
  r_n_370__54_,r_n_370__53_,r_n_370__52_,r_n_370__51_,r_n_370__50_,r_n_370__49_,
  r_n_370__48_,r_n_370__47_,r_n_370__46_,r_n_370__45_,r_n_370__44_,r_n_370__43_,r_n_370__42_,
  r_n_370__41_,r_n_370__40_,r_n_370__39_,r_n_370__38_,r_n_370__37_,r_n_370__36_,
  r_n_370__35_,r_n_370__34_,r_n_370__33_,r_n_370__32_,r_n_370__31_,r_n_370__30_,
  r_n_370__29_,r_n_370__28_,r_n_370__27_,r_n_370__26_,r_n_370__25_,r_n_370__24_,
  r_n_370__23_,r_n_370__22_,r_n_370__21_,r_n_370__20_,r_n_370__19_,r_n_370__18_,
  r_n_370__17_,r_n_370__16_,r_n_370__15_,r_n_370__14_,r_n_370__13_,r_n_370__12_,
  r_n_370__11_,r_n_370__10_,r_n_370__9_,r_n_370__8_,r_n_370__7_,r_n_370__6_,r_n_370__5_,
  r_n_370__4_,r_n_370__3_,r_n_370__2_,r_n_370__1_,r_n_370__0_,r_n_369__63_,
  r_n_369__62_,r_n_369__61_,r_n_369__60_,r_n_369__59_,r_n_369__58_,r_n_369__57_,r_n_369__56_,
  r_n_369__55_,r_n_369__54_,r_n_369__53_,r_n_369__52_,r_n_369__51_,r_n_369__50_,
  r_n_369__49_,r_n_369__48_,r_n_369__47_,r_n_369__46_,r_n_369__45_,r_n_369__44_,
  r_n_369__43_,r_n_369__42_,r_n_369__41_,r_n_369__40_,r_n_369__39_,r_n_369__38_,
  r_n_369__37_,r_n_369__36_,r_n_369__35_,r_n_369__34_,r_n_369__33_,r_n_369__32_,
  r_n_369__31_,r_n_369__30_,r_n_369__29_,r_n_369__28_,r_n_369__27_,r_n_369__26_,
  r_n_369__25_,r_n_369__24_,r_n_369__23_,r_n_369__22_,r_n_369__21_,r_n_369__20_,
  r_n_369__19_,r_n_369__18_,r_n_369__17_,r_n_369__16_,r_n_369__15_,r_n_369__14_,r_n_369__13_,
  r_n_369__12_,r_n_369__11_,r_n_369__10_,r_n_369__9_,r_n_369__8_,r_n_369__7_,
  r_n_369__6_,r_n_369__5_,r_n_369__4_,r_n_369__3_,r_n_369__2_,r_n_369__1_,r_n_369__0_,
  r_n_384__63_,r_n_384__62_,r_n_384__61_,r_n_384__60_,r_n_384__59_,r_n_384__58_,
  r_n_384__57_,r_n_384__56_,r_n_384__55_,r_n_384__54_,r_n_384__53_,r_n_384__52_,
  r_n_384__51_,r_n_384__50_,r_n_384__49_,r_n_384__48_,r_n_384__47_,r_n_384__46_,
  r_n_384__45_,r_n_384__44_,r_n_384__43_,r_n_384__42_,r_n_384__41_,r_n_384__40_,
  r_n_384__39_,r_n_384__38_,r_n_384__37_,r_n_384__36_,r_n_384__35_,r_n_384__34_,
  r_n_384__33_,r_n_384__32_,r_n_384__31_,r_n_384__30_,r_n_384__29_,r_n_384__28_,r_n_384__27_,
  r_n_384__26_,r_n_384__25_,r_n_384__24_,r_n_384__23_,r_n_384__22_,r_n_384__21_,
  r_n_384__20_,r_n_384__19_,r_n_384__18_,r_n_384__17_,r_n_384__16_,r_n_384__15_,
  r_n_384__14_,r_n_384__13_,r_n_384__12_,r_n_384__11_,r_n_384__10_,r_n_384__9_,
  r_n_384__8_,r_n_384__7_,r_n_384__6_,r_n_384__5_,r_n_384__4_,r_n_384__3_,r_n_384__2_,
  r_n_384__1_,r_n_384__0_,r_n_383__63_,r_n_383__62_,r_n_383__61_,r_n_383__60_,
  r_n_383__59_,r_n_383__58_,r_n_383__57_,r_n_383__56_,r_n_383__55_,r_n_383__54_,
  r_n_383__53_,r_n_383__52_,r_n_383__51_,r_n_383__50_,r_n_383__49_,r_n_383__48_,
  r_n_383__47_,r_n_383__46_,r_n_383__45_,r_n_383__44_,r_n_383__43_,r_n_383__42_,r_n_383__41_,
  r_n_383__40_,r_n_383__39_,r_n_383__38_,r_n_383__37_,r_n_383__36_,r_n_383__35_,
  r_n_383__34_,r_n_383__33_,r_n_383__32_,r_n_383__31_,r_n_383__30_,r_n_383__29_,
  r_n_383__28_,r_n_383__27_,r_n_383__26_,r_n_383__25_,r_n_383__24_,r_n_383__23_,
  r_n_383__22_,r_n_383__21_,r_n_383__20_,r_n_383__19_,r_n_383__18_,r_n_383__17_,
  r_n_383__16_,r_n_383__15_,r_n_383__14_,r_n_383__13_,r_n_383__12_,r_n_383__11_,
  r_n_383__10_,r_n_383__9_,r_n_383__8_,r_n_383__7_,r_n_383__6_,r_n_383__5_,r_n_383__4_,
  r_n_383__3_,r_n_383__2_,r_n_383__1_,r_n_383__0_,r_n_382__63_,r_n_382__62_,
  r_n_382__61_,r_n_382__60_,r_n_382__59_,r_n_382__58_,r_n_382__57_,r_n_382__56_,r_n_382__55_,
  r_n_382__54_,r_n_382__53_,r_n_382__52_,r_n_382__51_,r_n_382__50_,r_n_382__49_,
  r_n_382__48_,r_n_382__47_,r_n_382__46_,r_n_382__45_,r_n_382__44_,r_n_382__43_,
  r_n_382__42_,r_n_382__41_,r_n_382__40_,r_n_382__39_,r_n_382__38_,r_n_382__37_,
  r_n_382__36_,r_n_382__35_,r_n_382__34_,r_n_382__33_,r_n_382__32_,r_n_382__31_,
  r_n_382__30_,r_n_382__29_,r_n_382__28_,r_n_382__27_,r_n_382__26_,r_n_382__25_,
  r_n_382__24_,r_n_382__23_,r_n_382__22_,r_n_382__21_,r_n_382__20_,r_n_382__19_,r_n_382__18_,
  r_n_382__17_,r_n_382__16_,r_n_382__15_,r_n_382__14_,r_n_382__13_,r_n_382__12_,
  r_n_382__11_,r_n_382__10_,r_n_382__9_,r_n_382__8_,r_n_382__7_,r_n_382__6_,
  r_n_382__5_,r_n_382__4_,r_n_382__3_,r_n_382__2_,r_n_382__1_,r_n_382__0_,r_n_381__63_,
  r_n_381__62_,r_n_381__61_,r_n_381__60_,r_n_381__59_,r_n_381__58_,r_n_381__57_,
  r_n_381__56_,r_n_381__55_,r_n_381__54_,r_n_381__53_,r_n_381__52_,r_n_381__51_,
  r_n_381__50_,r_n_381__49_,r_n_381__48_,r_n_381__47_,r_n_381__46_,r_n_381__45_,
  r_n_381__44_,r_n_381__43_,r_n_381__42_,r_n_381__41_,r_n_381__40_,r_n_381__39_,
  r_n_381__38_,r_n_381__37_,r_n_381__36_,r_n_381__35_,r_n_381__34_,r_n_381__33_,r_n_381__32_,
  r_n_381__31_,r_n_381__30_,r_n_381__29_,r_n_381__28_,r_n_381__27_,r_n_381__26_,
  r_n_381__25_,r_n_381__24_,r_n_381__23_,r_n_381__22_,r_n_381__21_,r_n_381__20_,
  r_n_381__19_,r_n_381__18_,r_n_381__17_,r_n_381__16_,r_n_381__15_,r_n_381__14_,
  r_n_381__13_,r_n_381__12_,r_n_381__11_,r_n_381__10_,r_n_381__9_,r_n_381__8_,
  r_n_381__7_,r_n_381__6_,r_n_381__5_,r_n_381__4_,r_n_381__3_,r_n_381__2_,r_n_381__1_,
  r_n_381__0_,r_n_380__63_,r_n_380__62_,r_n_380__61_,r_n_380__60_,r_n_380__59_,
  r_n_380__58_,r_n_380__57_,r_n_380__56_,r_n_380__55_,r_n_380__54_,r_n_380__53_,
  r_n_380__52_,r_n_380__51_,r_n_380__50_,r_n_380__49_,r_n_380__48_,r_n_380__47_,r_n_380__46_,
  r_n_380__45_,r_n_380__44_,r_n_380__43_,r_n_380__42_,r_n_380__41_,r_n_380__40_,
  r_n_380__39_,r_n_380__38_,r_n_380__37_,r_n_380__36_,r_n_380__35_,r_n_380__34_,
  r_n_380__33_,r_n_380__32_,r_n_380__31_,r_n_380__30_,r_n_380__29_,r_n_380__28_,
  r_n_380__27_,r_n_380__26_,r_n_380__25_,r_n_380__24_,r_n_380__23_,r_n_380__22_,
  r_n_380__21_,r_n_380__20_,r_n_380__19_,r_n_380__18_,r_n_380__17_,r_n_380__16_,
  r_n_380__15_,r_n_380__14_,r_n_380__13_,r_n_380__12_,r_n_380__11_,r_n_380__10_,r_n_380__9_,
  r_n_380__8_,r_n_380__7_,r_n_380__6_,r_n_380__5_,r_n_380__4_,r_n_380__3_,
  r_n_380__2_,r_n_380__1_,r_n_380__0_,r_n_379__63_,r_n_379__62_,r_n_379__61_,r_n_379__60_,
  r_n_379__59_,r_n_379__58_,r_n_379__57_,r_n_379__56_,r_n_379__55_,r_n_379__54_,
  r_n_379__53_,r_n_379__52_,r_n_379__51_,r_n_379__50_,r_n_379__49_,r_n_379__48_,
  r_n_379__47_,r_n_379__46_,r_n_379__45_,r_n_379__44_,r_n_379__43_,r_n_379__42_,
  r_n_379__41_,r_n_379__40_,r_n_379__39_,r_n_379__38_,r_n_379__37_,r_n_379__36_,
  r_n_379__35_,r_n_379__34_,r_n_379__33_,r_n_379__32_,r_n_379__31_,r_n_379__30_,
  r_n_379__29_,r_n_379__28_,r_n_379__27_,r_n_379__26_,r_n_379__25_,r_n_379__24_,
  r_n_379__23_,r_n_379__22_,r_n_379__21_,r_n_379__20_,r_n_379__19_,r_n_379__18_,r_n_379__17_,
  r_n_379__16_,r_n_379__15_,r_n_379__14_,r_n_379__13_,r_n_379__12_,r_n_379__11_,
  r_n_379__10_,r_n_379__9_,r_n_379__8_,r_n_379__7_,r_n_379__6_,r_n_379__5_,
  r_n_379__4_,r_n_379__3_,r_n_379__2_,r_n_379__1_,r_n_379__0_,r_n_378__63_,r_n_378__62_,
  r_n_378__61_,r_n_378__60_,r_n_378__59_,r_n_378__58_,r_n_378__57_,r_n_378__56_,
  r_n_378__55_,r_n_378__54_,r_n_378__53_,r_n_378__52_,r_n_378__51_,r_n_378__50_,
  r_n_378__49_,r_n_378__48_,r_n_378__47_,r_n_378__46_,r_n_378__45_,r_n_378__44_,
  r_n_378__43_,r_n_378__42_,r_n_378__41_,r_n_378__40_,r_n_378__39_,r_n_378__38_,
  r_n_378__37_,r_n_378__36_,r_n_378__35_,r_n_378__34_,r_n_378__33_,r_n_378__32_,r_n_378__31_,
  r_n_378__30_,r_n_378__29_,r_n_378__28_,r_n_378__27_,r_n_378__26_,r_n_378__25_,
  r_n_378__24_,r_n_378__23_,r_n_378__22_,r_n_378__21_,r_n_378__20_,r_n_378__19_,
  r_n_378__18_,r_n_378__17_,r_n_378__16_,r_n_378__15_,r_n_378__14_,r_n_378__13_,
  r_n_378__12_,r_n_378__11_,r_n_378__10_,r_n_378__9_,r_n_378__8_,r_n_378__7_,r_n_378__6_,
  r_n_378__5_,r_n_378__4_,r_n_378__3_,r_n_378__2_,r_n_378__1_,r_n_378__0_,
  r_n_377__63_,r_n_377__62_,r_n_377__61_,r_n_377__60_,r_n_377__59_,r_n_377__58_,
  r_n_377__57_,r_n_377__56_,r_n_377__55_,r_n_377__54_,r_n_377__53_,r_n_377__52_,
  r_n_377__51_,r_n_377__50_,r_n_377__49_,r_n_377__48_,r_n_377__47_,r_n_377__46_,r_n_377__45_,
  r_n_377__44_,r_n_377__43_,r_n_377__42_,r_n_377__41_,r_n_377__40_,r_n_377__39_,
  r_n_377__38_,r_n_377__37_,r_n_377__36_,r_n_377__35_,r_n_377__34_,r_n_377__33_,
  r_n_377__32_,r_n_377__31_,r_n_377__30_,r_n_377__29_,r_n_377__28_,r_n_377__27_,
  r_n_377__26_,r_n_377__25_,r_n_377__24_,r_n_377__23_,r_n_377__22_,r_n_377__21_,
  r_n_377__20_,r_n_377__19_,r_n_377__18_,r_n_377__17_,r_n_377__16_,r_n_377__15_,
  r_n_377__14_,r_n_377__13_,r_n_377__12_,r_n_377__11_,r_n_377__10_,r_n_377__9_,r_n_377__8_,
  r_n_377__7_,r_n_377__6_,r_n_377__5_,r_n_377__4_,r_n_377__3_,r_n_377__2_,
  r_n_377__1_,r_n_377__0_,r_n_392__63_,r_n_392__62_,r_n_392__61_,r_n_392__60_,r_n_392__59_,
  r_n_392__58_,r_n_392__57_,r_n_392__56_,r_n_392__55_,r_n_392__54_,r_n_392__53_,
  r_n_392__52_,r_n_392__51_,r_n_392__50_,r_n_392__49_,r_n_392__48_,r_n_392__47_,
  r_n_392__46_,r_n_392__45_,r_n_392__44_,r_n_392__43_,r_n_392__42_,r_n_392__41_,
  r_n_392__40_,r_n_392__39_,r_n_392__38_,r_n_392__37_,r_n_392__36_,r_n_392__35_,
  r_n_392__34_,r_n_392__33_,r_n_392__32_,r_n_392__31_,r_n_392__30_,r_n_392__29_,
  r_n_392__28_,r_n_392__27_,r_n_392__26_,r_n_392__25_,r_n_392__24_,r_n_392__23_,r_n_392__22_,
  r_n_392__21_,r_n_392__20_,r_n_392__19_,r_n_392__18_,r_n_392__17_,r_n_392__16_,
  r_n_392__15_,r_n_392__14_,r_n_392__13_,r_n_392__12_,r_n_392__11_,r_n_392__10_,
  r_n_392__9_,r_n_392__8_,r_n_392__7_,r_n_392__6_,r_n_392__5_,r_n_392__4_,r_n_392__3_,
  r_n_392__2_,r_n_392__1_,r_n_392__0_,r_n_391__63_,r_n_391__62_,r_n_391__61_,
  r_n_391__60_,r_n_391__59_,r_n_391__58_,r_n_391__57_,r_n_391__56_,r_n_391__55_,
  r_n_391__54_,r_n_391__53_,r_n_391__52_,r_n_391__51_,r_n_391__50_,r_n_391__49_,
  r_n_391__48_,r_n_391__47_,r_n_391__46_,r_n_391__45_,r_n_391__44_,r_n_391__43_,
  r_n_391__42_,r_n_391__41_,r_n_391__40_,r_n_391__39_,r_n_391__38_,r_n_391__37_,r_n_391__36_,
  r_n_391__35_,r_n_391__34_,r_n_391__33_,r_n_391__32_,r_n_391__31_,r_n_391__30_,
  r_n_391__29_,r_n_391__28_,r_n_391__27_,r_n_391__26_,r_n_391__25_,r_n_391__24_,
  r_n_391__23_,r_n_391__22_,r_n_391__21_,r_n_391__20_,r_n_391__19_,r_n_391__18_,
  r_n_391__17_,r_n_391__16_,r_n_391__15_,r_n_391__14_,r_n_391__13_,r_n_391__12_,
  r_n_391__11_,r_n_391__10_,r_n_391__9_,r_n_391__8_,r_n_391__7_,r_n_391__6_,r_n_391__5_,
  r_n_391__4_,r_n_391__3_,r_n_391__2_,r_n_391__1_,r_n_391__0_,r_n_390__63_,
  r_n_390__62_,r_n_390__61_,r_n_390__60_,r_n_390__59_,r_n_390__58_,r_n_390__57_,
  r_n_390__56_,r_n_390__55_,r_n_390__54_,r_n_390__53_,r_n_390__52_,r_n_390__51_,r_n_390__50_,
  r_n_390__49_,r_n_390__48_,r_n_390__47_,r_n_390__46_,r_n_390__45_,r_n_390__44_,
  r_n_390__43_,r_n_390__42_,r_n_390__41_,r_n_390__40_,r_n_390__39_,r_n_390__38_,
  r_n_390__37_,r_n_390__36_,r_n_390__35_,r_n_390__34_,r_n_390__33_,r_n_390__32_,
  r_n_390__31_,r_n_390__30_,r_n_390__29_,r_n_390__28_,r_n_390__27_,r_n_390__26_,
  r_n_390__25_,r_n_390__24_,r_n_390__23_,r_n_390__22_,r_n_390__21_,r_n_390__20_,
  r_n_390__19_,r_n_390__18_,r_n_390__17_,r_n_390__16_,r_n_390__15_,r_n_390__14_,
  r_n_390__13_,r_n_390__12_,r_n_390__11_,r_n_390__10_,r_n_390__9_,r_n_390__8_,r_n_390__7_,
  r_n_390__6_,r_n_390__5_,r_n_390__4_,r_n_390__3_,r_n_390__2_,r_n_390__1_,r_n_390__0_,
  r_n_389__63_,r_n_389__62_,r_n_389__61_,r_n_389__60_,r_n_389__59_,r_n_389__58_,
  r_n_389__57_,r_n_389__56_,r_n_389__55_,r_n_389__54_,r_n_389__53_,r_n_389__52_,
  r_n_389__51_,r_n_389__50_,r_n_389__49_,r_n_389__48_,r_n_389__47_,r_n_389__46_,
  r_n_389__45_,r_n_389__44_,r_n_389__43_,r_n_389__42_,r_n_389__41_,r_n_389__40_,
  r_n_389__39_,r_n_389__38_,r_n_389__37_,r_n_389__36_,r_n_389__35_,r_n_389__34_,
  r_n_389__33_,r_n_389__32_,r_n_389__31_,r_n_389__30_,r_n_389__29_,r_n_389__28_,
  r_n_389__27_,r_n_389__26_,r_n_389__25_,r_n_389__24_,r_n_389__23_,r_n_389__22_,r_n_389__21_,
  r_n_389__20_,r_n_389__19_,r_n_389__18_,r_n_389__17_,r_n_389__16_,r_n_389__15_,
  r_n_389__14_,r_n_389__13_,r_n_389__12_,r_n_389__11_,r_n_389__10_,r_n_389__9_,
  r_n_389__8_,r_n_389__7_,r_n_389__6_,r_n_389__5_,r_n_389__4_,r_n_389__3_,r_n_389__2_,
  r_n_389__1_,r_n_389__0_,r_n_388__63_,r_n_388__62_,r_n_388__61_,r_n_388__60_,
  r_n_388__59_,r_n_388__58_,r_n_388__57_,r_n_388__56_,r_n_388__55_,r_n_388__54_,
  r_n_388__53_,r_n_388__52_,r_n_388__51_,r_n_388__50_,r_n_388__49_,r_n_388__48_,
  r_n_388__47_,r_n_388__46_,r_n_388__45_,r_n_388__44_,r_n_388__43_,r_n_388__42_,
  r_n_388__41_,r_n_388__40_,r_n_388__39_,r_n_388__38_,r_n_388__37_,r_n_388__36_,r_n_388__35_,
  r_n_388__34_,r_n_388__33_,r_n_388__32_,r_n_388__31_,r_n_388__30_,r_n_388__29_,
  r_n_388__28_,r_n_388__27_,r_n_388__26_,r_n_388__25_,r_n_388__24_,r_n_388__23_,
  r_n_388__22_,r_n_388__21_,r_n_388__20_,r_n_388__19_,r_n_388__18_,r_n_388__17_,
  r_n_388__16_,r_n_388__15_,r_n_388__14_,r_n_388__13_,r_n_388__12_,r_n_388__11_,
  r_n_388__10_,r_n_388__9_,r_n_388__8_,r_n_388__7_,r_n_388__6_,r_n_388__5_,r_n_388__4_,
  r_n_388__3_,r_n_388__2_,r_n_388__1_,r_n_388__0_,r_n_387__63_,r_n_387__62_,
  r_n_387__61_,r_n_387__60_,r_n_387__59_,r_n_387__58_,r_n_387__57_,r_n_387__56_,
  r_n_387__55_,r_n_387__54_,r_n_387__53_,r_n_387__52_,r_n_387__51_,r_n_387__50_,r_n_387__49_,
  r_n_387__48_,r_n_387__47_,r_n_387__46_,r_n_387__45_,r_n_387__44_,r_n_387__43_,
  r_n_387__42_,r_n_387__41_,r_n_387__40_,r_n_387__39_,r_n_387__38_,r_n_387__37_,
  r_n_387__36_,r_n_387__35_,r_n_387__34_,r_n_387__33_,r_n_387__32_,r_n_387__31_,
  r_n_387__30_,r_n_387__29_,r_n_387__28_,r_n_387__27_,r_n_387__26_,r_n_387__25_,
  r_n_387__24_,r_n_387__23_,r_n_387__22_,r_n_387__21_,r_n_387__20_,r_n_387__19_,
  r_n_387__18_,r_n_387__17_,r_n_387__16_,r_n_387__15_,r_n_387__14_,r_n_387__13_,r_n_387__12_,
  r_n_387__11_,r_n_387__10_,r_n_387__9_,r_n_387__8_,r_n_387__7_,r_n_387__6_,
  r_n_387__5_,r_n_387__4_,r_n_387__3_,r_n_387__2_,r_n_387__1_,r_n_387__0_,r_n_386__63_,
  r_n_386__62_,r_n_386__61_,r_n_386__60_,r_n_386__59_,r_n_386__58_,r_n_386__57_,
  r_n_386__56_,r_n_386__55_,r_n_386__54_,r_n_386__53_,r_n_386__52_,r_n_386__51_,
  r_n_386__50_,r_n_386__49_,r_n_386__48_,r_n_386__47_,r_n_386__46_,r_n_386__45_,
  r_n_386__44_,r_n_386__43_,r_n_386__42_,r_n_386__41_,r_n_386__40_,r_n_386__39_,
  r_n_386__38_,r_n_386__37_,r_n_386__36_,r_n_386__35_,r_n_386__34_,r_n_386__33_,
  r_n_386__32_,r_n_386__31_,r_n_386__30_,r_n_386__29_,r_n_386__28_,r_n_386__27_,r_n_386__26_,
  r_n_386__25_,r_n_386__24_,r_n_386__23_,r_n_386__22_,r_n_386__21_,r_n_386__20_,
  r_n_386__19_,r_n_386__18_,r_n_386__17_,r_n_386__16_,r_n_386__15_,r_n_386__14_,
  r_n_386__13_,r_n_386__12_,r_n_386__11_,r_n_386__10_,r_n_386__9_,r_n_386__8_,
  r_n_386__7_,r_n_386__6_,r_n_386__5_,r_n_386__4_,r_n_386__3_,r_n_386__2_,r_n_386__1_,
  r_n_386__0_,r_n_385__63_,r_n_385__62_,r_n_385__61_,r_n_385__60_,r_n_385__59_,
  r_n_385__58_,r_n_385__57_,r_n_385__56_,r_n_385__55_,r_n_385__54_,r_n_385__53_,
  r_n_385__52_,r_n_385__51_,r_n_385__50_,r_n_385__49_,r_n_385__48_,r_n_385__47_,
  r_n_385__46_,r_n_385__45_,r_n_385__44_,r_n_385__43_,r_n_385__42_,r_n_385__41_,r_n_385__40_,
  r_n_385__39_,r_n_385__38_,r_n_385__37_,r_n_385__36_,r_n_385__35_,r_n_385__34_,
  r_n_385__33_,r_n_385__32_,r_n_385__31_,r_n_385__30_,r_n_385__29_,r_n_385__28_,
  r_n_385__27_,r_n_385__26_,r_n_385__25_,r_n_385__24_,r_n_385__23_,r_n_385__22_,
  r_n_385__21_,r_n_385__20_,r_n_385__19_,r_n_385__18_,r_n_385__17_,r_n_385__16_,
  r_n_385__15_,r_n_385__14_,r_n_385__13_,r_n_385__12_,r_n_385__11_,r_n_385__10_,
  r_n_385__9_,r_n_385__8_,r_n_385__7_,r_n_385__6_,r_n_385__5_,r_n_385__4_,r_n_385__3_,
  r_n_385__2_,r_n_385__1_,r_n_385__0_,r_n_400__63_,r_n_400__62_,r_n_400__61_,
  r_n_400__60_,r_n_400__59_,r_n_400__58_,r_n_400__57_,r_n_400__56_,r_n_400__55_,r_n_400__54_,
  r_n_400__53_,r_n_400__52_,r_n_400__51_,r_n_400__50_,r_n_400__49_,r_n_400__48_,
  r_n_400__47_,r_n_400__46_,r_n_400__45_,r_n_400__44_,r_n_400__43_,r_n_400__42_,
  r_n_400__41_,r_n_400__40_,r_n_400__39_,r_n_400__38_,r_n_400__37_,r_n_400__36_,
  r_n_400__35_,r_n_400__34_,r_n_400__33_,r_n_400__32_,r_n_400__31_,r_n_400__30_,
  r_n_400__29_,r_n_400__28_,r_n_400__27_,r_n_400__26_,r_n_400__25_,r_n_400__24_,
  r_n_400__23_,r_n_400__22_,r_n_400__21_,r_n_400__20_,r_n_400__19_,r_n_400__18_,
  r_n_400__17_,r_n_400__16_,r_n_400__15_,r_n_400__14_,r_n_400__13_,r_n_400__12_,r_n_400__11_,
  r_n_400__10_,r_n_400__9_,r_n_400__8_,r_n_400__7_,r_n_400__6_,r_n_400__5_,
  r_n_400__4_,r_n_400__3_,r_n_400__2_,r_n_400__1_,r_n_400__0_,r_n_399__63_,r_n_399__62_,
  r_n_399__61_,r_n_399__60_,r_n_399__59_,r_n_399__58_,r_n_399__57_,r_n_399__56_,
  r_n_399__55_,r_n_399__54_,r_n_399__53_,r_n_399__52_,r_n_399__51_,r_n_399__50_,
  r_n_399__49_,r_n_399__48_,r_n_399__47_,r_n_399__46_,r_n_399__45_,r_n_399__44_,
  r_n_399__43_,r_n_399__42_,r_n_399__41_,r_n_399__40_,r_n_399__39_,r_n_399__38_,
  r_n_399__37_,r_n_399__36_,r_n_399__35_,r_n_399__34_,r_n_399__33_,r_n_399__32_,
  r_n_399__31_,r_n_399__30_,r_n_399__29_,r_n_399__28_,r_n_399__27_,r_n_399__26_,r_n_399__25_,
  r_n_399__24_,r_n_399__23_,r_n_399__22_,r_n_399__21_,r_n_399__20_,r_n_399__19_,
  r_n_399__18_,r_n_399__17_,r_n_399__16_,r_n_399__15_,r_n_399__14_,r_n_399__13_,
  r_n_399__12_,r_n_399__11_,r_n_399__10_,r_n_399__9_,r_n_399__8_,r_n_399__7_,
  r_n_399__6_,r_n_399__5_,r_n_399__4_,r_n_399__3_,r_n_399__2_,r_n_399__1_,r_n_399__0_,
  r_n_398__63_,r_n_398__62_,r_n_398__61_,r_n_398__60_,r_n_398__59_,r_n_398__58_,
  r_n_398__57_,r_n_398__56_,r_n_398__55_,r_n_398__54_,r_n_398__53_,r_n_398__52_,
  r_n_398__51_,r_n_398__50_,r_n_398__49_,r_n_398__48_,r_n_398__47_,r_n_398__46_,
  r_n_398__45_,r_n_398__44_,r_n_398__43_,r_n_398__42_,r_n_398__41_,r_n_398__40_,r_n_398__39_,
  r_n_398__38_,r_n_398__37_,r_n_398__36_,r_n_398__35_,r_n_398__34_,r_n_398__33_,
  r_n_398__32_,r_n_398__31_,r_n_398__30_,r_n_398__29_,r_n_398__28_,r_n_398__27_,
  r_n_398__26_,r_n_398__25_,r_n_398__24_,r_n_398__23_,r_n_398__22_,r_n_398__21_,
  r_n_398__20_,r_n_398__19_,r_n_398__18_,r_n_398__17_,r_n_398__16_,r_n_398__15_,
  r_n_398__14_,r_n_398__13_,r_n_398__12_,r_n_398__11_,r_n_398__10_,r_n_398__9_,r_n_398__8_,
  r_n_398__7_,r_n_398__6_,r_n_398__5_,r_n_398__4_,r_n_398__3_,r_n_398__2_,
  r_n_398__1_,r_n_398__0_,r_n_397__63_,r_n_397__62_,r_n_397__61_,r_n_397__60_,
  r_n_397__59_,r_n_397__58_,r_n_397__57_,r_n_397__56_,r_n_397__55_,r_n_397__54_,r_n_397__53_,
  r_n_397__52_,r_n_397__51_,r_n_397__50_,r_n_397__49_,r_n_397__48_,r_n_397__47_,
  r_n_397__46_,r_n_397__45_,r_n_397__44_,r_n_397__43_,r_n_397__42_,r_n_397__41_,
  r_n_397__40_,r_n_397__39_,r_n_397__38_,r_n_397__37_,r_n_397__36_,r_n_397__35_,
  r_n_397__34_,r_n_397__33_,r_n_397__32_,r_n_397__31_,r_n_397__30_,r_n_397__29_,
  r_n_397__28_,r_n_397__27_,r_n_397__26_,r_n_397__25_,r_n_397__24_,r_n_397__23_,
  r_n_397__22_,r_n_397__21_,r_n_397__20_,r_n_397__19_,r_n_397__18_,r_n_397__17_,r_n_397__16_,
  r_n_397__15_,r_n_397__14_,r_n_397__13_,r_n_397__12_,r_n_397__11_,r_n_397__10_,
  r_n_397__9_,r_n_397__8_,r_n_397__7_,r_n_397__6_,r_n_397__5_,r_n_397__4_,
  r_n_397__3_,r_n_397__2_,r_n_397__1_,r_n_397__0_,r_n_396__63_,r_n_396__62_,r_n_396__61_,
  r_n_396__60_,r_n_396__59_,r_n_396__58_,r_n_396__57_,r_n_396__56_,r_n_396__55_,
  r_n_396__54_,r_n_396__53_,r_n_396__52_,r_n_396__51_,r_n_396__50_,r_n_396__49_,
  r_n_396__48_,r_n_396__47_,r_n_396__46_,r_n_396__45_,r_n_396__44_,r_n_396__43_,
  r_n_396__42_,r_n_396__41_,r_n_396__40_,r_n_396__39_,r_n_396__38_,r_n_396__37_,
  r_n_396__36_,r_n_396__35_,r_n_396__34_,r_n_396__33_,r_n_396__32_,r_n_396__31_,r_n_396__30_,
  r_n_396__29_,r_n_396__28_,r_n_396__27_,r_n_396__26_,r_n_396__25_,r_n_396__24_,
  r_n_396__23_,r_n_396__22_,r_n_396__21_,r_n_396__20_,r_n_396__19_,r_n_396__18_,
  r_n_396__17_,r_n_396__16_,r_n_396__15_,r_n_396__14_,r_n_396__13_,r_n_396__12_,
  r_n_396__11_,r_n_396__10_,r_n_396__9_,r_n_396__8_,r_n_396__7_,r_n_396__6_,r_n_396__5_,
  r_n_396__4_,r_n_396__3_,r_n_396__2_,r_n_396__1_,r_n_396__0_,r_n_395__63_,
  r_n_395__62_,r_n_395__61_,r_n_395__60_,r_n_395__59_,r_n_395__58_,r_n_395__57_,
  r_n_395__56_,r_n_395__55_,r_n_395__54_,r_n_395__53_,r_n_395__52_,r_n_395__51_,
  r_n_395__50_,r_n_395__49_,r_n_395__48_,r_n_395__47_,r_n_395__46_,r_n_395__45_,r_n_395__44_,
  r_n_395__43_,r_n_395__42_,r_n_395__41_,r_n_395__40_,r_n_395__39_,r_n_395__38_,
  r_n_395__37_,r_n_395__36_,r_n_395__35_,r_n_395__34_,r_n_395__33_,r_n_395__32_,
  r_n_395__31_,r_n_395__30_,r_n_395__29_,r_n_395__28_,r_n_395__27_,r_n_395__26_,
  r_n_395__25_,r_n_395__24_,r_n_395__23_,r_n_395__22_,r_n_395__21_,r_n_395__20_,
  r_n_395__19_,r_n_395__18_,r_n_395__17_,r_n_395__16_,r_n_395__15_,r_n_395__14_,
  r_n_395__13_,r_n_395__12_,r_n_395__11_,r_n_395__10_,r_n_395__9_,r_n_395__8_,r_n_395__7_,
  r_n_395__6_,r_n_395__5_,r_n_395__4_,r_n_395__3_,r_n_395__2_,r_n_395__1_,
  r_n_395__0_,r_n_394__63_,r_n_394__62_,r_n_394__61_,r_n_394__60_,r_n_394__59_,r_n_394__58_,
  r_n_394__57_,r_n_394__56_,r_n_394__55_,r_n_394__54_,r_n_394__53_,r_n_394__52_,
  r_n_394__51_,r_n_394__50_,r_n_394__49_,r_n_394__48_,r_n_394__47_,r_n_394__46_,
  r_n_394__45_,r_n_394__44_,r_n_394__43_,r_n_394__42_,r_n_394__41_,r_n_394__40_,
  r_n_394__39_,r_n_394__38_,r_n_394__37_,r_n_394__36_,r_n_394__35_,r_n_394__34_,
  r_n_394__33_,r_n_394__32_,r_n_394__31_,r_n_394__30_,r_n_394__29_,r_n_394__28_,
  r_n_394__27_,r_n_394__26_,r_n_394__25_,r_n_394__24_,r_n_394__23_,r_n_394__22_,
  r_n_394__21_,r_n_394__20_,r_n_394__19_,r_n_394__18_,r_n_394__17_,r_n_394__16_,r_n_394__15_,
  r_n_394__14_,r_n_394__13_,r_n_394__12_,r_n_394__11_,r_n_394__10_,r_n_394__9_,
  r_n_394__8_,r_n_394__7_,r_n_394__6_,r_n_394__5_,r_n_394__4_,r_n_394__3_,r_n_394__2_,
  r_n_394__1_,r_n_394__0_,r_n_393__63_,r_n_393__62_,r_n_393__61_,r_n_393__60_,
  r_n_393__59_,r_n_393__58_,r_n_393__57_,r_n_393__56_,r_n_393__55_,r_n_393__54_,
  r_n_393__53_,r_n_393__52_,r_n_393__51_,r_n_393__50_,r_n_393__49_,r_n_393__48_,
  r_n_393__47_,r_n_393__46_,r_n_393__45_,r_n_393__44_,r_n_393__43_,r_n_393__42_,
  r_n_393__41_,r_n_393__40_,r_n_393__39_,r_n_393__38_,r_n_393__37_,r_n_393__36_,
  r_n_393__35_,r_n_393__34_,r_n_393__33_,r_n_393__32_,r_n_393__31_,r_n_393__30_,r_n_393__29_,
  r_n_393__28_,r_n_393__27_,r_n_393__26_,r_n_393__25_,r_n_393__24_,r_n_393__23_,
  r_n_393__22_,r_n_393__21_,r_n_393__20_,r_n_393__19_,r_n_393__18_,r_n_393__17_,
  r_n_393__16_,r_n_393__15_,r_n_393__14_,r_n_393__13_,r_n_393__12_,r_n_393__11_,
  r_n_393__10_,r_n_393__9_,r_n_393__8_,r_n_393__7_,r_n_393__6_,r_n_393__5_,r_n_393__4_,
  r_n_393__3_,r_n_393__2_,r_n_393__1_,r_n_393__0_,r_n_408__63_,r_n_408__62_,
  r_n_408__61_,r_n_408__60_,r_n_408__59_,r_n_408__58_,r_n_408__57_,r_n_408__56_,
  r_n_408__55_,r_n_408__54_,r_n_408__53_,r_n_408__52_,r_n_408__51_,r_n_408__50_,
  r_n_408__49_,r_n_408__48_,r_n_408__47_,r_n_408__46_,r_n_408__45_,r_n_408__44_,r_n_408__43_,
  r_n_408__42_,r_n_408__41_,r_n_408__40_,r_n_408__39_,r_n_408__38_,r_n_408__37_,
  r_n_408__36_,r_n_408__35_,r_n_408__34_,r_n_408__33_,r_n_408__32_,r_n_408__31_,
  r_n_408__30_,r_n_408__29_,r_n_408__28_,r_n_408__27_,r_n_408__26_,r_n_408__25_,
  r_n_408__24_,r_n_408__23_,r_n_408__22_,r_n_408__21_,r_n_408__20_,r_n_408__19_,
  r_n_408__18_,r_n_408__17_,r_n_408__16_,r_n_408__15_,r_n_408__14_,r_n_408__13_,
  r_n_408__12_,r_n_408__11_,r_n_408__10_,r_n_408__9_,r_n_408__8_,r_n_408__7_,r_n_408__6_,
  r_n_408__5_,r_n_408__4_,r_n_408__3_,r_n_408__2_,r_n_408__1_,r_n_408__0_,
  r_n_407__63_,r_n_407__62_,r_n_407__61_,r_n_407__60_,r_n_407__59_,r_n_407__58_,r_n_407__57_,
  r_n_407__56_,r_n_407__55_,r_n_407__54_,r_n_407__53_,r_n_407__52_,r_n_407__51_,
  r_n_407__50_,r_n_407__49_,r_n_407__48_,r_n_407__47_,r_n_407__46_,r_n_407__45_,
  r_n_407__44_,r_n_407__43_,r_n_407__42_,r_n_407__41_,r_n_407__40_,r_n_407__39_,
  r_n_407__38_,r_n_407__37_,r_n_407__36_,r_n_407__35_,r_n_407__34_,r_n_407__33_,
  r_n_407__32_,r_n_407__31_,r_n_407__30_,r_n_407__29_,r_n_407__28_,r_n_407__27_,
  r_n_407__26_,r_n_407__25_,r_n_407__24_,r_n_407__23_,r_n_407__22_,r_n_407__21_,r_n_407__20_,
  r_n_407__19_,r_n_407__18_,r_n_407__17_,r_n_407__16_,r_n_407__15_,r_n_407__14_,
  r_n_407__13_,r_n_407__12_,r_n_407__11_,r_n_407__10_,r_n_407__9_,r_n_407__8_,
  r_n_407__7_,r_n_407__6_,r_n_407__5_,r_n_407__4_,r_n_407__3_,r_n_407__2_,r_n_407__1_,
  r_n_407__0_,r_n_406__63_,r_n_406__62_,r_n_406__61_,r_n_406__60_,r_n_406__59_,
  r_n_406__58_,r_n_406__57_,r_n_406__56_,r_n_406__55_,r_n_406__54_,r_n_406__53_,
  r_n_406__52_,r_n_406__51_,r_n_406__50_,r_n_406__49_,r_n_406__48_,r_n_406__47_,
  r_n_406__46_,r_n_406__45_,r_n_406__44_,r_n_406__43_,r_n_406__42_,r_n_406__41_,
  r_n_406__40_,r_n_406__39_,r_n_406__38_,r_n_406__37_,r_n_406__36_,r_n_406__35_,r_n_406__34_,
  r_n_406__33_,r_n_406__32_,r_n_406__31_,r_n_406__30_,r_n_406__29_,r_n_406__28_,
  r_n_406__27_,r_n_406__26_,r_n_406__25_,r_n_406__24_,r_n_406__23_,r_n_406__22_,
  r_n_406__21_,r_n_406__20_,r_n_406__19_,r_n_406__18_,r_n_406__17_,r_n_406__16_,
  r_n_406__15_,r_n_406__14_,r_n_406__13_,r_n_406__12_,r_n_406__11_,r_n_406__10_,
  r_n_406__9_,r_n_406__8_,r_n_406__7_,r_n_406__6_,r_n_406__5_,r_n_406__4_,r_n_406__3_,
  r_n_406__2_,r_n_406__1_,r_n_406__0_,r_n_405__63_,r_n_405__62_,r_n_405__61_,
  r_n_405__60_,r_n_405__59_,r_n_405__58_,r_n_405__57_,r_n_405__56_,r_n_405__55_,
  r_n_405__54_,r_n_405__53_,r_n_405__52_,r_n_405__51_,r_n_405__50_,r_n_405__49_,r_n_405__48_,
  r_n_405__47_,r_n_405__46_,r_n_405__45_,r_n_405__44_,r_n_405__43_,r_n_405__42_,
  r_n_405__41_,r_n_405__40_,r_n_405__39_,r_n_405__38_,r_n_405__37_,r_n_405__36_,
  r_n_405__35_,r_n_405__34_,r_n_405__33_,r_n_405__32_,r_n_405__31_,r_n_405__30_,
  r_n_405__29_,r_n_405__28_,r_n_405__27_,r_n_405__26_,r_n_405__25_,r_n_405__24_,
  r_n_405__23_,r_n_405__22_,r_n_405__21_,r_n_405__20_,r_n_405__19_,r_n_405__18_,
  r_n_405__17_,r_n_405__16_,r_n_405__15_,r_n_405__14_,r_n_405__13_,r_n_405__12_,
  r_n_405__11_,r_n_405__10_,r_n_405__9_,r_n_405__8_,r_n_405__7_,r_n_405__6_,r_n_405__5_,
  r_n_405__4_,r_n_405__3_,r_n_405__2_,r_n_405__1_,r_n_405__0_,r_n_404__63_,r_n_404__62_,
  r_n_404__61_,r_n_404__60_,r_n_404__59_,r_n_404__58_,r_n_404__57_,r_n_404__56_,
  r_n_404__55_,r_n_404__54_,r_n_404__53_,r_n_404__52_,r_n_404__51_,r_n_404__50_,
  r_n_404__49_,r_n_404__48_,r_n_404__47_,r_n_404__46_,r_n_404__45_,r_n_404__44_,
  r_n_404__43_,r_n_404__42_,r_n_404__41_,r_n_404__40_,r_n_404__39_,r_n_404__38_,
  r_n_404__37_,r_n_404__36_,r_n_404__35_,r_n_404__34_,r_n_404__33_,r_n_404__32_,
  r_n_404__31_,r_n_404__30_,r_n_404__29_,r_n_404__28_,r_n_404__27_,r_n_404__26_,
  r_n_404__25_,r_n_404__24_,r_n_404__23_,r_n_404__22_,r_n_404__21_,r_n_404__20_,r_n_404__19_,
  r_n_404__18_,r_n_404__17_,r_n_404__16_,r_n_404__15_,r_n_404__14_,r_n_404__13_,
  r_n_404__12_,r_n_404__11_,r_n_404__10_,r_n_404__9_,r_n_404__8_,r_n_404__7_,
  r_n_404__6_,r_n_404__5_,r_n_404__4_,r_n_404__3_,r_n_404__2_,r_n_404__1_,r_n_404__0_,
  r_n_403__63_,r_n_403__62_,r_n_403__61_,r_n_403__60_,r_n_403__59_,r_n_403__58_,
  r_n_403__57_,r_n_403__56_,r_n_403__55_,r_n_403__54_,r_n_403__53_,r_n_403__52_,
  r_n_403__51_,r_n_403__50_,r_n_403__49_,r_n_403__48_,r_n_403__47_,r_n_403__46_,
  r_n_403__45_,r_n_403__44_,r_n_403__43_,r_n_403__42_,r_n_403__41_,r_n_403__40_,
  r_n_403__39_,r_n_403__38_,r_n_403__37_,r_n_403__36_,r_n_403__35_,r_n_403__34_,r_n_403__33_,
  r_n_403__32_,r_n_403__31_,r_n_403__30_,r_n_403__29_,r_n_403__28_,r_n_403__27_,
  r_n_403__26_,r_n_403__25_,r_n_403__24_,r_n_403__23_,r_n_403__22_,r_n_403__21_,
  r_n_403__20_,r_n_403__19_,r_n_403__18_,r_n_403__17_,r_n_403__16_,r_n_403__15_,
  r_n_403__14_,r_n_403__13_,r_n_403__12_,r_n_403__11_,r_n_403__10_,r_n_403__9_,
  r_n_403__8_,r_n_403__7_,r_n_403__6_,r_n_403__5_,r_n_403__4_,r_n_403__3_,r_n_403__2_,
  r_n_403__1_,r_n_403__0_,r_n_402__63_,r_n_402__62_,r_n_402__61_,r_n_402__60_,
  r_n_402__59_,r_n_402__58_,r_n_402__57_,r_n_402__56_,r_n_402__55_,r_n_402__54_,
  r_n_402__53_,r_n_402__52_,r_n_402__51_,r_n_402__50_,r_n_402__49_,r_n_402__48_,r_n_402__47_,
  r_n_402__46_,r_n_402__45_,r_n_402__44_,r_n_402__43_,r_n_402__42_,r_n_402__41_,
  r_n_402__40_,r_n_402__39_,r_n_402__38_,r_n_402__37_,r_n_402__36_,r_n_402__35_,
  r_n_402__34_,r_n_402__33_,r_n_402__32_,r_n_402__31_,r_n_402__30_,r_n_402__29_,
  r_n_402__28_,r_n_402__27_,r_n_402__26_,r_n_402__25_,r_n_402__24_,r_n_402__23_,
  r_n_402__22_,r_n_402__21_,r_n_402__20_,r_n_402__19_,r_n_402__18_,r_n_402__17_,
  r_n_402__16_,r_n_402__15_,r_n_402__14_,r_n_402__13_,r_n_402__12_,r_n_402__11_,r_n_402__10_,
  r_n_402__9_,r_n_402__8_,r_n_402__7_,r_n_402__6_,r_n_402__5_,r_n_402__4_,
  r_n_402__3_,r_n_402__2_,r_n_402__1_,r_n_402__0_,r_n_401__63_,r_n_401__62_,r_n_401__61_,
  r_n_401__60_,r_n_401__59_,r_n_401__58_,r_n_401__57_,r_n_401__56_,r_n_401__55_,
  r_n_401__54_,r_n_401__53_,r_n_401__52_,r_n_401__51_,r_n_401__50_,r_n_401__49_,
  r_n_401__48_,r_n_401__47_,r_n_401__46_,r_n_401__45_,r_n_401__44_,r_n_401__43_,
  r_n_401__42_,r_n_401__41_,r_n_401__40_,r_n_401__39_,r_n_401__38_,r_n_401__37_,
  r_n_401__36_,r_n_401__35_,r_n_401__34_,r_n_401__33_,r_n_401__32_,r_n_401__31_,
  r_n_401__30_,r_n_401__29_,r_n_401__28_,r_n_401__27_,r_n_401__26_,r_n_401__25_,r_n_401__24_,
  r_n_401__23_,r_n_401__22_,r_n_401__21_,r_n_401__20_,r_n_401__19_,r_n_401__18_,
  r_n_401__17_,r_n_401__16_,r_n_401__15_,r_n_401__14_,r_n_401__13_,r_n_401__12_,
  r_n_401__11_,r_n_401__10_,r_n_401__9_,r_n_401__8_,r_n_401__7_,r_n_401__6_,
  r_n_401__5_,r_n_401__4_,r_n_401__3_,r_n_401__2_,r_n_401__1_,r_n_401__0_,r_n_416__63_,
  r_n_416__62_,r_n_416__61_,r_n_416__60_,r_n_416__59_,r_n_416__58_,r_n_416__57_,
  r_n_416__56_,r_n_416__55_,r_n_416__54_,r_n_416__53_,r_n_416__52_,r_n_416__51_,
  r_n_416__50_,r_n_416__49_,r_n_416__48_,r_n_416__47_,r_n_416__46_,r_n_416__45_,
  r_n_416__44_,r_n_416__43_,r_n_416__42_,r_n_416__41_,r_n_416__40_,r_n_416__39_,r_n_416__38_,
  r_n_416__37_,r_n_416__36_,r_n_416__35_,r_n_416__34_,r_n_416__33_,r_n_416__32_,
  r_n_416__31_,r_n_416__30_,r_n_416__29_,r_n_416__28_,r_n_416__27_,r_n_416__26_,
  r_n_416__25_,r_n_416__24_,r_n_416__23_,r_n_416__22_,r_n_416__21_,r_n_416__20_,
  r_n_416__19_,r_n_416__18_,r_n_416__17_,r_n_416__16_,r_n_416__15_,r_n_416__14_,
  r_n_416__13_,r_n_416__12_,r_n_416__11_,r_n_416__10_,r_n_416__9_,r_n_416__8_,r_n_416__7_,
  r_n_416__6_,r_n_416__5_,r_n_416__4_,r_n_416__3_,r_n_416__2_,r_n_416__1_,
  r_n_416__0_,r_n_415__63_,r_n_415__62_,r_n_415__61_,r_n_415__60_,r_n_415__59_,
  r_n_415__58_,r_n_415__57_,r_n_415__56_,r_n_415__55_,r_n_415__54_,r_n_415__53_,r_n_415__52_,
  r_n_415__51_,r_n_415__50_,r_n_415__49_,r_n_415__48_,r_n_415__47_,r_n_415__46_,
  r_n_415__45_,r_n_415__44_,r_n_415__43_,r_n_415__42_,r_n_415__41_,r_n_415__40_,
  r_n_415__39_,r_n_415__38_,r_n_415__37_,r_n_415__36_,r_n_415__35_,r_n_415__34_,
  r_n_415__33_,r_n_415__32_,r_n_415__31_,r_n_415__30_,r_n_415__29_,r_n_415__28_,
  r_n_415__27_,r_n_415__26_,r_n_415__25_,r_n_415__24_,r_n_415__23_,r_n_415__22_,
  r_n_415__21_,r_n_415__20_,r_n_415__19_,r_n_415__18_,r_n_415__17_,r_n_415__16_,
  r_n_415__15_,r_n_415__14_,r_n_415__13_,r_n_415__12_,r_n_415__11_,r_n_415__10_,r_n_415__9_,
  r_n_415__8_,r_n_415__7_,r_n_415__6_,r_n_415__5_,r_n_415__4_,r_n_415__3_,
  r_n_415__2_,r_n_415__1_,r_n_415__0_,r_n_414__63_,r_n_414__62_,r_n_414__61_,r_n_414__60_,
  r_n_414__59_,r_n_414__58_,r_n_414__57_,r_n_414__56_,r_n_414__55_,r_n_414__54_,
  r_n_414__53_,r_n_414__52_,r_n_414__51_,r_n_414__50_,r_n_414__49_,r_n_414__48_,
  r_n_414__47_,r_n_414__46_,r_n_414__45_,r_n_414__44_,r_n_414__43_,r_n_414__42_,
  r_n_414__41_,r_n_414__40_,r_n_414__39_,r_n_414__38_,r_n_414__37_,r_n_414__36_,
  r_n_414__35_,r_n_414__34_,r_n_414__33_,r_n_414__32_,r_n_414__31_,r_n_414__30_,
  r_n_414__29_,r_n_414__28_,r_n_414__27_,r_n_414__26_,r_n_414__25_,r_n_414__24_,r_n_414__23_,
  r_n_414__22_,r_n_414__21_,r_n_414__20_,r_n_414__19_,r_n_414__18_,r_n_414__17_,
  r_n_414__16_,r_n_414__15_,r_n_414__14_,r_n_414__13_,r_n_414__12_,r_n_414__11_,
  r_n_414__10_,r_n_414__9_,r_n_414__8_,r_n_414__7_,r_n_414__6_,r_n_414__5_,r_n_414__4_,
  r_n_414__3_,r_n_414__2_,r_n_414__1_,r_n_414__0_,r_n_413__63_,r_n_413__62_,
  r_n_413__61_,r_n_413__60_,r_n_413__59_,r_n_413__58_,r_n_413__57_,r_n_413__56_,
  r_n_413__55_,r_n_413__54_,r_n_413__53_,r_n_413__52_,r_n_413__51_,r_n_413__50_,
  r_n_413__49_,r_n_413__48_,r_n_413__47_,r_n_413__46_,r_n_413__45_,r_n_413__44_,
  r_n_413__43_,r_n_413__42_,r_n_413__41_,r_n_413__40_,r_n_413__39_,r_n_413__38_,r_n_413__37_,
  r_n_413__36_,r_n_413__35_,r_n_413__34_,r_n_413__33_,r_n_413__32_,r_n_413__31_,
  r_n_413__30_,r_n_413__29_,r_n_413__28_,r_n_413__27_,r_n_413__26_,r_n_413__25_,
  r_n_413__24_,r_n_413__23_,r_n_413__22_,r_n_413__21_,r_n_413__20_,r_n_413__19_,
  r_n_413__18_,r_n_413__17_,r_n_413__16_,r_n_413__15_,r_n_413__14_,r_n_413__13_,
  r_n_413__12_,r_n_413__11_,r_n_413__10_,r_n_413__9_,r_n_413__8_,r_n_413__7_,r_n_413__6_,
  r_n_413__5_,r_n_413__4_,r_n_413__3_,r_n_413__2_,r_n_413__1_,r_n_413__0_,
  r_n_412__63_,r_n_412__62_,r_n_412__61_,r_n_412__60_,r_n_412__59_,r_n_412__58_,
  r_n_412__57_,r_n_412__56_,r_n_412__55_,r_n_412__54_,r_n_412__53_,r_n_412__52_,r_n_412__51_,
  r_n_412__50_,r_n_412__49_,r_n_412__48_,r_n_412__47_,r_n_412__46_,r_n_412__45_,
  r_n_412__44_,r_n_412__43_,r_n_412__42_,r_n_412__41_,r_n_412__40_,r_n_412__39_,
  r_n_412__38_,r_n_412__37_,r_n_412__36_,r_n_412__35_,r_n_412__34_,r_n_412__33_,
  r_n_412__32_,r_n_412__31_,r_n_412__30_,r_n_412__29_,r_n_412__28_,r_n_412__27_,
  r_n_412__26_,r_n_412__25_,r_n_412__24_,r_n_412__23_,r_n_412__22_,r_n_412__21_,
  r_n_412__20_,r_n_412__19_,r_n_412__18_,r_n_412__17_,r_n_412__16_,r_n_412__15_,r_n_412__14_,
  r_n_412__13_,r_n_412__12_,r_n_412__11_,r_n_412__10_,r_n_412__9_,r_n_412__8_,
  r_n_412__7_,r_n_412__6_,r_n_412__5_,r_n_412__4_,r_n_412__3_,r_n_412__2_,r_n_412__1_,
  r_n_412__0_,r_n_411__63_,r_n_411__62_,r_n_411__61_,r_n_411__60_,r_n_411__59_,
  r_n_411__58_,r_n_411__57_,r_n_411__56_,r_n_411__55_,r_n_411__54_,r_n_411__53_,
  r_n_411__52_,r_n_411__51_,r_n_411__50_,r_n_411__49_,r_n_411__48_,r_n_411__47_,
  r_n_411__46_,r_n_411__45_,r_n_411__44_,r_n_411__43_,r_n_411__42_,r_n_411__41_,
  r_n_411__40_,r_n_411__39_,r_n_411__38_,r_n_411__37_,r_n_411__36_,r_n_411__35_,
  r_n_411__34_,r_n_411__33_,r_n_411__32_,r_n_411__31_,r_n_411__30_,r_n_411__29_,r_n_411__28_,
  r_n_411__27_,r_n_411__26_,r_n_411__25_,r_n_411__24_,r_n_411__23_,r_n_411__22_,
  r_n_411__21_,r_n_411__20_,r_n_411__19_,r_n_411__18_,r_n_411__17_,r_n_411__16_,
  r_n_411__15_,r_n_411__14_,r_n_411__13_,r_n_411__12_,r_n_411__11_,r_n_411__10_,
  r_n_411__9_,r_n_411__8_,r_n_411__7_,r_n_411__6_,r_n_411__5_,r_n_411__4_,r_n_411__3_,
  r_n_411__2_,r_n_411__1_,r_n_411__0_,r_n_410__63_,r_n_410__62_,r_n_410__61_,
  r_n_410__60_,r_n_410__59_,r_n_410__58_,r_n_410__57_,r_n_410__56_,r_n_410__55_,
  r_n_410__54_,r_n_410__53_,r_n_410__52_,r_n_410__51_,r_n_410__50_,r_n_410__49_,
  r_n_410__48_,r_n_410__47_,r_n_410__46_,r_n_410__45_,r_n_410__44_,r_n_410__43_,r_n_410__42_,
  r_n_410__41_,r_n_410__40_,r_n_410__39_,r_n_410__38_,r_n_410__37_,r_n_410__36_,
  r_n_410__35_,r_n_410__34_,r_n_410__33_,r_n_410__32_,r_n_410__31_,r_n_410__30_,
  r_n_410__29_,r_n_410__28_,r_n_410__27_,r_n_410__26_,r_n_410__25_,r_n_410__24_,
  r_n_410__23_,r_n_410__22_,r_n_410__21_,r_n_410__20_,r_n_410__19_,r_n_410__18_,
  r_n_410__17_,r_n_410__16_,r_n_410__15_,r_n_410__14_,r_n_410__13_,r_n_410__12_,
  r_n_410__11_,r_n_410__10_,r_n_410__9_,r_n_410__8_,r_n_410__7_,r_n_410__6_,r_n_410__5_,
  r_n_410__4_,r_n_410__3_,r_n_410__2_,r_n_410__1_,r_n_410__0_,r_n_409__63_,
  r_n_409__62_,r_n_409__61_,r_n_409__60_,r_n_409__59_,r_n_409__58_,r_n_409__57_,r_n_409__56_,
  r_n_409__55_,r_n_409__54_,r_n_409__53_,r_n_409__52_,r_n_409__51_,r_n_409__50_,
  r_n_409__49_,r_n_409__48_,r_n_409__47_,r_n_409__46_,r_n_409__45_,r_n_409__44_,
  r_n_409__43_,r_n_409__42_,r_n_409__41_,r_n_409__40_,r_n_409__39_,r_n_409__38_,
  r_n_409__37_,r_n_409__36_,r_n_409__35_,r_n_409__34_,r_n_409__33_,r_n_409__32_,
  r_n_409__31_,r_n_409__30_,r_n_409__29_,r_n_409__28_,r_n_409__27_,r_n_409__26_,
  r_n_409__25_,r_n_409__24_,r_n_409__23_,r_n_409__22_,r_n_409__21_,r_n_409__20_,
  r_n_409__19_,r_n_409__18_,r_n_409__17_,r_n_409__16_,r_n_409__15_,r_n_409__14_,r_n_409__13_,
  r_n_409__12_,r_n_409__11_,r_n_409__10_,r_n_409__9_,r_n_409__8_,r_n_409__7_,
  r_n_409__6_,r_n_409__5_,r_n_409__4_,r_n_409__3_,r_n_409__2_,r_n_409__1_,r_n_409__0_,
  r_n_424__63_,r_n_424__62_,r_n_424__61_,r_n_424__60_,r_n_424__59_,r_n_424__58_,
  r_n_424__57_,r_n_424__56_,r_n_424__55_,r_n_424__54_,r_n_424__53_,r_n_424__52_,
  r_n_424__51_,r_n_424__50_,r_n_424__49_,r_n_424__48_,r_n_424__47_,r_n_424__46_,
  r_n_424__45_,r_n_424__44_,r_n_424__43_,r_n_424__42_,r_n_424__41_,r_n_424__40_,
  r_n_424__39_,r_n_424__38_,r_n_424__37_,r_n_424__36_,r_n_424__35_,r_n_424__34_,
  r_n_424__33_,r_n_424__32_,r_n_424__31_,r_n_424__30_,r_n_424__29_,r_n_424__28_,r_n_424__27_,
  r_n_424__26_,r_n_424__25_,r_n_424__24_,r_n_424__23_,r_n_424__22_,r_n_424__21_,
  r_n_424__20_,r_n_424__19_,r_n_424__18_,r_n_424__17_,r_n_424__16_,r_n_424__15_,
  r_n_424__14_,r_n_424__13_,r_n_424__12_,r_n_424__11_,r_n_424__10_,r_n_424__9_,
  r_n_424__8_,r_n_424__7_,r_n_424__6_,r_n_424__5_,r_n_424__4_,r_n_424__3_,r_n_424__2_,
  r_n_424__1_,r_n_424__0_,r_n_423__63_,r_n_423__62_,r_n_423__61_,r_n_423__60_,
  r_n_423__59_,r_n_423__58_,r_n_423__57_,r_n_423__56_,r_n_423__55_,r_n_423__54_,
  r_n_423__53_,r_n_423__52_,r_n_423__51_,r_n_423__50_,r_n_423__49_,r_n_423__48_,
  r_n_423__47_,r_n_423__46_,r_n_423__45_,r_n_423__44_,r_n_423__43_,r_n_423__42_,r_n_423__41_,
  r_n_423__40_,r_n_423__39_,r_n_423__38_,r_n_423__37_,r_n_423__36_,r_n_423__35_,
  r_n_423__34_,r_n_423__33_,r_n_423__32_,r_n_423__31_,r_n_423__30_,r_n_423__29_,
  r_n_423__28_,r_n_423__27_,r_n_423__26_,r_n_423__25_,r_n_423__24_,r_n_423__23_,
  r_n_423__22_,r_n_423__21_,r_n_423__20_,r_n_423__19_,r_n_423__18_,r_n_423__17_,
  r_n_423__16_,r_n_423__15_,r_n_423__14_,r_n_423__13_,r_n_423__12_,r_n_423__11_,
  r_n_423__10_,r_n_423__9_,r_n_423__8_,r_n_423__7_,r_n_423__6_,r_n_423__5_,r_n_423__4_,
  r_n_423__3_,r_n_423__2_,r_n_423__1_,r_n_423__0_,r_n_422__63_,r_n_422__62_,
  r_n_422__61_,r_n_422__60_,r_n_422__59_,r_n_422__58_,r_n_422__57_,r_n_422__56_,r_n_422__55_,
  r_n_422__54_,r_n_422__53_,r_n_422__52_,r_n_422__51_,r_n_422__50_,r_n_422__49_,
  r_n_422__48_,r_n_422__47_,r_n_422__46_,r_n_422__45_,r_n_422__44_,r_n_422__43_,
  r_n_422__42_,r_n_422__41_,r_n_422__40_,r_n_422__39_,r_n_422__38_,r_n_422__37_,
  r_n_422__36_,r_n_422__35_,r_n_422__34_,r_n_422__33_,r_n_422__32_,r_n_422__31_,
  r_n_422__30_,r_n_422__29_,r_n_422__28_,r_n_422__27_,r_n_422__26_,r_n_422__25_,
  r_n_422__24_,r_n_422__23_,r_n_422__22_,r_n_422__21_,r_n_422__20_,r_n_422__19_,r_n_422__18_,
  r_n_422__17_,r_n_422__16_,r_n_422__15_,r_n_422__14_,r_n_422__13_,r_n_422__12_,
  r_n_422__11_,r_n_422__10_,r_n_422__9_,r_n_422__8_,r_n_422__7_,r_n_422__6_,
  r_n_422__5_,r_n_422__4_,r_n_422__3_,r_n_422__2_,r_n_422__1_,r_n_422__0_,r_n_421__63_,
  r_n_421__62_,r_n_421__61_,r_n_421__60_,r_n_421__59_,r_n_421__58_,r_n_421__57_,
  r_n_421__56_,r_n_421__55_,r_n_421__54_,r_n_421__53_,r_n_421__52_,r_n_421__51_,
  r_n_421__50_,r_n_421__49_,r_n_421__48_,r_n_421__47_,r_n_421__46_,r_n_421__45_,
  r_n_421__44_,r_n_421__43_,r_n_421__42_,r_n_421__41_,r_n_421__40_,r_n_421__39_,
  r_n_421__38_,r_n_421__37_,r_n_421__36_,r_n_421__35_,r_n_421__34_,r_n_421__33_,r_n_421__32_,
  r_n_421__31_,r_n_421__30_,r_n_421__29_,r_n_421__28_,r_n_421__27_,r_n_421__26_,
  r_n_421__25_,r_n_421__24_,r_n_421__23_,r_n_421__22_,r_n_421__21_,r_n_421__20_,
  r_n_421__19_,r_n_421__18_,r_n_421__17_,r_n_421__16_,r_n_421__15_,r_n_421__14_,
  r_n_421__13_,r_n_421__12_,r_n_421__11_,r_n_421__10_,r_n_421__9_,r_n_421__8_,
  r_n_421__7_,r_n_421__6_,r_n_421__5_,r_n_421__4_,r_n_421__3_,r_n_421__2_,r_n_421__1_,
  r_n_421__0_,r_n_420__63_,r_n_420__62_,r_n_420__61_,r_n_420__60_,r_n_420__59_,
  r_n_420__58_,r_n_420__57_,r_n_420__56_,r_n_420__55_,r_n_420__54_,r_n_420__53_,
  r_n_420__52_,r_n_420__51_,r_n_420__50_,r_n_420__49_,r_n_420__48_,r_n_420__47_,r_n_420__46_,
  r_n_420__45_,r_n_420__44_,r_n_420__43_,r_n_420__42_,r_n_420__41_,r_n_420__40_,
  r_n_420__39_,r_n_420__38_,r_n_420__37_,r_n_420__36_,r_n_420__35_,r_n_420__34_,
  r_n_420__33_,r_n_420__32_,r_n_420__31_,r_n_420__30_,r_n_420__29_,r_n_420__28_,
  r_n_420__27_,r_n_420__26_,r_n_420__25_,r_n_420__24_,r_n_420__23_,r_n_420__22_,
  r_n_420__21_,r_n_420__20_,r_n_420__19_,r_n_420__18_,r_n_420__17_,r_n_420__16_,
  r_n_420__15_,r_n_420__14_,r_n_420__13_,r_n_420__12_,r_n_420__11_,r_n_420__10_,r_n_420__9_,
  r_n_420__8_,r_n_420__7_,r_n_420__6_,r_n_420__5_,r_n_420__4_,r_n_420__3_,
  r_n_420__2_,r_n_420__1_,r_n_420__0_,r_n_419__63_,r_n_419__62_,r_n_419__61_,r_n_419__60_,
  r_n_419__59_,r_n_419__58_,r_n_419__57_,r_n_419__56_,r_n_419__55_,r_n_419__54_,
  r_n_419__53_,r_n_419__52_,r_n_419__51_,r_n_419__50_,r_n_419__49_,r_n_419__48_,
  r_n_419__47_,r_n_419__46_,r_n_419__45_,r_n_419__44_,r_n_419__43_,r_n_419__42_,
  r_n_419__41_,r_n_419__40_,r_n_419__39_,r_n_419__38_,r_n_419__37_,r_n_419__36_,
  r_n_419__35_,r_n_419__34_,r_n_419__33_,r_n_419__32_,r_n_419__31_,r_n_419__30_,
  r_n_419__29_,r_n_419__28_,r_n_419__27_,r_n_419__26_,r_n_419__25_,r_n_419__24_,
  r_n_419__23_,r_n_419__22_,r_n_419__21_,r_n_419__20_,r_n_419__19_,r_n_419__18_,r_n_419__17_,
  r_n_419__16_,r_n_419__15_,r_n_419__14_,r_n_419__13_,r_n_419__12_,r_n_419__11_,
  r_n_419__10_,r_n_419__9_,r_n_419__8_,r_n_419__7_,r_n_419__6_,r_n_419__5_,
  r_n_419__4_,r_n_419__3_,r_n_419__2_,r_n_419__1_,r_n_419__0_,r_n_418__63_,r_n_418__62_,
  r_n_418__61_,r_n_418__60_,r_n_418__59_,r_n_418__58_,r_n_418__57_,r_n_418__56_,
  r_n_418__55_,r_n_418__54_,r_n_418__53_,r_n_418__52_,r_n_418__51_,r_n_418__50_,
  r_n_418__49_,r_n_418__48_,r_n_418__47_,r_n_418__46_,r_n_418__45_,r_n_418__44_,
  r_n_418__43_,r_n_418__42_,r_n_418__41_,r_n_418__40_,r_n_418__39_,r_n_418__38_,
  r_n_418__37_,r_n_418__36_,r_n_418__35_,r_n_418__34_,r_n_418__33_,r_n_418__32_,r_n_418__31_,
  r_n_418__30_,r_n_418__29_,r_n_418__28_,r_n_418__27_,r_n_418__26_,r_n_418__25_,
  r_n_418__24_,r_n_418__23_,r_n_418__22_,r_n_418__21_,r_n_418__20_,r_n_418__19_,
  r_n_418__18_,r_n_418__17_,r_n_418__16_,r_n_418__15_,r_n_418__14_,r_n_418__13_,
  r_n_418__12_,r_n_418__11_,r_n_418__10_,r_n_418__9_,r_n_418__8_,r_n_418__7_,r_n_418__6_,
  r_n_418__5_,r_n_418__4_,r_n_418__3_,r_n_418__2_,r_n_418__1_,r_n_418__0_,
  r_n_417__63_,r_n_417__62_,r_n_417__61_,r_n_417__60_,r_n_417__59_,r_n_417__58_,
  r_n_417__57_,r_n_417__56_,r_n_417__55_,r_n_417__54_,r_n_417__53_,r_n_417__52_,
  r_n_417__51_,r_n_417__50_,r_n_417__49_,r_n_417__48_,r_n_417__47_,r_n_417__46_,r_n_417__45_,
  r_n_417__44_,r_n_417__43_,r_n_417__42_,r_n_417__41_,r_n_417__40_,r_n_417__39_,
  r_n_417__38_,r_n_417__37_,r_n_417__36_,r_n_417__35_,r_n_417__34_,r_n_417__33_,
  r_n_417__32_,r_n_417__31_,r_n_417__30_,r_n_417__29_,r_n_417__28_,r_n_417__27_,
  r_n_417__26_,r_n_417__25_,r_n_417__24_,r_n_417__23_,r_n_417__22_,r_n_417__21_,
  r_n_417__20_,r_n_417__19_,r_n_417__18_,r_n_417__17_,r_n_417__16_,r_n_417__15_,
  r_n_417__14_,r_n_417__13_,r_n_417__12_,r_n_417__11_,r_n_417__10_,r_n_417__9_,r_n_417__8_,
  r_n_417__7_,r_n_417__6_,r_n_417__5_,r_n_417__4_,r_n_417__3_,r_n_417__2_,
  r_n_417__1_,r_n_417__0_,r_n_432__63_,r_n_432__62_,r_n_432__61_,r_n_432__60_,r_n_432__59_,
  r_n_432__58_,r_n_432__57_,r_n_432__56_,r_n_432__55_,r_n_432__54_,r_n_432__53_,
  r_n_432__52_,r_n_432__51_,r_n_432__50_,r_n_432__49_,r_n_432__48_,r_n_432__47_,
  r_n_432__46_,r_n_432__45_,r_n_432__44_,r_n_432__43_,r_n_432__42_,r_n_432__41_,
  r_n_432__40_,r_n_432__39_,r_n_432__38_,r_n_432__37_,r_n_432__36_,r_n_432__35_,
  r_n_432__34_,r_n_432__33_,r_n_432__32_,r_n_432__31_,r_n_432__30_,r_n_432__29_,
  r_n_432__28_,r_n_432__27_,r_n_432__26_,r_n_432__25_,r_n_432__24_,r_n_432__23_,r_n_432__22_,
  r_n_432__21_,r_n_432__20_,r_n_432__19_,r_n_432__18_,r_n_432__17_,r_n_432__16_,
  r_n_432__15_,r_n_432__14_,r_n_432__13_,r_n_432__12_,r_n_432__11_,r_n_432__10_,
  r_n_432__9_,r_n_432__8_,r_n_432__7_,r_n_432__6_,r_n_432__5_,r_n_432__4_,r_n_432__3_,
  r_n_432__2_,r_n_432__1_,r_n_432__0_,r_n_431__63_,r_n_431__62_,r_n_431__61_,
  r_n_431__60_,r_n_431__59_,r_n_431__58_,r_n_431__57_,r_n_431__56_,r_n_431__55_,
  r_n_431__54_,r_n_431__53_,r_n_431__52_,r_n_431__51_,r_n_431__50_,r_n_431__49_,
  r_n_431__48_,r_n_431__47_,r_n_431__46_,r_n_431__45_,r_n_431__44_,r_n_431__43_,
  r_n_431__42_,r_n_431__41_,r_n_431__40_,r_n_431__39_,r_n_431__38_,r_n_431__37_,r_n_431__36_,
  r_n_431__35_,r_n_431__34_,r_n_431__33_,r_n_431__32_,r_n_431__31_,r_n_431__30_,
  r_n_431__29_,r_n_431__28_,r_n_431__27_,r_n_431__26_,r_n_431__25_,r_n_431__24_,
  r_n_431__23_,r_n_431__22_,r_n_431__21_,r_n_431__20_,r_n_431__19_,r_n_431__18_,
  r_n_431__17_,r_n_431__16_,r_n_431__15_,r_n_431__14_,r_n_431__13_,r_n_431__12_,
  r_n_431__11_,r_n_431__10_,r_n_431__9_,r_n_431__8_,r_n_431__7_,r_n_431__6_,r_n_431__5_,
  r_n_431__4_,r_n_431__3_,r_n_431__2_,r_n_431__1_,r_n_431__0_,r_n_430__63_,
  r_n_430__62_,r_n_430__61_,r_n_430__60_,r_n_430__59_,r_n_430__58_,r_n_430__57_,
  r_n_430__56_,r_n_430__55_,r_n_430__54_,r_n_430__53_,r_n_430__52_,r_n_430__51_,r_n_430__50_,
  r_n_430__49_,r_n_430__48_,r_n_430__47_,r_n_430__46_,r_n_430__45_,r_n_430__44_,
  r_n_430__43_,r_n_430__42_,r_n_430__41_,r_n_430__40_,r_n_430__39_,r_n_430__38_,
  r_n_430__37_,r_n_430__36_,r_n_430__35_,r_n_430__34_,r_n_430__33_,r_n_430__32_,
  r_n_430__31_,r_n_430__30_,r_n_430__29_,r_n_430__28_,r_n_430__27_,r_n_430__26_,
  r_n_430__25_,r_n_430__24_,r_n_430__23_,r_n_430__22_,r_n_430__21_,r_n_430__20_,
  r_n_430__19_,r_n_430__18_,r_n_430__17_,r_n_430__16_,r_n_430__15_,r_n_430__14_,
  r_n_430__13_,r_n_430__12_,r_n_430__11_,r_n_430__10_,r_n_430__9_,r_n_430__8_,r_n_430__7_,
  r_n_430__6_,r_n_430__5_,r_n_430__4_,r_n_430__3_,r_n_430__2_,r_n_430__1_,r_n_430__0_,
  r_n_429__63_,r_n_429__62_,r_n_429__61_,r_n_429__60_,r_n_429__59_,r_n_429__58_,
  r_n_429__57_,r_n_429__56_,r_n_429__55_,r_n_429__54_,r_n_429__53_,r_n_429__52_,
  r_n_429__51_,r_n_429__50_,r_n_429__49_,r_n_429__48_,r_n_429__47_,r_n_429__46_,
  r_n_429__45_,r_n_429__44_,r_n_429__43_,r_n_429__42_,r_n_429__41_,r_n_429__40_,
  r_n_429__39_,r_n_429__38_,r_n_429__37_,r_n_429__36_,r_n_429__35_,r_n_429__34_,
  r_n_429__33_,r_n_429__32_,r_n_429__31_,r_n_429__30_,r_n_429__29_,r_n_429__28_,
  r_n_429__27_,r_n_429__26_,r_n_429__25_,r_n_429__24_,r_n_429__23_,r_n_429__22_,r_n_429__21_,
  r_n_429__20_,r_n_429__19_,r_n_429__18_,r_n_429__17_,r_n_429__16_,r_n_429__15_,
  r_n_429__14_,r_n_429__13_,r_n_429__12_,r_n_429__11_,r_n_429__10_,r_n_429__9_,
  r_n_429__8_,r_n_429__7_,r_n_429__6_,r_n_429__5_,r_n_429__4_,r_n_429__3_,r_n_429__2_,
  r_n_429__1_,r_n_429__0_,r_n_428__63_,r_n_428__62_,r_n_428__61_,r_n_428__60_,
  r_n_428__59_,r_n_428__58_,r_n_428__57_,r_n_428__56_,r_n_428__55_,r_n_428__54_,
  r_n_428__53_,r_n_428__52_,r_n_428__51_,r_n_428__50_,r_n_428__49_,r_n_428__48_,
  r_n_428__47_,r_n_428__46_,r_n_428__45_,r_n_428__44_,r_n_428__43_,r_n_428__42_,
  r_n_428__41_,r_n_428__40_,r_n_428__39_,r_n_428__38_,r_n_428__37_,r_n_428__36_,r_n_428__35_,
  r_n_428__34_,r_n_428__33_,r_n_428__32_,r_n_428__31_,r_n_428__30_,r_n_428__29_,
  r_n_428__28_,r_n_428__27_,r_n_428__26_,r_n_428__25_,r_n_428__24_,r_n_428__23_,
  r_n_428__22_,r_n_428__21_,r_n_428__20_,r_n_428__19_,r_n_428__18_,r_n_428__17_,
  r_n_428__16_,r_n_428__15_,r_n_428__14_,r_n_428__13_,r_n_428__12_,r_n_428__11_,
  r_n_428__10_,r_n_428__9_,r_n_428__8_,r_n_428__7_,r_n_428__6_,r_n_428__5_,r_n_428__4_,
  r_n_428__3_,r_n_428__2_,r_n_428__1_,r_n_428__0_,r_n_427__63_,r_n_427__62_,
  r_n_427__61_,r_n_427__60_,r_n_427__59_,r_n_427__58_,r_n_427__57_,r_n_427__56_,
  r_n_427__55_,r_n_427__54_,r_n_427__53_,r_n_427__52_,r_n_427__51_,r_n_427__50_,r_n_427__49_,
  r_n_427__48_,r_n_427__47_,r_n_427__46_,r_n_427__45_,r_n_427__44_,r_n_427__43_,
  r_n_427__42_,r_n_427__41_,r_n_427__40_,r_n_427__39_,r_n_427__38_,r_n_427__37_,
  r_n_427__36_,r_n_427__35_,r_n_427__34_,r_n_427__33_,r_n_427__32_,r_n_427__31_,
  r_n_427__30_,r_n_427__29_,r_n_427__28_,r_n_427__27_,r_n_427__26_,r_n_427__25_,
  r_n_427__24_,r_n_427__23_,r_n_427__22_,r_n_427__21_,r_n_427__20_,r_n_427__19_,
  r_n_427__18_,r_n_427__17_,r_n_427__16_,r_n_427__15_,r_n_427__14_,r_n_427__13_,r_n_427__12_,
  r_n_427__11_,r_n_427__10_,r_n_427__9_,r_n_427__8_,r_n_427__7_,r_n_427__6_,
  r_n_427__5_,r_n_427__4_,r_n_427__3_,r_n_427__2_,r_n_427__1_,r_n_427__0_,r_n_426__63_,
  r_n_426__62_,r_n_426__61_,r_n_426__60_,r_n_426__59_,r_n_426__58_,r_n_426__57_,
  r_n_426__56_,r_n_426__55_,r_n_426__54_,r_n_426__53_,r_n_426__52_,r_n_426__51_,
  r_n_426__50_,r_n_426__49_,r_n_426__48_,r_n_426__47_,r_n_426__46_,r_n_426__45_,
  r_n_426__44_,r_n_426__43_,r_n_426__42_,r_n_426__41_,r_n_426__40_,r_n_426__39_,
  r_n_426__38_,r_n_426__37_,r_n_426__36_,r_n_426__35_,r_n_426__34_,r_n_426__33_,
  r_n_426__32_,r_n_426__31_,r_n_426__30_,r_n_426__29_,r_n_426__28_,r_n_426__27_,r_n_426__26_,
  r_n_426__25_,r_n_426__24_,r_n_426__23_,r_n_426__22_,r_n_426__21_,r_n_426__20_,
  r_n_426__19_,r_n_426__18_,r_n_426__17_,r_n_426__16_,r_n_426__15_,r_n_426__14_,
  r_n_426__13_,r_n_426__12_,r_n_426__11_,r_n_426__10_,r_n_426__9_,r_n_426__8_,
  r_n_426__7_,r_n_426__6_,r_n_426__5_,r_n_426__4_,r_n_426__3_,r_n_426__2_,r_n_426__1_,
  r_n_426__0_,r_n_425__63_,r_n_425__62_,r_n_425__61_,r_n_425__60_,r_n_425__59_,
  r_n_425__58_,r_n_425__57_,r_n_425__56_,r_n_425__55_,r_n_425__54_,r_n_425__53_,
  r_n_425__52_,r_n_425__51_,r_n_425__50_,r_n_425__49_,r_n_425__48_,r_n_425__47_,
  r_n_425__46_,r_n_425__45_,r_n_425__44_,r_n_425__43_,r_n_425__42_,r_n_425__41_,r_n_425__40_,
  r_n_425__39_,r_n_425__38_,r_n_425__37_,r_n_425__36_,r_n_425__35_,r_n_425__34_,
  r_n_425__33_,r_n_425__32_,r_n_425__31_,r_n_425__30_,r_n_425__29_,r_n_425__28_,
  r_n_425__27_,r_n_425__26_,r_n_425__25_,r_n_425__24_,r_n_425__23_,r_n_425__22_,
  r_n_425__21_,r_n_425__20_,r_n_425__19_,r_n_425__18_,r_n_425__17_,r_n_425__16_,
  r_n_425__15_,r_n_425__14_,r_n_425__13_,r_n_425__12_,r_n_425__11_,r_n_425__10_,
  r_n_425__9_,r_n_425__8_,r_n_425__7_,r_n_425__6_,r_n_425__5_,r_n_425__4_,r_n_425__3_,
  r_n_425__2_,r_n_425__1_,r_n_425__0_,r_n_440__63_,r_n_440__62_,r_n_440__61_,
  r_n_440__60_,r_n_440__59_,r_n_440__58_,r_n_440__57_,r_n_440__56_,r_n_440__55_,r_n_440__54_,
  r_n_440__53_,r_n_440__52_,r_n_440__51_,r_n_440__50_,r_n_440__49_,r_n_440__48_,
  r_n_440__47_,r_n_440__46_,r_n_440__45_,r_n_440__44_,r_n_440__43_,r_n_440__42_,
  r_n_440__41_,r_n_440__40_,r_n_440__39_,r_n_440__38_,r_n_440__37_,r_n_440__36_,
  r_n_440__35_,r_n_440__34_,r_n_440__33_,r_n_440__32_,r_n_440__31_,r_n_440__30_,
  r_n_440__29_,r_n_440__28_,r_n_440__27_,r_n_440__26_,r_n_440__25_,r_n_440__24_,
  r_n_440__23_,r_n_440__22_,r_n_440__21_,r_n_440__20_,r_n_440__19_,r_n_440__18_,
  r_n_440__17_,r_n_440__16_,r_n_440__15_,r_n_440__14_,r_n_440__13_,r_n_440__12_,r_n_440__11_,
  r_n_440__10_,r_n_440__9_,r_n_440__8_,r_n_440__7_,r_n_440__6_,r_n_440__5_,
  r_n_440__4_,r_n_440__3_,r_n_440__2_,r_n_440__1_,r_n_440__0_,r_n_439__63_,r_n_439__62_,
  r_n_439__61_,r_n_439__60_,r_n_439__59_,r_n_439__58_,r_n_439__57_,r_n_439__56_,
  r_n_439__55_,r_n_439__54_,r_n_439__53_,r_n_439__52_,r_n_439__51_,r_n_439__50_,
  r_n_439__49_,r_n_439__48_,r_n_439__47_,r_n_439__46_,r_n_439__45_,r_n_439__44_,
  r_n_439__43_,r_n_439__42_,r_n_439__41_,r_n_439__40_,r_n_439__39_,r_n_439__38_,
  r_n_439__37_,r_n_439__36_,r_n_439__35_,r_n_439__34_,r_n_439__33_,r_n_439__32_,
  r_n_439__31_,r_n_439__30_,r_n_439__29_,r_n_439__28_,r_n_439__27_,r_n_439__26_,r_n_439__25_,
  r_n_439__24_,r_n_439__23_,r_n_439__22_,r_n_439__21_,r_n_439__20_,r_n_439__19_,
  r_n_439__18_,r_n_439__17_,r_n_439__16_,r_n_439__15_,r_n_439__14_,r_n_439__13_,
  r_n_439__12_,r_n_439__11_,r_n_439__10_,r_n_439__9_,r_n_439__8_,r_n_439__7_,
  r_n_439__6_,r_n_439__5_,r_n_439__4_,r_n_439__3_,r_n_439__2_,r_n_439__1_,r_n_439__0_,
  r_n_438__63_,r_n_438__62_,r_n_438__61_,r_n_438__60_,r_n_438__59_,r_n_438__58_,
  r_n_438__57_,r_n_438__56_,r_n_438__55_,r_n_438__54_,r_n_438__53_,r_n_438__52_,
  r_n_438__51_,r_n_438__50_,r_n_438__49_,r_n_438__48_,r_n_438__47_,r_n_438__46_,
  r_n_438__45_,r_n_438__44_,r_n_438__43_,r_n_438__42_,r_n_438__41_,r_n_438__40_,r_n_438__39_,
  r_n_438__38_,r_n_438__37_,r_n_438__36_,r_n_438__35_,r_n_438__34_,r_n_438__33_,
  r_n_438__32_,r_n_438__31_,r_n_438__30_,r_n_438__29_,r_n_438__28_,r_n_438__27_,
  r_n_438__26_,r_n_438__25_,r_n_438__24_,r_n_438__23_,r_n_438__22_,r_n_438__21_,
  r_n_438__20_,r_n_438__19_,r_n_438__18_,r_n_438__17_,r_n_438__16_,r_n_438__15_,
  r_n_438__14_,r_n_438__13_,r_n_438__12_,r_n_438__11_,r_n_438__10_,r_n_438__9_,r_n_438__8_,
  r_n_438__7_,r_n_438__6_,r_n_438__5_,r_n_438__4_,r_n_438__3_,r_n_438__2_,
  r_n_438__1_,r_n_438__0_,r_n_437__63_,r_n_437__62_,r_n_437__61_,r_n_437__60_,
  r_n_437__59_,r_n_437__58_,r_n_437__57_,r_n_437__56_,r_n_437__55_,r_n_437__54_,r_n_437__53_,
  r_n_437__52_,r_n_437__51_,r_n_437__50_,r_n_437__49_,r_n_437__48_,r_n_437__47_,
  r_n_437__46_,r_n_437__45_,r_n_437__44_,r_n_437__43_,r_n_437__42_,r_n_437__41_,
  r_n_437__40_,r_n_437__39_,r_n_437__38_,r_n_437__37_,r_n_437__36_,r_n_437__35_,
  r_n_437__34_,r_n_437__33_,r_n_437__32_,r_n_437__31_,r_n_437__30_,r_n_437__29_,
  r_n_437__28_,r_n_437__27_,r_n_437__26_,r_n_437__25_,r_n_437__24_,r_n_437__23_,
  r_n_437__22_,r_n_437__21_,r_n_437__20_,r_n_437__19_,r_n_437__18_,r_n_437__17_,r_n_437__16_,
  r_n_437__15_,r_n_437__14_,r_n_437__13_,r_n_437__12_,r_n_437__11_,r_n_437__10_,
  r_n_437__9_,r_n_437__8_,r_n_437__7_,r_n_437__6_,r_n_437__5_,r_n_437__4_,
  r_n_437__3_,r_n_437__2_,r_n_437__1_,r_n_437__0_,r_n_436__63_,r_n_436__62_,r_n_436__61_,
  r_n_436__60_,r_n_436__59_,r_n_436__58_,r_n_436__57_,r_n_436__56_,r_n_436__55_,
  r_n_436__54_,r_n_436__53_,r_n_436__52_,r_n_436__51_,r_n_436__50_,r_n_436__49_,
  r_n_436__48_,r_n_436__47_,r_n_436__46_,r_n_436__45_,r_n_436__44_,r_n_436__43_,
  r_n_436__42_,r_n_436__41_,r_n_436__40_,r_n_436__39_,r_n_436__38_,r_n_436__37_,
  r_n_436__36_,r_n_436__35_,r_n_436__34_,r_n_436__33_,r_n_436__32_,r_n_436__31_,r_n_436__30_,
  r_n_436__29_,r_n_436__28_,r_n_436__27_,r_n_436__26_,r_n_436__25_,r_n_436__24_,
  r_n_436__23_,r_n_436__22_,r_n_436__21_,r_n_436__20_,r_n_436__19_,r_n_436__18_,
  r_n_436__17_,r_n_436__16_,r_n_436__15_,r_n_436__14_,r_n_436__13_,r_n_436__12_,
  r_n_436__11_,r_n_436__10_,r_n_436__9_,r_n_436__8_,r_n_436__7_,r_n_436__6_,r_n_436__5_,
  r_n_436__4_,r_n_436__3_,r_n_436__2_,r_n_436__1_,r_n_436__0_,r_n_435__63_,
  r_n_435__62_,r_n_435__61_,r_n_435__60_,r_n_435__59_,r_n_435__58_,r_n_435__57_,
  r_n_435__56_,r_n_435__55_,r_n_435__54_,r_n_435__53_,r_n_435__52_,r_n_435__51_,
  r_n_435__50_,r_n_435__49_,r_n_435__48_,r_n_435__47_,r_n_435__46_,r_n_435__45_,r_n_435__44_,
  r_n_435__43_,r_n_435__42_,r_n_435__41_,r_n_435__40_,r_n_435__39_,r_n_435__38_,
  r_n_435__37_,r_n_435__36_,r_n_435__35_,r_n_435__34_,r_n_435__33_,r_n_435__32_,
  r_n_435__31_,r_n_435__30_,r_n_435__29_,r_n_435__28_,r_n_435__27_,r_n_435__26_,
  r_n_435__25_,r_n_435__24_,r_n_435__23_,r_n_435__22_,r_n_435__21_,r_n_435__20_,
  r_n_435__19_,r_n_435__18_,r_n_435__17_,r_n_435__16_,r_n_435__15_,r_n_435__14_,
  r_n_435__13_,r_n_435__12_,r_n_435__11_,r_n_435__10_,r_n_435__9_,r_n_435__8_,r_n_435__7_,
  r_n_435__6_,r_n_435__5_,r_n_435__4_,r_n_435__3_,r_n_435__2_,r_n_435__1_,
  r_n_435__0_,r_n_434__63_,r_n_434__62_,r_n_434__61_,r_n_434__60_,r_n_434__59_,r_n_434__58_,
  r_n_434__57_,r_n_434__56_,r_n_434__55_,r_n_434__54_,r_n_434__53_,r_n_434__52_,
  r_n_434__51_,r_n_434__50_,r_n_434__49_,r_n_434__48_,r_n_434__47_,r_n_434__46_,
  r_n_434__45_,r_n_434__44_,r_n_434__43_,r_n_434__42_,r_n_434__41_,r_n_434__40_,
  r_n_434__39_,r_n_434__38_,r_n_434__37_,r_n_434__36_,r_n_434__35_,r_n_434__34_,
  r_n_434__33_,r_n_434__32_,r_n_434__31_,r_n_434__30_,r_n_434__29_,r_n_434__28_,
  r_n_434__27_,r_n_434__26_,r_n_434__25_,r_n_434__24_,r_n_434__23_,r_n_434__22_,
  r_n_434__21_,r_n_434__20_,r_n_434__19_,r_n_434__18_,r_n_434__17_,r_n_434__16_,r_n_434__15_,
  r_n_434__14_,r_n_434__13_,r_n_434__12_,r_n_434__11_,r_n_434__10_,r_n_434__9_,
  r_n_434__8_,r_n_434__7_,r_n_434__6_,r_n_434__5_,r_n_434__4_,r_n_434__3_,r_n_434__2_,
  r_n_434__1_,r_n_434__0_,r_n_433__63_,r_n_433__62_,r_n_433__61_,r_n_433__60_,
  r_n_433__59_,r_n_433__58_,r_n_433__57_,r_n_433__56_,r_n_433__55_,r_n_433__54_,
  r_n_433__53_,r_n_433__52_,r_n_433__51_,r_n_433__50_,r_n_433__49_,r_n_433__48_,
  r_n_433__47_,r_n_433__46_,r_n_433__45_,r_n_433__44_,r_n_433__43_,r_n_433__42_,
  r_n_433__41_,r_n_433__40_,r_n_433__39_,r_n_433__38_,r_n_433__37_,r_n_433__36_,
  r_n_433__35_,r_n_433__34_,r_n_433__33_,r_n_433__32_,r_n_433__31_,r_n_433__30_,r_n_433__29_,
  r_n_433__28_,r_n_433__27_,r_n_433__26_,r_n_433__25_,r_n_433__24_,r_n_433__23_,
  r_n_433__22_,r_n_433__21_,r_n_433__20_,r_n_433__19_,r_n_433__18_,r_n_433__17_,
  r_n_433__16_,r_n_433__15_,r_n_433__14_,r_n_433__13_,r_n_433__12_,r_n_433__11_,
  r_n_433__10_,r_n_433__9_,r_n_433__8_,r_n_433__7_,r_n_433__6_,r_n_433__5_,r_n_433__4_,
  r_n_433__3_,r_n_433__2_,r_n_433__1_,r_n_433__0_,r_n_448__63_,r_n_448__62_,
  r_n_448__61_,r_n_448__60_,r_n_448__59_,r_n_448__58_,r_n_448__57_,r_n_448__56_,
  r_n_448__55_,r_n_448__54_,r_n_448__53_,r_n_448__52_,r_n_448__51_,r_n_448__50_,
  r_n_448__49_,r_n_448__48_,r_n_448__47_,r_n_448__46_,r_n_448__45_,r_n_448__44_,r_n_448__43_,
  r_n_448__42_,r_n_448__41_,r_n_448__40_,r_n_448__39_,r_n_448__38_,r_n_448__37_,
  r_n_448__36_,r_n_448__35_,r_n_448__34_,r_n_448__33_,r_n_448__32_,r_n_448__31_,
  r_n_448__30_,r_n_448__29_,r_n_448__28_,r_n_448__27_,r_n_448__26_,r_n_448__25_,
  r_n_448__24_,r_n_448__23_,r_n_448__22_,r_n_448__21_,r_n_448__20_,r_n_448__19_,
  r_n_448__18_,r_n_448__17_,r_n_448__16_,r_n_448__15_,r_n_448__14_,r_n_448__13_,
  r_n_448__12_,r_n_448__11_,r_n_448__10_,r_n_448__9_,r_n_448__8_,r_n_448__7_,r_n_448__6_,
  r_n_448__5_,r_n_448__4_,r_n_448__3_,r_n_448__2_,r_n_448__1_,r_n_448__0_,
  r_n_447__63_,r_n_447__62_,r_n_447__61_,r_n_447__60_,r_n_447__59_,r_n_447__58_,r_n_447__57_,
  r_n_447__56_,r_n_447__55_,r_n_447__54_,r_n_447__53_,r_n_447__52_,r_n_447__51_,
  r_n_447__50_,r_n_447__49_,r_n_447__48_,r_n_447__47_,r_n_447__46_,r_n_447__45_,
  r_n_447__44_,r_n_447__43_,r_n_447__42_,r_n_447__41_,r_n_447__40_,r_n_447__39_,
  r_n_447__38_,r_n_447__37_,r_n_447__36_,r_n_447__35_,r_n_447__34_,r_n_447__33_,
  r_n_447__32_,r_n_447__31_,r_n_447__30_,r_n_447__29_,r_n_447__28_,r_n_447__27_,
  r_n_447__26_,r_n_447__25_,r_n_447__24_,r_n_447__23_,r_n_447__22_,r_n_447__21_,r_n_447__20_,
  r_n_447__19_,r_n_447__18_,r_n_447__17_,r_n_447__16_,r_n_447__15_,r_n_447__14_,
  r_n_447__13_,r_n_447__12_,r_n_447__11_,r_n_447__10_,r_n_447__9_,r_n_447__8_,
  r_n_447__7_,r_n_447__6_,r_n_447__5_,r_n_447__4_,r_n_447__3_,r_n_447__2_,r_n_447__1_,
  r_n_447__0_,r_n_446__63_,r_n_446__62_,r_n_446__61_,r_n_446__60_,r_n_446__59_,
  r_n_446__58_,r_n_446__57_,r_n_446__56_,r_n_446__55_,r_n_446__54_,r_n_446__53_,
  r_n_446__52_,r_n_446__51_,r_n_446__50_,r_n_446__49_,r_n_446__48_,r_n_446__47_,
  r_n_446__46_,r_n_446__45_,r_n_446__44_,r_n_446__43_,r_n_446__42_,r_n_446__41_,
  r_n_446__40_,r_n_446__39_,r_n_446__38_,r_n_446__37_,r_n_446__36_,r_n_446__35_,r_n_446__34_,
  r_n_446__33_,r_n_446__32_,r_n_446__31_,r_n_446__30_,r_n_446__29_,r_n_446__28_,
  r_n_446__27_,r_n_446__26_,r_n_446__25_,r_n_446__24_,r_n_446__23_,r_n_446__22_,
  r_n_446__21_,r_n_446__20_,r_n_446__19_,r_n_446__18_,r_n_446__17_,r_n_446__16_,
  r_n_446__15_,r_n_446__14_,r_n_446__13_,r_n_446__12_,r_n_446__11_,r_n_446__10_,
  r_n_446__9_,r_n_446__8_,r_n_446__7_,r_n_446__6_,r_n_446__5_,r_n_446__4_,r_n_446__3_,
  r_n_446__2_,r_n_446__1_,r_n_446__0_,r_n_445__63_,r_n_445__62_,r_n_445__61_,
  r_n_445__60_,r_n_445__59_,r_n_445__58_,r_n_445__57_,r_n_445__56_,r_n_445__55_,
  r_n_445__54_,r_n_445__53_,r_n_445__52_,r_n_445__51_,r_n_445__50_,r_n_445__49_,r_n_445__48_,
  r_n_445__47_,r_n_445__46_,r_n_445__45_,r_n_445__44_,r_n_445__43_,r_n_445__42_,
  r_n_445__41_,r_n_445__40_,r_n_445__39_,r_n_445__38_,r_n_445__37_,r_n_445__36_,
  r_n_445__35_,r_n_445__34_,r_n_445__33_,r_n_445__32_,r_n_445__31_,r_n_445__30_,
  r_n_445__29_,r_n_445__28_,r_n_445__27_,r_n_445__26_,r_n_445__25_,r_n_445__24_,
  r_n_445__23_,r_n_445__22_,r_n_445__21_,r_n_445__20_,r_n_445__19_,r_n_445__18_,
  r_n_445__17_,r_n_445__16_,r_n_445__15_,r_n_445__14_,r_n_445__13_,r_n_445__12_,
  r_n_445__11_,r_n_445__10_,r_n_445__9_,r_n_445__8_,r_n_445__7_,r_n_445__6_,r_n_445__5_,
  r_n_445__4_,r_n_445__3_,r_n_445__2_,r_n_445__1_,r_n_445__0_,r_n_444__63_,r_n_444__62_,
  r_n_444__61_,r_n_444__60_,r_n_444__59_,r_n_444__58_,r_n_444__57_,r_n_444__56_,
  r_n_444__55_,r_n_444__54_,r_n_444__53_,r_n_444__52_,r_n_444__51_,r_n_444__50_,
  r_n_444__49_,r_n_444__48_,r_n_444__47_,r_n_444__46_,r_n_444__45_,r_n_444__44_,
  r_n_444__43_,r_n_444__42_,r_n_444__41_,r_n_444__40_,r_n_444__39_,r_n_444__38_,
  r_n_444__37_,r_n_444__36_,r_n_444__35_,r_n_444__34_,r_n_444__33_,r_n_444__32_,
  r_n_444__31_,r_n_444__30_,r_n_444__29_,r_n_444__28_,r_n_444__27_,r_n_444__26_,
  r_n_444__25_,r_n_444__24_,r_n_444__23_,r_n_444__22_,r_n_444__21_,r_n_444__20_,r_n_444__19_,
  r_n_444__18_,r_n_444__17_,r_n_444__16_,r_n_444__15_,r_n_444__14_,r_n_444__13_,
  r_n_444__12_,r_n_444__11_,r_n_444__10_,r_n_444__9_,r_n_444__8_,r_n_444__7_,
  r_n_444__6_,r_n_444__5_,r_n_444__4_,r_n_444__3_,r_n_444__2_,r_n_444__1_,r_n_444__0_,
  r_n_443__63_,r_n_443__62_,r_n_443__61_,r_n_443__60_,r_n_443__59_,r_n_443__58_,
  r_n_443__57_,r_n_443__56_,r_n_443__55_,r_n_443__54_,r_n_443__53_,r_n_443__52_,
  r_n_443__51_,r_n_443__50_,r_n_443__49_,r_n_443__48_,r_n_443__47_,r_n_443__46_,
  r_n_443__45_,r_n_443__44_,r_n_443__43_,r_n_443__42_,r_n_443__41_,r_n_443__40_,
  r_n_443__39_,r_n_443__38_,r_n_443__37_,r_n_443__36_,r_n_443__35_,r_n_443__34_,r_n_443__33_,
  r_n_443__32_,r_n_443__31_,r_n_443__30_,r_n_443__29_,r_n_443__28_,r_n_443__27_,
  r_n_443__26_,r_n_443__25_,r_n_443__24_,r_n_443__23_,r_n_443__22_,r_n_443__21_,
  r_n_443__20_,r_n_443__19_,r_n_443__18_,r_n_443__17_,r_n_443__16_,r_n_443__15_,
  r_n_443__14_,r_n_443__13_,r_n_443__12_,r_n_443__11_,r_n_443__10_,r_n_443__9_,
  r_n_443__8_,r_n_443__7_,r_n_443__6_,r_n_443__5_,r_n_443__4_,r_n_443__3_,r_n_443__2_,
  r_n_443__1_,r_n_443__0_,r_n_442__63_,r_n_442__62_,r_n_442__61_,r_n_442__60_,
  r_n_442__59_,r_n_442__58_,r_n_442__57_,r_n_442__56_,r_n_442__55_,r_n_442__54_,
  r_n_442__53_,r_n_442__52_,r_n_442__51_,r_n_442__50_,r_n_442__49_,r_n_442__48_,r_n_442__47_,
  r_n_442__46_,r_n_442__45_,r_n_442__44_,r_n_442__43_,r_n_442__42_,r_n_442__41_,
  r_n_442__40_,r_n_442__39_,r_n_442__38_,r_n_442__37_,r_n_442__36_,r_n_442__35_,
  r_n_442__34_,r_n_442__33_,r_n_442__32_,r_n_442__31_,r_n_442__30_,r_n_442__29_,
  r_n_442__28_,r_n_442__27_,r_n_442__26_,r_n_442__25_,r_n_442__24_,r_n_442__23_,
  r_n_442__22_,r_n_442__21_,r_n_442__20_,r_n_442__19_,r_n_442__18_,r_n_442__17_,
  r_n_442__16_,r_n_442__15_,r_n_442__14_,r_n_442__13_,r_n_442__12_,r_n_442__11_,r_n_442__10_,
  r_n_442__9_,r_n_442__8_,r_n_442__7_,r_n_442__6_,r_n_442__5_,r_n_442__4_,
  r_n_442__3_,r_n_442__2_,r_n_442__1_,r_n_442__0_,r_n_441__63_,r_n_441__62_,r_n_441__61_,
  r_n_441__60_,r_n_441__59_,r_n_441__58_,r_n_441__57_,r_n_441__56_,r_n_441__55_,
  r_n_441__54_,r_n_441__53_,r_n_441__52_,r_n_441__51_,r_n_441__50_,r_n_441__49_,
  r_n_441__48_,r_n_441__47_,r_n_441__46_,r_n_441__45_,r_n_441__44_,r_n_441__43_,
  r_n_441__42_,r_n_441__41_,r_n_441__40_,r_n_441__39_,r_n_441__38_,r_n_441__37_,
  r_n_441__36_,r_n_441__35_,r_n_441__34_,r_n_441__33_,r_n_441__32_,r_n_441__31_,
  r_n_441__30_,r_n_441__29_,r_n_441__28_,r_n_441__27_,r_n_441__26_,r_n_441__25_,r_n_441__24_,
  r_n_441__23_,r_n_441__22_,r_n_441__21_,r_n_441__20_,r_n_441__19_,r_n_441__18_,
  r_n_441__17_,r_n_441__16_,r_n_441__15_,r_n_441__14_,r_n_441__13_,r_n_441__12_,
  r_n_441__11_,r_n_441__10_,r_n_441__9_,r_n_441__8_,r_n_441__7_,r_n_441__6_,
  r_n_441__5_,r_n_441__4_,r_n_441__3_,r_n_441__2_,r_n_441__1_,r_n_441__0_,r_n_456__63_,
  r_n_456__62_,r_n_456__61_,r_n_456__60_,r_n_456__59_,r_n_456__58_,r_n_456__57_,
  r_n_456__56_,r_n_456__55_,r_n_456__54_,r_n_456__53_,r_n_456__52_,r_n_456__51_,
  r_n_456__50_,r_n_456__49_,r_n_456__48_,r_n_456__47_,r_n_456__46_,r_n_456__45_,
  r_n_456__44_,r_n_456__43_,r_n_456__42_,r_n_456__41_,r_n_456__40_,r_n_456__39_,r_n_456__38_,
  r_n_456__37_,r_n_456__36_,r_n_456__35_,r_n_456__34_,r_n_456__33_,r_n_456__32_,
  r_n_456__31_,r_n_456__30_,r_n_456__29_,r_n_456__28_,r_n_456__27_,r_n_456__26_,
  r_n_456__25_,r_n_456__24_,r_n_456__23_,r_n_456__22_,r_n_456__21_,r_n_456__20_,
  r_n_456__19_,r_n_456__18_,r_n_456__17_,r_n_456__16_,r_n_456__15_,r_n_456__14_,
  r_n_456__13_,r_n_456__12_,r_n_456__11_,r_n_456__10_,r_n_456__9_,r_n_456__8_,r_n_456__7_,
  r_n_456__6_,r_n_456__5_,r_n_456__4_,r_n_456__3_,r_n_456__2_,r_n_456__1_,
  r_n_456__0_,r_n_455__63_,r_n_455__62_,r_n_455__61_,r_n_455__60_,r_n_455__59_,
  r_n_455__58_,r_n_455__57_,r_n_455__56_,r_n_455__55_,r_n_455__54_,r_n_455__53_,r_n_455__52_,
  r_n_455__51_,r_n_455__50_,r_n_455__49_,r_n_455__48_,r_n_455__47_,r_n_455__46_,
  r_n_455__45_,r_n_455__44_,r_n_455__43_,r_n_455__42_,r_n_455__41_,r_n_455__40_,
  r_n_455__39_,r_n_455__38_,r_n_455__37_,r_n_455__36_,r_n_455__35_,r_n_455__34_,
  r_n_455__33_,r_n_455__32_,r_n_455__31_,r_n_455__30_,r_n_455__29_,r_n_455__28_,
  r_n_455__27_,r_n_455__26_,r_n_455__25_,r_n_455__24_,r_n_455__23_,r_n_455__22_,
  r_n_455__21_,r_n_455__20_,r_n_455__19_,r_n_455__18_,r_n_455__17_,r_n_455__16_,
  r_n_455__15_,r_n_455__14_,r_n_455__13_,r_n_455__12_,r_n_455__11_,r_n_455__10_,r_n_455__9_,
  r_n_455__8_,r_n_455__7_,r_n_455__6_,r_n_455__5_,r_n_455__4_,r_n_455__3_,
  r_n_455__2_,r_n_455__1_,r_n_455__0_,r_n_454__63_,r_n_454__62_,r_n_454__61_,r_n_454__60_,
  r_n_454__59_,r_n_454__58_,r_n_454__57_,r_n_454__56_,r_n_454__55_,r_n_454__54_,
  r_n_454__53_,r_n_454__52_,r_n_454__51_,r_n_454__50_,r_n_454__49_,r_n_454__48_,
  r_n_454__47_,r_n_454__46_,r_n_454__45_,r_n_454__44_,r_n_454__43_,r_n_454__42_,
  r_n_454__41_,r_n_454__40_,r_n_454__39_,r_n_454__38_,r_n_454__37_,r_n_454__36_,
  r_n_454__35_,r_n_454__34_,r_n_454__33_,r_n_454__32_,r_n_454__31_,r_n_454__30_,
  r_n_454__29_,r_n_454__28_,r_n_454__27_,r_n_454__26_,r_n_454__25_,r_n_454__24_,r_n_454__23_,
  r_n_454__22_,r_n_454__21_,r_n_454__20_,r_n_454__19_,r_n_454__18_,r_n_454__17_,
  r_n_454__16_,r_n_454__15_,r_n_454__14_,r_n_454__13_,r_n_454__12_,r_n_454__11_,
  r_n_454__10_,r_n_454__9_,r_n_454__8_,r_n_454__7_,r_n_454__6_,r_n_454__5_,r_n_454__4_,
  r_n_454__3_,r_n_454__2_,r_n_454__1_,r_n_454__0_,r_n_453__63_,r_n_453__62_,
  r_n_453__61_,r_n_453__60_,r_n_453__59_,r_n_453__58_,r_n_453__57_,r_n_453__56_,
  r_n_453__55_,r_n_453__54_,r_n_453__53_,r_n_453__52_,r_n_453__51_,r_n_453__50_,
  r_n_453__49_,r_n_453__48_,r_n_453__47_,r_n_453__46_,r_n_453__45_,r_n_453__44_,
  r_n_453__43_,r_n_453__42_,r_n_453__41_,r_n_453__40_,r_n_453__39_,r_n_453__38_,r_n_453__37_,
  r_n_453__36_,r_n_453__35_,r_n_453__34_,r_n_453__33_,r_n_453__32_,r_n_453__31_,
  r_n_453__30_,r_n_453__29_,r_n_453__28_,r_n_453__27_,r_n_453__26_,r_n_453__25_,
  r_n_453__24_,r_n_453__23_,r_n_453__22_,r_n_453__21_,r_n_453__20_,r_n_453__19_,
  r_n_453__18_,r_n_453__17_,r_n_453__16_,r_n_453__15_,r_n_453__14_,r_n_453__13_,
  r_n_453__12_,r_n_453__11_,r_n_453__10_,r_n_453__9_,r_n_453__8_,r_n_453__7_,r_n_453__6_,
  r_n_453__5_,r_n_453__4_,r_n_453__3_,r_n_453__2_,r_n_453__1_,r_n_453__0_,
  r_n_452__63_,r_n_452__62_,r_n_452__61_,r_n_452__60_,r_n_452__59_,r_n_452__58_,
  r_n_452__57_,r_n_452__56_,r_n_452__55_,r_n_452__54_,r_n_452__53_,r_n_452__52_,r_n_452__51_,
  r_n_452__50_,r_n_452__49_,r_n_452__48_,r_n_452__47_,r_n_452__46_,r_n_452__45_,
  r_n_452__44_,r_n_452__43_,r_n_452__42_,r_n_452__41_,r_n_452__40_,r_n_452__39_,
  r_n_452__38_,r_n_452__37_,r_n_452__36_,r_n_452__35_,r_n_452__34_,r_n_452__33_,
  r_n_452__32_,r_n_452__31_,r_n_452__30_,r_n_452__29_,r_n_452__28_,r_n_452__27_,
  r_n_452__26_,r_n_452__25_,r_n_452__24_,r_n_452__23_,r_n_452__22_,r_n_452__21_,
  r_n_452__20_,r_n_452__19_,r_n_452__18_,r_n_452__17_,r_n_452__16_,r_n_452__15_,r_n_452__14_,
  r_n_452__13_,r_n_452__12_,r_n_452__11_,r_n_452__10_,r_n_452__9_,r_n_452__8_,
  r_n_452__7_,r_n_452__6_,r_n_452__5_,r_n_452__4_,r_n_452__3_,r_n_452__2_,r_n_452__1_,
  r_n_452__0_,r_n_451__63_,r_n_451__62_,r_n_451__61_,r_n_451__60_,r_n_451__59_,
  r_n_451__58_,r_n_451__57_,r_n_451__56_,r_n_451__55_,r_n_451__54_,r_n_451__53_,
  r_n_451__52_,r_n_451__51_,r_n_451__50_,r_n_451__49_,r_n_451__48_,r_n_451__47_,
  r_n_451__46_,r_n_451__45_,r_n_451__44_,r_n_451__43_,r_n_451__42_,r_n_451__41_,
  r_n_451__40_,r_n_451__39_,r_n_451__38_,r_n_451__37_,r_n_451__36_,r_n_451__35_,
  r_n_451__34_,r_n_451__33_,r_n_451__32_,r_n_451__31_,r_n_451__30_,r_n_451__29_,r_n_451__28_,
  r_n_451__27_,r_n_451__26_,r_n_451__25_,r_n_451__24_,r_n_451__23_,r_n_451__22_,
  r_n_451__21_,r_n_451__20_,r_n_451__19_,r_n_451__18_,r_n_451__17_,r_n_451__16_,
  r_n_451__15_,r_n_451__14_,r_n_451__13_,r_n_451__12_,r_n_451__11_,r_n_451__10_,
  r_n_451__9_,r_n_451__8_,r_n_451__7_,r_n_451__6_,r_n_451__5_,r_n_451__4_,r_n_451__3_,
  r_n_451__2_,r_n_451__1_,r_n_451__0_,r_n_450__63_,r_n_450__62_,r_n_450__61_,
  r_n_450__60_,r_n_450__59_,r_n_450__58_,r_n_450__57_,r_n_450__56_,r_n_450__55_,
  r_n_450__54_,r_n_450__53_,r_n_450__52_,r_n_450__51_,r_n_450__50_,r_n_450__49_,
  r_n_450__48_,r_n_450__47_,r_n_450__46_,r_n_450__45_,r_n_450__44_,r_n_450__43_,r_n_450__42_,
  r_n_450__41_,r_n_450__40_,r_n_450__39_,r_n_450__38_,r_n_450__37_,r_n_450__36_,
  r_n_450__35_,r_n_450__34_,r_n_450__33_,r_n_450__32_,r_n_450__31_,r_n_450__30_,
  r_n_450__29_,r_n_450__28_,r_n_450__27_,r_n_450__26_,r_n_450__25_,r_n_450__24_,
  r_n_450__23_,r_n_450__22_,r_n_450__21_,r_n_450__20_,r_n_450__19_,r_n_450__18_,
  r_n_450__17_,r_n_450__16_,r_n_450__15_,r_n_450__14_,r_n_450__13_,r_n_450__12_,
  r_n_450__11_,r_n_450__10_,r_n_450__9_,r_n_450__8_,r_n_450__7_,r_n_450__6_,r_n_450__5_,
  r_n_450__4_,r_n_450__3_,r_n_450__2_,r_n_450__1_,r_n_450__0_,r_n_449__63_,
  r_n_449__62_,r_n_449__61_,r_n_449__60_,r_n_449__59_,r_n_449__58_,r_n_449__57_,r_n_449__56_,
  r_n_449__55_,r_n_449__54_,r_n_449__53_,r_n_449__52_,r_n_449__51_,r_n_449__50_,
  r_n_449__49_,r_n_449__48_,r_n_449__47_,r_n_449__46_,r_n_449__45_,r_n_449__44_,
  r_n_449__43_,r_n_449__42_,r_n_449__41_,r_n_449__40_,r_n_449__39_,r_n_449__38_,
  r_n_449__37_,r_n_449__36_,r_n_449__35_,r_n_449__34_,r_n_449__33_,r_n_449__32_,
  r_n_449__31_,r_n_449__30_,r_n_449__29_,r_n_449__28_,r_n_449__27_,r_n_449__26_,
  r_n_449__25_,r_n_449__24_,r_n_449__23_,r_n_449__22_,r_n_449__21_,r_n_449__20_,
  r_n_449__19_,r_n_449__18_,r_n_449__17_,r_n_449__16_,r_n_449__15_,r_n_449__14_,r_n_449__13_,
  r_n_449__12_,r_n_449__11_,r_n_449__10_,r_n_449__9_,r_n_449__8_,r_n_449__7_,
  r_n_449__6_,r_n_449__5_,r_n_449__4_,r_n_449__3_,r_n_449__2_,r_n_449__1_,r_n_449__0_,
  r_n_464__63_,r_n_464__62_,r_n_464__61_,r_n_464__60_,r_n_464__59_,r_n_464__58_,
  r_n_464__57_,r_n_464__56_,r_n_464__55_,r_n_464__54_,r_n_464__53_,r_n_464__52_,
  r_n_464__51_,r_n_464__50_,r_n_464__49_,r_n_464__48_,r_n_464__47_,r_n_464__46_,
  r_n_464__45_,r_n_464__44_,r_n_464__43_,r_n_464__42_,r_n_464__41_,r_n_464__40_,
  r_n_464__39_,r_n_464__38_,r_n_464__37_,r_n_464__36_,r_n_464__35_,r_n_464__34_,
  r_n_464__33_,r_n_464__32_,r_n_464__31_,r_n_464__30_,r_n_464__29_,r_n_464__28_,r_n_464__27_,
  r_n_464__26_,r_n_464__25_,r_n_464__24_,r_n_464__23_,r_n_464__22_,r_n_464__21_,
  r_n_464__20_,r_n_464__19_,r_n_464__18_,r_n_464__17_,r_n_464__16_,r_n_464__15_,
  r_n_464__14_,r_n_464__13_,r_n_464__12_,r_n_464__11_,r_n_464__10_,r_n_464__9_,
  r_n_464__8_,r_n_464__7_,r_n_464__6_,r_n_464__5_,r_n_464__4_,r_n_464__3_,r_n_464__2_,
  r_n_464__1_,r_n_464__0_,r_n_463__63_,r_n_463__62_,r_n_463__61_,r_n_463__60_,
  r_n_463__59_,r_n_463__58_,r_n_463__57_,r_n_463__56_,r_n_463__55_,r_n_463__54_,
  r_n_463__53_,r_n_463__52_,r_n_463__51_,r_n_463__50_,r_n_463__49_,r_n_463__48_,
  r_n_463__47_,r_n_463__46_,r_n_463__45_,r_n_463__44_,r_n_463__43_,r_n_463__42_,r_n_463__41_,
  r_n_463__40_,r_n_463__39_,r_n_463__38_,r_n_463__37_,r_n_463__36_,r_n_463__35_,
  r_n_463__34_,r_n_463__33_,r_n_463__32_,r_n_463__31_,r_n_463__30_,r_n_463__29_,
  r_n_463__28_,r_n_463__27_,r_n_463__26_,r_n_463__25_,r_n_463__24_,r_n_463__23_,
  r_n_463__22_,r_n_463__21_,r_n_463__20_,r_n_463__19_,r_n_463__18_,r_n_463__17_,
  r_n_463__16_,r_n_463__15_,r_n_463__14_,r_n_463__13_,r_n_463__12_,r_n_463__11_,
  r_n_463__10_,r_n_463__9_,r_n_463__8_,r_n_463__7_,r_n_463__6_,r_n_463__5_,r_n_463__4_,
  r_n_463__3_,r_n_463__2_,r_n_463__1_,r_n_463__0_,r_n_462__63_,r_n_462__62_,
  r_n_462__61_,r_n_462__60_,r_n_462__59_,r_n_462__58_,r_n_462__57_,r_n_462__56_,r_n_462__55_,
  r_n_462__54_,r_n_462__53_,r_n_462__52_,r_n_462__51_,r_n_462__50_,r_n_462__49_,
  r_n_462__48_,r_n_462__47_,r_n_462__46_,r_n_462__45_,r_n_462__44_,r_n_462__43_,
  r_n_462__42_,r_n_462__41_,r_n_462__40_,r_n_462__39_,r_n_462__38_,r_n_462__37_,
  r_n_462__36_,r_n_462__35_,r_n_462__34_,r_n_462__33_,r_n_462__32_,r_n_462__31_,
  r_n_462__30_,r_n_462__29_,r_n_462__28_,r_n_462__27_,r_n_462__26_,r_n_462__25_,
  r_n_462__24_,r_n_462__23_,r_n_462__22_,r_n_462__21_,r_n_462__20_,r_n_462__19_,r_n_462__18_,
  r_n_462__17_,r_n_462__16_,r_n_462__15_,r_n_462__14_,r_n_462__13_,r_n_462__12_,
  r_n_462__11_,r_n_462__10_,r_n_462__9_,r_n_462__8_,r_n_462__7_,r_n_462__6_,
  r_n_462__5_,r_n_462__4_,r_n_462__3_,r_n_462__2_,r_n_462__1_,r_n_462__0_,r_n_461__63_,
  r_n_461__62_,r_n_461__61_,r_n_461__60_,r_n_461__59_,r_n_461__58_,r_n_461__57_,
  r_n_461__56_,r_n_461__55_,r_n_461__54_,r_n_461__53_,r_n_461__52_,r_n_461__51_,
  r_n_461__50_,r_n_461__49_,r_n_461__48_,r_n_461__47_,r_n_461__46_,r_n_461__45_,
  r_n_461__44_,r_n_461__43_,r_n_461__42_,r_n_461__41_,r_n_461__40_,r_n_461__39_,
  r_n_461__38_,r_n_461__37_,r_n_461__36_,r_n_461__35_,r_n_461__34_,r_n_461__33_,r_n_461__32_,
  r_n_461__31_,r_n_461__30_,r_n_461__29_,r_n_461__28_,r_n_461__27_,r_n_461__26_,
  r_n_461__25_,r_n_461__24_,r_n_461__23_,r_n_461__22_,r_n_461__21_,r_n_461__20_,
  r_n_461__19_,r_n_461__18_,r_n_461__17_,r_n_461__16_,r_n_461__15_,r_n_461__14_,
  r_n_461__13_,r_n_461__12_,r_n_461__11_,r_n_461__10_,r_n_461__9_,r_n_461__8_,
  r_n_461__7_,r_n_461__6_,r_n_461__5_,r_n_461__4_,r_n_461__3_,r_n_461__2_,r_n_461__1_,
  r_n_461__0_,r_n_460__63_,r_n_460__62_,r_n_460__61_,r_n_460__60_,r_n_460__59_,
  r_n_460__58_,r_n_460__57_,r_n_460__56_,r_n_460__55_,r_n_460__54_,r_n_460__53_,
  r_n_460__52_,r_n_460__51_,r_n_460__50_,r_n_460__49_,r_n_460__48_,r_n_460__47_,r_n_460__46_,
  r_n_460__45_,r_n_460__44_,r_n_460__43_,r_n_460__42_,r_n_460__41_,r_n_460__40_,
  r_n_460__39_,r_n_460__38_,r_n_460__37_,r_n_460__36_,r_n_460__35_,r_n_460__34_,
  r_n_460__33_,r_n_460__32_,r_n_460__31_,r_n_460__30_,r_n_460__29_,r_n_460__28_,
  r_n_460__27_,r_n_460__26_,r_n_460__25_,r_n_460__24_,r_n_460__23_,r_n_460__22_,
  r_n_460__21_,r_n_460__20_,r_n_460__19_,r_n_460__18_,r_n_460__17_,r_n_460__16_,
  r_n_460__15_,r_n_460__14_,r_n_460__13_,r_n_460__12_,r_n_460__11_,r_n_460__10_,r_n_460__9_,
  r_n_460__8_,r_n_460__7_,r_n_460__6_,r_n_460__5_,r_n_460__4_,r_n_460__3_,
  r_n_460__2_,r_n_460__1_,r_n_460__0_,r_n_459__63_,r_n_459__62_,r_n_459__61_,r_n_459__60_,
  r_n_459__59_,r_n_459__58_,r_n_459__57_,r_n_459__56_,r_n_459__55_,r_n_459__54_,
  r_n_459__53_,r_n_459__52_,r_n_459__51_,r_n_459__50_,r_n_459__49_,r_n_459__48_,
  r_n_459__47_,r_n_459__46_,r_n_459__45_,r_n_459__44_,r_n_459__43_,r_n_459__42_,
  r_n_459__41_,r_n_459__40_,r_n_459__39_,r_n_459__38_,r_n_459__37_,r_n_459__36_,
  r_n_459__35_,r_n_459__34_,r_n_459__33_,r_n_459__32_,r_n_459__31_,r_n_459__30_,
  r_n_459__29_,r_n_459__28_,r_n_459__27_,r_n_459__26_,r_n_459__25_,r_n_459__24_,
  r_n_459__23_,r_n_459__22_,r_n_459__21_,r_n_459__20_,r_n_459__19_,r_n_459__18_,r_n_459__17_,
  r_n_459__16_,r_n_459__15_,r_n_459__14_,r_n_459__13_,r_n_459__12_,r_n_459__11_,
  r_n_459__10_,r_n_459__9_,r_n_459__8_,r_n_459__7_,r_n_459__6_,r_n_459__5_,
  r_n_459__4_,r_n_459__3_,r_n_459__2_,r_n_459__1_,r_n_459__0_,r_n_458__63_,r_n_458__62_,
  r_n_458__61_,r_n_458__60_,r_n_458__59_,r_n_458__58_,r_n_458__57_,r_n_458__56_,
  r_n_458__55_,r_n_458__54_,r_n_458__53_,r_n_458__52_,r_n_458__51_,r_n_458__50_,
  r_n_458__49_,r_n_458__48_,r_n_458__47_,r_n_458__46_,r_n_458__45_,r_n_458__44_,
  r_n_458__43_,r_n_458__42_,r_n_458__41_,r_n_458__40_,r_n_458__39_,r_n_458__38_,
  r_n_458__37_,r_n_458__36_,r_n_458__35_,r_n_458__34_,r_n_458__33_,r_n_458__32_,r_n_458__31_,
  r_n_458__30_,r_n_458__29_,r_n_458__28_,r_n_458__27_,r_n_458__26_,r_n_458__25_,
  r_n_458__24_,r_n_458__23_,r_n_458__22_,r_n_458__21_,r_n_458__20_,r_n_458__19_,
  r_n_458__18_,r_n_458__17_,r_n_458__16_,r_n_458__15_,r_n_458__14_,r_n_458__13_,
  r_n_458__12_,r_n_458__11_,r_n_458__10_,r_n_458__9_,r_n_458__8_,r_n_458__7_,r_n_458__6_,
  r_n_458__5_,r_n_458__4_,r_n_458__3_,r_n_458__2_,r_n_458__1_,r_n_458__0_,
  r_n_457__63_,r_n_457__62_,r_n_457__61_,r_n_457__60_,r_n_457__59_,r_n_457__58_,
  r_n_457__57_,r_n_457__56_,r_n_457__55_,r_n_457__54_,r_n_457__53_,r_n_457__52_,
  r_n_457__51_,r_n_457__50_,r_n_457__49_,r_n_457__48_,r_n_457__47_,r_n_457__46_,r_n_457__45_,
  r_n_457__44_,r_n_457__43_,r_n_457__42_,r_n_457__41_,r_n_457__40_,r_n_457__39_,
  r_n_457__38_,r_n_457__37_,r_n_457__36_,r_n_457__35_,r_n_457__34_,r_n_457__33_,
  r_n_457__32_,r_n_457__31_,r_n_457__30_,r_n_457__29_,r_n_457__28_,r_n_457__27_,
  r_n_457__26_,r_n_457__25_,r_n_457__24_,r_n_457__23_,r_n_457__22_,r_n_457__21_,
  r_n_457__20_,r_n_457__19_,r_n_457__18_,r_n_457__17_,r_n_457__16_,r_n_457__15_,
  r_n_457__14_,r_n_457__13_,r_n_457__12_,r_n_457__11_,r_n_457__10_,r_n_457__9_,r_n_457__8_,
  r_n_457__7_,r_n_457__6_,r_n_457__5_,r_n_457__4_,r_n_457__3_,r_n_457__2_,
  r_n_457__1_,r_n_457__0_,r_n_472__63_,r_n_472__62_,r_n_472__61_,r_n_472__60_,r_n_472__59_,
  r_n_472__58_,r_n_472__57_,r_n_472__56_,r_n_472__55_,r_n_472__54_,r_n_472__53_,
  r_n_472__52_,r_n_472__51_,r_n_472__50_,r_n_472__49_,r_n_472__48_,r_n_472__47_,
  r_n_472__46_,r_n_472__45_,r_n_472__44_,r_n_472__43_,r_n_472__42_,r_n_472__41_,
  r_n_472__40_,r_n_472__39_,r_n_472__38_,r_n_472__37_,r_n_472__36_,r_n_472__35_,
  r_n_472__34_,r_n_472__33_,r_n_472__32_,r_n_472__31_,r_n_472__30_,r_n_472__29_,
  r_n_472__28_,r_n_472__27_,r_n_472__26_,r_n_472__25_,r_n_472__24_,r_n_472__23_,r_n_472__22_,
  r_n_472__21_,r_n_472__20_,r_n_472__19_,r_n_472__18_,r_n_472__17_,r_n_472__16_,
  r_n_472__15_,r_n_472__14_,r_n_472__13_,r_n_472__12_,r_n_472__11_,r_n_472__10_,
  r_n_472__9_,r_n_472__8_,r_n_472__7_,r_n_472__6_,r_n_472__5_,r_n_472__4_,r_n_472__3_,
  r_n_472__2_,r_n_472__1_,r_n_472__0_,r_n_471__63_,r_n_471__62_,r_n_471__61_,
  r_n_471__60_,r_n_471__59_,r_n_471__58_,r_n_471__57_,r_n_471__56_,r_n_471__55_,
  r_n_471__54_,r_n_471__53_,r_n_471__52_,r_n_471__51_,r_n_471__50_,r_n_471__49_,
  r_n_471__48_,r_n_471__47_,r_n_471__46_,r_n_471__45_,r_n_471__44_,r_n_471__43_,
  r_n_471__42_,r_n_471__41_,r_n_471__40_,r_n_471__39_,r_n_471__38_,r_n_471__37_,r_n_471__36_,
  r_n_471__35_,r_n_471__34_,r_n_471__33_,r_n_471__32_,r_n_471__31_,r_n_471__30_,
  r_n_471__29_,r_n_471__28_,r_n_471__27_,r_n_471__26_,r_n_471__25_,r_n_471__24_,
  r_n_471__23_,r_n_471__22_,r_n_471__21_,r_n_471__20_,r_n_471__19_,r_n_471__18_,
  r_n_471__17_,r_n_471__16_,r_n_471__15_,r_n_471__14_,r_n_471__13_,r_n_471__12_,
  r_n_471__11_,r_n_471__10_,r_n_471__9_,r_n_471__8_,r_n_471__7_,r_n_471__6_,r_n_471__5_,
  r_n_471__4_,r_n_471__3_,r_n_471__2_,r_n_471__1_,r_n_471__0_,r_n_470__63_,
  r_n_470__62_,r_n_470__61_,r_n_470__60_,r_n_470__59_,r_n_470__58_,r_n_470__57_,
  r_n_470__56_,r_n_470__55_,r_n_470__54_,r_n_470__53_,r_n_470__52_,r_n_470__51_,r_n_470__50_,
  r_n_470__49_,r_n_470__48_,r_n_470__47_,r_n_470__46_,r_n_470__45_,r_n_470__44_,
  r_n_470__43_,r_n_470__42_,r_n_470__41_,r_n_470__40_,r_n_470__39_,r_n_470__38_,
  r_n_470__37_,r_n_470__36_,r_n_470__35_,r_n_470__34_,r_n_470__33_,r_n_470__32_,
  r_n_470__31_,r_n_470__30_,r_n_470__29_,r_n_470__28_,r_n_470__27_,r_n_470__26_,
  r_n_470__25_,r_n_470__24_,r_n_470__23_,r_n_470__22_,r_n_470__21_,r_n_470__20_,
  r_n_470__19_,r_n_470__18_,r_n_470__17_,r_n_470__16_,r_n_470__15_,r_n_470__14_,
  r_n_470__13_,r_n_470__12_,r_n_470__11_,r_n_470__10_,r_n_470__9_,r_n_470__8_,r_n_470__7_,
  r_n_470__6_,r_n_470__5_,r_n_470__4_,r_n_470__3_,r_n_470__2_,r_n_470__1_,r_n_470__0_,
  r_n_469__63_,r_n_469__62_,r_n_469__61_,r_n_469__60_,r_n_469__59_,r_n_469__58_,
  r_n_469__57_,r_n_469__56_,r_n_469__55_,r_n_469__54_,r_n_469__53_,r_n_469__52_,
  r_n_469__51_,r_n_469__50_,r_n_469__49_,r_n_469__48_,r_n_469__47_,r_n_469__46_,
  r_n_469__45_,r_n_469__44_,r_n_469__43_,r_n_469__42_,r_n_469__41_,r_n_469__40_,
  r_n_469__39_,r_n_469__38_,r_n_469__37_,r_n_469__36_,r_n_469__35_,r_n_469__34_,
  r_n_469__33_,r_n_469__32_,r_n_469__31_,r_n_469__30_,r_n_469__29_,r_n_469__28_,
  r_n_469__27_,r_n_469__26_,r_n_469__25_,r_n_469__24_,r_n_469__23_,r_n_469__22_,r_n_469__21_,
  r_n_469__20_,r_n_469__19_,r_n_469__18_,r_n_469__17_,r_n_469__16_,r_n_469__15_,
  r_n_469__14_,r_n_469__13_,r_n_469__12_,r_n_469__11_,r_n_469__10_,r_n_469__9_,
  r_n_469__8_,r_n_469__7_,r_n_469__6_,r_n_469__5_,r_n_469__4_,r_n_469__3_,r_n_469__2_,
  r_n_469__1_,r_n_469__0_,r_n_468__63_,r_n_468__62_,r_n_468__61_,r_n_468__60_,
  r_n_468__59_,r_n_468__58_,r_n_468__57_,r_n_468__56_,r_n_468__55_,r_n_468__54_,
  r_n_468__53_,r_n_468__52_,r_n_468__51_,r_n_468__50_,r_n_468__49_,r_n_468__48_,
  r_n_468__47_,r_n_468__46_,r_n_468__45_,r_n_468__44_,r_n_468__43_,r_n_468__42_,
  r_n_468__41_,r_n_468__40_,r_n_468__39_,r_n_468__38_,r_n_468__37_,r_n_468__36_,r_n_468__35_,
  r_n_468__34_,r_n_468__33_,r_n_468__32_,r_n_468__31_,r_n_468__30_,r_n_468__29_,
  r_n_468__28_,r_n_468__27_,r_n_468__26_,r_n_468__25_,r_n_468__24_,r_n_468__23_,
  r_n_468__22_,r_n_468__21_,r_n_468__20_,r_n_468__19_,r_n_468__18_,r_n_468__17_,
  r_n_468__16_,r_n_468__15_,r_n_468__14_,r_n_468__13_,r_n_468__12_,r_n_468__11_,
  r_n_468__10_,r_n_468__9_,r_n_468__8_,r_n_468__7_,r_n_468__6_,r_n_468__5_,r_n_468__4_,
  r_n_468__3_,r_n_468__2_,r_n_468__1_,r_n_468__0_,r_n_467__63_,r_n_467__62_,
  r_n_467__61_,r_n_467__60_,r_n_467__59_,r_n_467__58_,r_n_467__57_,r_n_467__56_,
  r_n_467__55_,r_n_467__54_,r_n_467__53_,r_n_467__52_,r_n_467__51_,r_n_467__50_,r_n_467__49_,
  r_n_467__48_,r_n_467__47_,r_n_467__46_,r_n_467__45_,r_n_467__44_,r_n_467__43_,
  r_n_467__42_,r_n_467__41_,r_n_467__40_,r_n_467__39_,r_n_467__38_,r_n_467__37_,
  r_n_467__36_,r_n_467__35_,r_n_467__34_,r_n_467__33_,r_n_467__32_,r_n_467__31_,
  r_n_467__30_,r_n_467__29_,r_n_467__28_,r_n_467__27_,r_n_467__26_,r_n_467__25_,
  r_n_467__24_,r_n_467__23_,r_n_467__22_,r_n_467__21_,r_n_467__20_,r_n_467__19_,
  r_n_467__18_,r_n_467__17_,r_n_467__16_,r_n_467__15_,r_n_467__14_,r_n_467__13_,r_n_467__12_,
  r_n_467__11_,r_n_467__10_,r_n_467__9_,r_n_467__8_,r_n_467__7_,r_n_467__6_,
  r_n_467__5_,r_n_467__4_,r_n_467__3_,r_n_467__2_,r_n_467__1_,r_n_467__0_,r_n_466__63_,
  r_n_466__62_,r_n_466__61_,r_n_466__60_,r_n_466__59_,r_n_466__58_,r_n_466__57_,
  r_n_466__56_,r_n_466__55_,r_n_466__54_,r_n_466__53_,r_n_466__52_,r_n_466__51_,
  r_n_466__50_,r_n_466__49_,r_n_466__48_,r_n_466__47_,r_n_466__46_,r_n_466__45_,
  r_n_466__44_,r_n_466__43_,r_n_466__42_,r_n_466__41_,r_n_466__40_,r_n_466__39_,
  r_n_466__38_,r_n_466__37_,r_n_466__36_,r_n_466__35_,r_n_466__34_,r_n_466__33_,
  r_n_466__32_,r_n_466__31_,r_n_466__30_,r_n_466__29_,r_n_466__28_,r_n_466__27_,r_n_466__26_,
  r_n_466__25_,r_n_466__24_,r_n_466__23_,r_n_466__22_,r_n_466__21_,r_n_466__20_,
  r_n_466__19_,r_n_466__18_,r_n_466__17_,r_n_466__16_,r_n_466__15_,r_n_466__14_,
  r_n_466__13_,r_n_466__12_,r_n_466__11_,r_n_466__10_,r_n_466__9_,r_n_466__8_,
  r_n_466__7_,r_n_466__6_,r_n_466__5_,r_n_466__4_,r_n_466__3_,r_n_466__2_,r_n_466__1_,
  r_n_466__0_,r_n_465__63_,r_n_465__62_,r_n_465__61_,r_n_465__60_,r_n_465__59_,
  r_n_465__58_,r_n_465__57_,r_n_465__56_,r_n_465__55_,r_n_465__54_,r_n_465__53_,
  r_n_465__52_,r_n_465__51_,r_n_465__50_,r_n_465__49_,r_n_465__48_,r_n_465__47_,
  r_n_465__46_,r_n_465__45_,r_n_465__44_,r_n_465__43_,r_n_465__42_,r_n_465__41_,r_n_465__40_,
  r_n_465__39_,r_n_465__38_,r_n_465__37_,r_n_465__36_,r_n_465__35_,r_n_465__34_,
  r_n_465__33_,r_n_465__32_,r_n_465__31_,r_n_465__30_,r_n_465__29_,r_n_465__28_,
  r_n_465__27_,r_n_465__26_,r_n_465__25_,r_n_465__24_,r_n_465__23_,r_n_465__22_,
  r_n_465__21_,r_n_465__20_,r_n_465__19_,r_n_465__18_,r_n_465__17_,r_n_465__16_,
  r_n_465__15_,r_n_465__14_,r_n_465__13_,r_n_465__12_,r_n_465__11_,r_n_465__10_,
  r_n_465__9_,r_n_465__8_,r_n_465__7_,r_n_465__6_,r_n_465__5_,r_n_465__4_,r_n_465__3_,
  r_n_465__2_,r_n_465__1_,r_n_465__0_,r_n_480__63_,r_n_480__62_,r_n_480__61_,
  r_n_480__60_,r_n_480__59_,r_n_480__58_,r_n_480__57_,r_n_480__56_,r_n_480__55_,r_n_480__54_,
  r_n_480__53_,r_n_480__52_,r_n_480__51_,r_n_480__50_,r_n_480__49_,r_n_480__48_,
  r_n_480__47_,r_n_480__46_,r_n_480__45_,r_n_480__44_,r_n_480__43_,r_n_480__42_,
  r_n_480__41_,r_n_480__40_,r_n_480__39_,r_n_480__38_,r_n_480__37_,r_n_480__36_,
  r_n_480__35_,r_n_480__34_,r_n_480__33_,r_n_480__32_,r_n_480__31_,r_n_480__30_,
  r_n_480__29_,r_n_480__28_,r_n_480__27_,r_n_480__26_,r_n_480__25_,r_n_480__24_,
  r_n_480__23_,r_n_480__22_,r_n_480__21_,r_n_480__20_,r_n_480__19_,r_n_480__18_,
  r_n_480__17_,r_n_480__16_,r_n_480__15_,r_n_480__14_,r_n_480__13_,r_n_480__12_,r_n_480__11_,
  r_n_480__10_,r_n_480__9_,r_n_480__8_,r_n_480__7_,r_n_480__6_,r_n_480__5_,
  r_n_480__4_,r_n_480__3_,r_n_480__2_,r_n_480__1_,r_n_480__0_,r_n_479__63_,r_n_479__62_,
  r_n_479__61_,r_n_479__60_,r_n_479__59_,r_n_479__58_,r_n_479__57_,r_n_479__56_,
  r_n_479__55_,r_n_479__54_,r_n_479__53_,r_n_479__52_,r_n_479__51_,r_n_479__50_,
  r_n_479__49_,r_n_479__48_,r_n_479__47_,r_n_479__46_,r_n_479__45_,r_n_479__44_,
  r_n_479__43_,r_n_479__42_,r_n_479__41_,r_n_479__40_,r_n_479__39_,r_n_479__38_,
  r_n_479__37_,r_n_479__36_,r_n_479__35_,r_n_479__34_,r_n_479__33_,r_n_479__32_,
  r_n_479__31_,r_n_479__30_,r_n_479__29_,r_n_479__28_,r_n_479__27_,r_n_479__26_,r_n_479__25_,
  r_n_479__24_,r_n_479__23_,r_n_479__22_,r_n_479__21_,r_n_479__20_,r_n_479__19_,
  r_n_479__18_,r_n_479__17_,r_n_479__16_,r_n_479__15_,r_n_479__14_,r_n_479__13_,
  r_n_479__12_,r_n_479__11_,r_n_479__10_,r_n_479__9_,r_n_479__8_,r_n_479__7_,
  r_n_479__6_,r_n_479__5_,r_n_479__4_,r_n_479__3_,r_n_479__2_,r_n_479__1_,r_n_479__0_,
  r_n_478__63_,r_n_478__62_,r_n_478__61_,r_n_478__60_,r_n_478__59_,r_n_478__58_,
  r_n_478__57_,r_n_478__56_,r_n_478__55_,r_n_478__54_,r_n_478__53_,r_n_478__52_,
  r_n_478__51_,r_n_478__50_,r_n_478__49_,r_n_478__48_,r_n_478__47_,r_n_478__46_,
  r_n_478__45_,r_n_478__44_,r_n_478__43_,r_n_478__42_,r_n_478__41_,r_n_478__40_,r_n_478__39_,
  r_n_478__38_,r_n_478__37_,r_n_478__36_,r_n_478__35_,r_n_478__34_,r_n_478__33_,
  r_n_478__32_,r_n_478__31_,r_n_478__30_,r_n_478__29_,r_n_478__28_,r_n_478__27_,
  r_n_478__26_,r_n_478__25_,r_n_478__24_,r_n_478__23_,r_n_478__22_,r_n_478__21_,
  r_n_478__20_,r_n_478__19_,r_n_478__18_,r_n_478__17_,r_n_478__16_,r_n_478__15_,
  r_n_478__14_,r_n_478__13_,r_n_478__12_,r_n_478__11_,r_n_478__10_,r_n_478__9_,r_n_478__8_,
  r_n_478__7_,r_n_478__6_,r_n_478__5_,r_n_478__4_,r_n_478__3_,r_n_478__2_,
  r_n_478__1_,r_n_478__0_,r_n_477__63_,r_n_477__62_,r_n_477__61_,r_n_477__60_,
  r_n_477__59_,r_n_477__58_,r_n_477__57_,r_n_477__56_,r_n_477__55_,r_n_477__54_,r_n_477__53_,
  r_n_477__52_,r_n_477__51_,r_n_477__50_,r_n_477__49_,r_n_477__48_,r_n_477__47_,
  r_n_477__46_,r_n_477__45_,r_n_477__44_,r_n_477__43_,r_n_477__42_,r_n_477__41_,
  r_n_477__40_,r_n_477__39_,r_n_477__38_,r_n_477__37_,r_n_477__36_,r_n_477__35_,
  r_n_477__34_,r_n_477__33_,r_n_477__32_,r_n_477__31_,r_n_477__30_,r_n_477__29_,
  r_n_477__28_,r_n_477__27_,r_n_477__26_,r_n_477__25_,r_n_477__24_,r_n_477__23_,
  r_n_477__22_,r_n_477__21_,r_n_477__20_,r_n_477__19_,r_n_477__18_,r_n_477__17_,r_n_477__16_,
  r_n_477__15_,r_n_477__14_,r_n_477__13_,r_n_477__12_,r_n_477__11_,r_n_477__10_,
  r_n_477__9_,r_n_477__8_,r_n_477__7_,r_n_477__6_,r_n_477__5_,r_n_477__4_,
  r_n_477__3_,r_n_477__2_,r_n_477__1_,r_n_477__0_,r_n_476__63_,r_n_476__62_,r_n_476__61_,
  r_n_476__60_,r_n_476__59_,r_n_476__58_,r_n_476__57_,r_n_476__56_,r_n_476__55_,
  r_n_476__54_,r_n_476__53_,r_n_476__52_,r_n_476__51_,r_n_476__50_,r_n_476__49_,
  r_n_476__48_,r_n_476__47_,r_n_476__46_,r_n_476__45_,r_n_476__44_,r_n_476__43_,
  r_n_476__42_,r_n_476__41_,r_n_476__40_,r_n_476__39_,r_n_476__38_,r_n_476__37_,
  r_n_476__36_,r_n_476__35_,r_n_476__34_,r_n_476__33_,r_n_476__32_,r_n_476__31_,r_n_476__30_,
  r_n_476__29_,r_n_476__28_,r_n_476__27_,r_n_476__26_,r_n_476__25_,r_n_476__24_,
  r_n_476__23_,r_n_476__22_,r_n_476__21_,r_n_476__20_,r_n_476__19_,r_n_476__18_,
  r_n_476__17_,r_n_476__16_,r_n_476__15_,r_n_476__14_,r_n_476__13_,r_n_476__12_,
  r_n_476__11_,r_n_476__10_,r_n_476__9_,r_n_476__8_,r_n_476__7_,r_n_476__6_,r_n_476__5_,
  r_n_476__4_,r_n_476__3_,r_n_476__2_,r_n_476__1_,r_n_476__0_,r_n_475__63_,
  r_n_475__62_,r_n_475__61_,r_n_475__60_,r_n_475__59_,r_n_475__58_,r_n_475__57_,
  r_n_475__56_,r_n_475__55_,r_n_475__54_,r_n_475__53_,r_n_475__52_,r_n_475__51_,
  r_n_475__50_,r_n_475__49_,r_n_475__48_,r_n_475__47_,r_n_475__46_,r_n_475__45_,r_n_475__44_,
  r_n_475__43_,r_n_475__42_,r_n_475__41_,r_n_475__40_,r_n_475__39_,r_n_475__38_,
  r_n_475__37_,r_n_475__36_,r_n_475__35_,r_n_475__34_,r_n_475__33_,r_n_475__32_,
  r_n_475__31_,r_n_475__30_,r_n_475__29_,r_n_475__28_,r_n_475__27_,r_n_475__26_,
  r_n_475__25_,r_n_475__24_,r_n_475__23_,r_n_475__22_,r_n_475__21_,r_n_475__20_,
  r_n_475__19_,r_n_475__18_,r_n_475__17_,r_n_475__16_,r_n_475__15_,r_n_475__14_,
  r_n_475__13_,r_n_475__12_,r_n_475__11_,r_n_475__10_,r_n_475__9_,r_n_475__8_,r_n_475__7_,
  r_n_475__6_,r_n_475__5_,r_n_475__4_,r_n_475__3_,r_n_475__2_,r_n_475__1_,
  r_n_475__0_,r_n_474__63_,r_n_474__62_,r_n_474__61_,r_n_474__60_,r_n_474__59_,r_n_474__58_,
  r_n_474__57_,r_n_474__56_,r_n_474__55_,r_n_474__54_,r_n_474__53_,r_n_474__52_,
  r_n_474__51_,r_n_474__50_,r_n_474__49_,r_n_474__48_,r_n_474__47_,r_n_474__46_,
  r_n_474__45_,r_n_474__44_,r_n_474__43_,r_n_474__42_,r_n_474__41_,r_n_474__40_,
  r_n_474__39_,r_n_474__38_,r_n_474__37_,r_n_474__36_,r_n_474__35_,r_n_474__34_,
  r_n_474__33_,r_n_474__32_,r_n_474__31_,r_n_474__30_,r_n_474__29_,r_n_474__28_,
  r_n_474__27_,r_n_474__26_,r_n_474__25_,r_n_474__24_,r_n_474__23_,r_n_474__22_,
  r_n_474__21_,r_n_474__20_,r_n_474__19_,r_n_474__18_,r_n_474__17_,r_n_474__16_,r_n_474__15_,
  r_n_474__14_,r_n_474__13_,r_n_474__12_,r_n_474__11_,r_n_474__10_,r_n_474__9_,
  r_n_474__8_,r_n_474__7_,r_n_474__6_,r_n_474__5_,r_n_474__4_,r_n_474__3_,r_n_474__2_,
  r_n_474__1_,r_n_474__0_,r_n_473__63_,r_n_473__62_,r_n_473__61_,r_n_473__60_,
  r_n_473__59_,r_n_473__58_,r_n_473__57_,r_n_473__56_,r_n_473__55_,r_n_473__54_,
  r_n_473__53_,r_n_473__52_,r_n_473__51_,r_n_473__50_,r_n_473__49_,r_n_473__48_,
  r_n_473__47_,r_n_473__46_,r_n_473__45_,r_n_473__44_,r_n_473__43_,r_n_473__42_,
  r_n_473__41_,r_n_473__40_,r_n_473__39_,r_n_473__38_,r_n_473__37_,r_n_473__36_,
  r_n_473__35_,r_n_473__34_,r_n_473__33_,r_n_473__32_,r_n_473__31_,r_n_473__30_,r_n_473__29_,
  r_n_473__28_,r_n_473__27_,r_n_473__26_,r_n_473__25_,r_n_473__24_,r_n_473__23_,
  r_n_473__22_,r_n_473__21_,r_n_473__20_,r_n_473__19_,r_n_473__18_,r_n_473__17_,
  r_n_473__16_,r_n_473__15_,r_n_473__14_,r_n_473__13_,r_n_473__12_,r_n_473__11_,
  r_n_473__10_,r_n_473__9_,r_n_473__8_,r_n_473__7_,r_n_473__6_,r_n_473__5_,r_n_473__4_,
  r_n_473__3_,r_n_473__2_,r_n_473__1_,r_n_473__0_,r_n_488__63_,r_n_488__62_,
  r_n_488__61_,r_n_488__60_,r_n_488__59_,r_n_488__58_,r_n_488__57_,r_n_488__56_,
  r_n_488__55_,r_n_488__54_,r_n_488__53_,r_n_488__52_,r_n_488__51_,r_n_488__50_,
  r_n_488__49_,r_n_488__48_,r_n_488__47_,r_n_488__46_,r_n_488__45_,r_n_488__44_,r_n_488__43_,
  r_n_488__42_,r_n_488__41_,r_n_488__40_,r_n_488__39_,r_n_488__38_,r_n_488__37_,
  r_n_488__36_,r_n_488__35_,r_n_488__34_,r_n_488__33_,r_n_488__32_,r_n_488__31_,
  r_n_488__30_,r_n_488__29_,r_n_488__28_,r_n_488__27_,r_n_488__26_,r_n_488__25_,
  r_n_488__24_,r_n_488__23_,r_n_488__22_,r_n_488__21_,r_n_488__20_,r_n_488__19_,
  r_n_488__18_,r_n_488__17_,r_n_488__16_,r_n_488__15_,r_n_488__14_,r_n_488__13_,
  r_n_488__12_,r_n_488__11_,r_n_488__10_,r_n_488__9_,r_n_488__8_,r_n_488__7_,r_n_488__6_,
  r_n_488__5_,r_n_488__4_,r_n_488__3_,r_n_488__2_,r_n_488__1_,r_n_488__0_,
  r_n_487__63_,r_n_487__62_,r_n_487__61_,r_n_487__60_,r_n_487__59_,r_n_487__58_,r_n_487__57_,
  r_n_487__56_,r_n_487__55_,r_n_487__54_,r_n_487__53_,r_n_487__52_,r_n_487__51_,
  r_n_487__50_,r_n_487__49_,r_n_487__48_,r_n_487__47_,r_n_487__46_,r_n_487__45_,
  r_n_487__44_,r_n_487__43_,r_n_487__42_,r_n_487__41_,r_n_487__40_,r_n_487__39_,
  r_n_487__38_,r_n_487__37_,r_n_487__36_,r_n_487__35_,r_n_487__34_,r_n_487__33_,
  r_n_487__32_,r_n_487__31_,r_n_487__30_,r_n_487__29_,r_n_487__28_,r_n_487__27_,
  r_n_487__26_,r_n_487__25_,r_n_487__24_,r_n_487__23_,r_n_487__22_,r_n_487__21_,r_n_487__20_,
  r_n_487__19_,r_n_487__18_,r_n_487__17_,r_n_487__16_,r_n_487__15_,r_n_487__14_,
  r_n_487__13_,r_n_487__12_,r_n_487__11_,r_n_487__10_,r_n_487__9_,r_n_487__8_,
  r_n_487__7_,r_n_487__6_,r_n_487__5_,r_n_487__4_,r_n_487__3_,r_n_487__2_,r_n_487__1_,
  r_n_487__0_,r_n_486__63_,r_n_486__62_,r_n_486__61_,r_n_486__60_,r_n_486__59_,
  r_n_486__58_,r_n_486__57_,r_n_486__56_,r_n_486__55_,r_n_486__54_,r_n_486__53_,
  r_n_486__52_,r_n_486__51_,r_n_486__50_,r_n_486__49_,r_n_486__48_,r_n_486__47_,
  r_n_486__46_,r_n_486__45_,r_n_486__44_,r_n_486__43_,r_n_486__42_,r_n_486__41_,
  r_n_486__40_,r_n_486__39_,r_n_486__38_,r_n_486__37_,r_n_486__36_,r_n_486__35_,r_n_486__34_,
  r_n_486__33_,r_n_486__32_,r_n_486__31_,r_n_486__30_,r_n_486__29_,r_n_486__28_,
  r_n_486__27_,r_n_486__26_,r_n_486__25_,r_n_486__24_,r_n_486__23_,r_n_486__22_,
  r_n_486__21_,r_n_486__20_,r_n_486__19_,r_n_486__18_,r_n_486__17_,r_n_486__16_,
  r_n_486__15_,r_n_486__14_,r_n_486__13_,r_n_486__12_,r_n_486__11_,r_n_486__10_,
  r_n_486__9_,r_n_486__8_,r_n_486__7_,r_n_486__6_,r_n_486__5_,r_n_486__4_,r_n_486__3_,
  r_n_486__2_,r_n_486__1_,r_n_486__0_,r_n_485__63_,r_n_485__62_,r_n_485__61_,
  r_n_485__60_,r_n_485__59_,r_n_485__58_,r_n_485__57_,r_n_485__56_,r_n_485__55_,
  r_n_485__54_,r_n_485__53_,r_n_485__52_,r_n_485__51_,r_n_485__50_,r_n_485__49_,r_n_485__48_,
  r_n_485__47_,r_n_485__46_,r_n_485__45_,r_n_485__44_,r_n_485__43_,r_n_485__42_,
  r_n_485__41_,r_n_485__40_,r_n_485__39_,r_n_485__38_,r_n_485__37_,r_n_485__36_,
  r_n_485__35_,r_n_485__34_,r_n_485__33_,r_n_485__32_,r_n_485__31_,r_n_485__30_,
  r_n_485__29_,r_n_485__28_,r_n_485__27_,r_n_485__26_,r_n_485__25_,r_n_485__24_,
  r_n_485__23_,r_n_485__22_,r_n_485__21_,r_n_485__20_,r_n_485__19_,r_n_485__18_,
  r_n_485__17_,r_n_485__16_,r_n_485__15_,r_n_485__14_,r_n_485__13_,r_n_485__12_,
  r_n_485__11_,r_n_485__10_,r_n_485__9_,r_n_485__8_,r_n_485__7_,r_n_485__6_,r_n_485__5_,
  r_n_485__4_,r_n_485__3_,r_n_485__2_,r_n_485__1_,r_n_485__0_,r_n_484__63_,r_n_484__62_,
  r_n_484__61_,r_n_484__60_,r_n_484__59_,r_n_484__58_,r_n_484__57_,r_n_484__56_,
  r_n_484__55_,r_n_484__54_,r_n_484__53_,r_n_484__52_,r_n_484__51_,r_n_484__50_,
  r_n_484__49_,r_n_484__48_,r_n_484__47_,r_n_484__46_,r_n_484__45_,r_n_484__44_,
  r_n_484__43_,r_n_484__42_,r_n_484__41_,r_n_484__40_,r_n_484__39_,r_n_484__38_,
  r_n_484__37_,r_n_484__36_,r_n_484__35_,r_n_484__34_,r_n_484__33_,r_n_484__32_,
  r_n_484__31_,r_n_484__30_,r_n_484__29_,r_n_484__28_,r_n_484__27_,r_n_484__26_,
  r_n_484__25_,r_n_484__24_,r_n_484__23_,r_n_484__22_,r_n_484__21_,r_n_484__20_,r_n_484__19_,
  r_n_484__18_,r_n_484__17_,r_n_484__16_,r_n_484__15_,r_n_484__14_,r_n_484__13_,
  r_n_484__12_,r_n_484__11_,r_n_484__10_,r_n_484__9_,r_n_484__8_,r_n_484__7_,
  r_n_484__6_,r_n_484__5_,r_n_484__4_,r_n_484__3_,r_n_484__2_,r_n_484__1_,r_n_484__0_,
  r_n_483__63_,r_n_483__62_,r_n_483__61_,r_n_483__60_,r_n_483__59_,r_n_483__58_,
  r_n_483__57_,r_n_483__56_,r_n_483__55_,r_n_483__54_,r_n_483__53_,r_n_483__52_,
  r_n_483__51_,r_n_483__50_,r_n_483__49_,r_n_483__48_,r_n_483__47_,r_n_483__46_,
  r_n_483__45_,r_n_483__44_,r_n_483__43_,r_n_483__42_,r_n_483__41_,r_n_483__40_,
  r_n_483__39_,r_n_483__38_,r_n_483__37_,r_n_483__36_,r_n_483__35_,r_n_483__34_,r_n_483__33_,
  r_n_483__32_,r_n_483__31_,r_n_483__30_,r_n_483__29_,r_n_483__28_,r_n_483__27_,
  r_n_483__26_,r_n_483__25_,r_n_483__24_,r_n_483__23_,r_n_483__22_,r_n_483__21_,
  r_n_483__20_,r_n_483__19_,r_n_483__18_,r_n_483__17_,r_n_483__16_,r_n_483__15_,
  r_n_483__14_,r_n_483__13_,r_n_483__12_,r_n_483__11_,r_n_483__10_,r_n_483__9_,
  r_n_483__8_,r_n_483__7_,r_n_483__6_,r_n_483__5_,r_n_483__4_,r_n_483__3_,r_n_483__2_,
  r_n_483__1_,r_n_483__0_,r_n_482__63_,r_n_482__62_,r_n_482__61_,r_n_482__60_,
  r_n_482__59_,r_n_482__58_,r_n_482__57_,r_n_482__56_,r_n_482__55_,r_n_482__54_,
  r_n_482__53_,r_n_482__52_,r_n_482__51_,r_n_482__50_,r_n_482__49_,r_n_482__48_,r_n_482__47_,
  r_n_482__46_,r_n_482__45_,r_n_482__44_,r_n_482__43_,r_n_482__42_,r_n_482__41_,
  r_n_482__40_,r_n_482__39_,r_n_482__38_,r_n_482__37_,r_n_482__36_,r_n_482__35_,
  r_n_482__34_,r_n_482__33_,r_n_482__32_,r_n_482__31_,r_n_482__30_,r_n_482__29_,
  r_n_482__28_,r_n_482__27_,r_n_482__26_,r_n_482__25_,r_n_482__24_,r_n_482__23_,
  r_n_482__22_,r_n_482__21_,r_n_482__20_,r_n_482__19_,r_n_482__18_,r_n_482__17_,
  r_n_482__16_,r_n_482__15_,r_n_482__14_,r_n_482__13_,r_n_482__12_,r_n_482__11_,r_n_482__10_,
  r_n_482__9_,r_n_482__8_,r_n_482__7_,r_n_482__6_,r_n_482__5_,r_n_482__4_,
  r_n_482__3_,r_n_482__2_,r_n_482__1_,r_n_482__0_,r_n_481__63_,r_n_481__62_,r_n_481__61_,
  r_n_481__60_,r_n_481__59_,r_n_481__58_,r_n_481__57_,r_n_481__56_,r_n_481__55_,
  r_n_481__54_,r_n_481__53_,r_n_481__52_,r_n_481__51_,r_n_481__50_,r_n_481__49_,
  r_n_481__48_,r_n_481__47_,r_n_481__46_,r_n_481__45_,r_n_481__44_,r_n_481__43_,
  r_n_481__42_,r_n_481__41_,r_n_481__40_,r_n_481__39_,r_n_481__38_,r_n_481__37_,
  r_n_481__36_,r_n_481__35_,r_n_481__34_,r_n_481__33_,r_n_481__32_,r_n_481__31_,
  r_n_481__30_,r_n_481__29_,r_n_481__28_,r_n_481__27_,r_n_481__26_,r_n_481__25_,r_n_481__24_,
  r_n_481__23_,r_n_481__22_,r_n_481__21_,r_n_481__20_,r_n_481__19_,r_n_481__18_,
  r_n_481__17_,r_n_481__16_,r_n_481__15_,r_n_481__14_,r_n_481__13_,r_n_481__12_,
  r_n_481__11_,r_n_481__10_,r_n_481__9_,r_n_481__8_,r_n_481__7_,r_n_481__6_,
  r_n_481__5_,r_n_481__4_,r_n_481__3_,r_n_481__2_,r_n_481__1_,r_n_481__0_,r_n_496__63_,
  r_n_496__62_,r_n_496__61_,r_n_496__60_,r_n_496__59_,r_n_496__58_,r_n_496__57_,
  r_n_496__56_,r_n_496__55_,r_n_496__54_,r_n_496__53_,r_n_496__52_,r_n_496__51_,
  r_n_496__50_,r_n_496__49_,r_n_496__48_,r_n_496__47_,r_n_496__46_,r_n_496__45_,
  r_n_496__44_,r_n_496__43_,r_n_496__42_,r_n_496__41_,r_n_496__40_,r_n_496__39_,r_n_496__38_,
  r_n_496__37_,r_n_496__36_,r_n_496__35_,r_n_496__34_,r_n_496__33_,r_n_496__32_,
  r_n_496__31_,r_n_496__30_,r_n_496__29_,r_n_496__28_,r_n_496__27_,r_n_496__26_,
  r_n_496__25_,r_n_496__24_,r_n_496__23_,r_n_496__22_,r_n_496__21_,r_n_496__20_,
  r_n_496__19_,r_n_496__18_,r_n_496__17_,r_n_496__16_,r_n_496__15_,r_n_496__14_,
  r_n_496__13_,r_n_496__12_,r_n_496__11_,r_n_496__10_,r_n_496__9_,r_n_496__8_,r_n_496__7_,
  r_n_496__6_,r_n_496__5_,r_n_496__4_,r_n_496__3_,r_n_496__2_,r_n_496__1_,
  r_n_496__0_,r_n_495__63_,r_n_495__62_,r_n_495__61_,r_n_495__60_,r_n_495__59_,
  r_n_495__58_,r_n_495__57_,r_n_495__56_,r_n_495__55_,r_n_495__54_,r_n_495__53_,r_n_495__52_,
  r_n_495__51_,r_n_495__50_,r_n_495__49_,r_n_495__48_,r_n_495__47_,r_n_495__46_,
  r_n_495__45_,r_n_495__44_,r_n_495__43_,r_n_495__42_,r_n_495__41_,r_n_495__40_,
  r_n_495__39_,r_n_495__38_,r_n_495__37_,r_n_495__36_,r_n_495__35_,r_n_495__34_,
  r_n_495__33_,r_n_495__32_,r_n_495__31_,r_n_495__30_,r_n_495__29_,r_n_495__28_,
  r_n_495__27_,r_n_495__26_,r_n_495__25_,r_n_495__24_,r_n_495__23_,r_n_495__22_,
  r_n_495__21_,r_n_495__20_,r_n_495__19_,r_n_495__18_,r_n_495__17_,r_n_495__16_,
  r_n_495__15_,r_n_495__14_,r_n_495__13_,r_n_495__12_,r_n_495__11_,r_n_495__10_,r_n_495__9_,
  r_n_495__8_,r_n_495__7_,r_n_495__6_,r_n_495__5_,r_n_495__4_,r_n_495__3_,
  r_n_495__2_,r_n_495__1_,r_n_495__0_,r_n_494__63_,r_n_494__62_,r_n_494__61_,r_n_494__60_,
  r_n_494__59_,r_n_494__58_,r_n_494__57_,r_n_494__56_,r_n_494__55_,r_n_494__54_,
  r_n_494__53_,r_n_494__52_,r_n_494__51_,r_n_494__50_,r_n_494__49_,r_n_494__48_,
  r_n_494__47_,r_n_494__46_,r_n_494__45_,r_n_494__44_,r_n_494__43_,r_n_494__42_,
  r_n_494__41_,r_n_494__40_,r_n_494__39_,r_n_494__38_,r_n_494__37_,r_n_494__36_,
  r_n_494__35_,r_n_494__34_,r_n_494__33_,r_n_494__32_,r_n_494__31_,r_n_494__30_,
  r_n_494__29_,r_n_494__28_,r_n_494__27_,r_n_494__26_,r_n_494__25_,r_n_494__24_,r_n_494__23_,
  r_n_494__22_,r_n_494__21_,r_n_494__20_,r_n_494__19_,r_n_494__18_,r_n_494__17_,
  r_n_494__16_,r_n_494__15_,r_n_494__14_,r_n_494__13_,r_n_494__12_,r_n_494__11_,
  r_n_494__10_,r_n_494__9_,r_n_494__8_,r_n_494__7_,r_n_494__6_,r_n_494__5_,r_n_494__4_,
  r_n_494__3_,r_n_494__2_,r_n_494__1_,r_n_494__0_,r_n_493__63_,r_n_493__62_,
  r_n_493__61_,r_n_493__60_,r_n_493__59_,r_n_493__58_,r_n_493__57_,r_n_493__56_,
  r_n_493__55_,r_n_493__54_,r_n_493__53_,r_n_493__52_,r_n_493__51_,r_n_493__50_,
  r_n_493__49_,r_n_493__48_,r_n_493__47_,r_n_493__46_,r_n_493__45_,r_n_493__44_,
  r_n_493__43_,r_n_493__42_,r_n_493__41_,r_n_493__40_,r_n_493__39_,r_n_493__38_,r_n_493__37_,
  r_n_493__36_,r_n_493__35_,r_n_493__34_,r_n_493__33_,r_n_493__32_,r_n_493__31_,
  r_n_493__30_,r_n_493__29_,r_n_493__28_,r_n_493__27_,r_n_493__26_,r_n_493__25_,
  r_n_493__24_,r_n_493__23_,r_n_493__22_,r_n_493__21_,r_n_493__20_,r_n_493__19_,
  r_n_493__18_,r_n_493__17_,r_n_493__16_,r_n_493__15_,r_n_493__14_,r_n_493__13_,
  r_n_493__12_,r_n_493__11_,r_n_493__10_,r_n_493__9_,r_n_493__8_,r_n_493__7_,r_n_493__6_,
  r_n_493__5_,r_n_493__4_,r_n_493__3_,r_n_493__2_,r_n_493__1_,r_n_493__0_,
  r_n_492__63_,r_n_492__62_,r_n_492__61_,r_n_492__60_,r_n_492__59_,r_n_492__58_,
  r_n_492__57_,r_n_492__56_,r_n_492__55_,r_n_492__54_,r_n_492__53_,r_n_492__52_,r_n_492__51_,
  r_n_492__50_,r_n_492__49_,r_n_492__48_,r_n_492__47_,r_n_492__46_,r_n_492__45_,
  r_n_492__44_,r_n_492__43_,r_n_492__42_,r_n_492__41_,r_n_492__40_,r_n_492__39_,
  r_n_492__38_,r_n_492__37_,r_n_492__36_,r_n_492__35_,r_n_492__34_,r_n_492__33_,
  r_n_492__32_,r_n_492__31_,r_n_492__30_,r_n_492__29_,r_n_492__28_,r_n_492__27_,
  r_n_492__26_,r_n_492__25_,r_n_492__24_,r_n_492__23_,r_n_492__22_,r_n_492__21_,
  r_n_492__20_,r_n_492__19_,r_n_492__18_,r_n_492__17_,r_n_492__16_,r_n_492__15_,r_n_492__14_,
  r_n_492__13_,r_n_492__12_,r_n_492__11_,r_n_492__10_,r_n_492__9_,r_n_492__8_,
  r_n_492__7_,r_n_492__6_,r_n_492__5_,r_n_492__4_,r_n_492__3_,r_n_492__2_,r_n_492__1_,
  r_n_492__0_,r_n_491__63_,r_n_491__62_,r_n_491__61_,r_n_491__60_,r_n_491__59_,
  r_n_491__58_,r_n_491__57_,r_n_491__56_,r_n_491__55_,r_n_491__54_,r_n_491__53_,
  r_n_491__52_,r_n_491__51_,r_n_491__50_,r_n_491__49_,r_n_491__48_,r_n_491__47_,
  r_n_491__46_,r_n_491__45_,r_n_491__44_,r_n_491__43_,r_n_491__42_,r_n_491__41_,
  r_n_491__40_,r_n_491__39_,r_n_491__38_,r_n_491__37_,r_n_491__36_,r_n_491__35_,
  r_n_491__34_,r_n_491__33_,r_n_491__32_,r_n_491__31_,r_n_491__30_,r_n_491__29_,r_n_491__28_,
  r_n_491__27_,r_n_491__26_,r_n_491__25_,r_n_491__24_,r_n_491__23_,r_n_491__22_,
  r_n_491__21_,r_n_491__20_,r_n_491__19_,r_n_491__18_,r_n_491__17_,r_n_491__16_,
  r_n_491__15_,r_n_491__14_,r_n_491__13_,r_n_491__12_,r_n_491__11_,r_n_491__10_,
  r_n_491__9_,r_n_491__8_,r_n_491__7_,r_n_491__6_,r_n_491__5_,r_n_491__4_,r_n_491__3_,
  r_n_491__2_,r_n_491__1_,r_n_491__0_,r_n_490__63_,r_n_490__62_,r_n_490__61_,
  r_n_490__60_,r_n_490__59_,r_n_490__58_,r_n_490__57_,r_n_490__56_,r_n_490__55_,
  r_n_490__54_,r_n_490__53_,r_n_490__52_,r_n_490__51_,r_n_490__50_,r_n_490__49_,
  r_n_490__48_,r_n_490__47_,r_n_490__46_,r_n_490__45_,r_n_490__44_,r_n_490__43_,r_n_490__42_,
  r_n_490__41_,r_n_490__40_,r_n_490__39_,r_n_490__38_,r_n_490__37_,r_n_490__36_,
  r_n_490__35_,r_n_490__34_,r_n_490__33_,r_n_490__32_,r_n_490__31_,r_n_490__30_,
  r_n_490__29_,r_n_490__28_,r_n_490__27_,r_n_490__26_,r_n_490__25_,r_n_490__24_,
  r_n_490__23_,r_n_490__22_,r_n_490__21_,r_n_490__20_,r_n_490__19_,r_n_490__18_,
  r_n_490__17_,r_n_490__16_,r_n_490__15_,r_n_490__14_,r_n_490__13_,r_n_490__12_,
  r_n_490__11_,r_n_490__10_,r_n_490__9_,r_n_490__8_,r_n_490__7_,r_n_490__6_,r_n_490__5_,
  r_n_490__4_,r_n_490__3_,r_n_490__2_,r_n_490__1_,r_n_490__0_,r_n_489__63_,
  r_n_489__62_,r_n_489__61_,r_n_489__60_,r_n_489__59_,r_n_489__58_,r_n_489__57_,r_n_489__56_,
  r_n_489__55_,r_n_489__54_,r_n_489__53_,r_n_489__52_,r_n_489__51_,r_n_489__50_,
  r_n_489__49_,r_n_489__48_,r_n_489__47_,r_n_489__46_,r_n_489__45_,r_n_489__44_,
  r_n_489__43_,r_n_489__42_,r_n_489__41_,r_n_489__40_,r_n_489__39_,r_n_489__38_,
  r_n_489__37_,r_n_489__36_,r_n_489__35_,r_n_489__34_,r_n_489__33_,r_n_489__32_,
  r_n_489__31_,r_n_489__30_,r_n_489__29_,r_n_489__28_,r_n_489__27_,r_n_489__26_,
  r_n_489__25_,r_n_489__24_,r_n_489__23_,r_n_489__22_,r_n_489__21_,r_n_489__20_,
  r_n_489__19_,r_n_489__18_,r_n_489__17_,r_n_489__16_,r_n_489__15_,r_n_489__14_,r_n_489__13_,
  r_n_489__12_,r_n_489__11_,r_n_489__10_,r_n_489__9_,r_n_489__8_,r_n_489__7_,
  r_n_489__6_,r_n_489__5_,r_n_489__4_,r_n_489__3_,r_n_489__2_,r_n_489__1_,r_n_489__0_,
  r_n_504__63_,r_n_504__62_,r_n_504__61_,r_n_504__60_,r_n_504__59_,r_n_504__58_,
  r_n_504__57_,r_n_504__56_,r_n_504__55_,r_n_504__54_,r_n_504__53_,r_n_504__52_,
  r_n_504__51_,r_n_504__50_,r_n_504__49_,r_n_504__48_,r_n_504__47_,r_n_504__46_,
  r_n_504__45_,r_n_504__44_,r_n_504__43_,r_n_504__42_,r_n_504__41_,r_n_504__40_,
  r_n_504__39_,r_n_504__38_,r_n_504__37_,r_n_504__36_,r_n_504__35_,r_n_504__34_,
  r_n_504__33_,r_n_504__32_,r_n_504__31_,r_n_504__30_,r_n_504__29_,r_n_504__28_,r_n_504__27_,
  r_n_504__26_,r_n_504__25_,r_n_504__24_,r_n_504__23_,r_n_504__22_,r_n_504__21_,
  r_n_504__20_,r_n_504__19_,r_n_504__18_,r_n_504__17_,r_n_504__16_,r_n_504__15_,
  r_n_504__14_,r_n_504__13_,r_n_504__12_,r_n_504__11_,r_n_504__10_,r_n_504__9_,
  r_n_504__8_,r_n_504__7_,r_n_504__6_,r_n_504__5_,r_n_504__4_,r_n_504__3_,r_n_504__2_,
  r_n_504__1_,r_n_504__0_,r_n_503__63_,r_n_503__62_,r_n_503__61_,r_n_503__60_,
  r_n_503__59_,r_n_503__58_,r_n_503__57_,r_n_503__56_,r_n_503__55_,r_n_503__54_,
  r_n_503__53_,r_n_503__52_,r_n_503__51_,r_n_503__50_,r_n_503__49_,r_n_503__48_,
  r_n_503__47_,r_n_503__46_,r_n_503__45_,r_n_503__44_,r_n_503__43_,r_n_503__42_,r_n_503__41_,
  r_n_503__40_,r_n_503__39_,r_n_503__38_,r_n_503__37_,r_n_503__36_,r_n_503__35_,
  r_n_503__34_,r_n_503__33_,r_n_503__32_,r_n_503__31_,r_n_503__30_,r_n_503__29_,
  r_n_503__28_,r_n_503__27_,r_n_503__26_,r_n_503__25_,r_n_503__24_,r_n_503__23_,
  r_n_503__22_,r_n_503__21_,r_n_503__20_,r_n_503__19_,r_n_503__18_,r_n_503__17_,
  r_n_503__16_,r_n_503__15_,r_n_503__14_,r_n_503__13_,r_n_503__12_,r_n_503__11_,
  r_n_503__10_,r_n_503__9_,r_n_503__8_,r_n_503__7_,r_n_503__6_,r_n_503__5_,r_n_503__4_,
  r_n_503__3_,r_n_503__2_,r_n_503__1_,r_n_503__0_,r_n_502__63_,r_n_502__62_,
  r_n_502__61_,r_n_502__60_,r_n_502__59_,r_n_502__58_,r_n_502__57_,r_n_502__56_,r_n_502__55_,
  r_n_502__54_,r_n_502__53_,r_n_502__52_,r_n_502__51_,r_n_502__50_,r_n_502__49_,
  r_n_502__48_,r_n_502__47_,r_n_502__46_,r_n_502__45_,r_n_502__44_,r_n_502__43_,
  r_n_502__42_,r_n_502__41_,r_n_502__40_,r_n_502__39_,r_n_502__38_,r_n_502__37_,
  r_n_502__36_,r_n_502__35_,r_n_502__34_,r_n_502__33_,r_n_502__32_,r_n_502__31_,
  r_n_502__30_,r_n_502__29_,r_n_502__28_,r_n_502__27_,r_n_502__26_,r_n_502__25_,
  r_n_502__24_,r_n_502__23_,r_n_502__22_,r_n_502__21_,r_n_502__20_,r_n_502__19_,r_n_502__18_,
  r_n_502__17_,r_n_502__16_,r_n_502__15_,r_n_502__14_,r_n_502__13_,r_n_502__12_,
  r_n_502__11_,r_n_502__10_,r_n_502__9_,r_n_502__8_,r_n_502__7_,r_n_502__6_,
  r_n_502__5_,r_n_502__4_,r_n_502__3_,r_n_502__2_,r_n_502__1_,r_n_502__0_,r_n_501__63_,
  r_n_501__62_,r_n_501__61_,r_n_501__60_,r_n_501__59_,r_n_501__58_,r_n_501__57_,
  r_n_501__56_,r_n_501__55_,r_n_501__54_,r_n_501__53_,r_n_501__52_,r_n_501__51_,
  r_n_501__50_,r_n_501__49_,r_n_501__48_,r_n_501__47_,r_n_501__46_,r_n_501__45_,
  r_n_501__44_,r_n_501__43_,r_n_501__42_,r_n_501__41_,r_n_501__40_,r_n_501__39_,
  r_n_501__38_,r_n_501__37_,r_n_501__36_,r_n_501__35_,r_n_501__34_,r_n_501__33_,r_n_501__32_,
  r_n_501__31_,r_n_501__30_,r_n_501__29_,r_n_501__28_,r_n_501__27_,r_n_501__26_,
  r_n_501__25_,r_n_501__24_,r_n_501__23_,r_n_501__22_,r_n_501__21_,r_n_501__20_,
  r_n_501__19_,r_n_501__18_,r_n_501__17_,r_n_501__16_,r_n_501__15_,r_n_501__14_,
  r_n_501__13_,r_n_501__12_,r_n_501__11_,r_n_501__10_,r_n_501__9_,r_n_501__8_,
  r_n_501__7_,r_n_501__6_,r_n_501__5_,r_n_501__4_,r_n_501__3_,r_n_501__2_,r_n_501__1_,
  r_n_501__0_,r_n_500__63_,r_n_500__62_,r_n_500__61_,r_n_500__60_,r_n_500__59_,
  r_n_500__58_,r_n_500__57_,r_n_500__56_,r_n_500__55_,r_n_500__54_,r_n_500__53_,
  r_n_500__52_,r_n_500__51_,r_n_500__50_,r_n_500__49_,r_n_500__48_,r_n_500__47_,r_n_500__46_,
  r_n_500__45_,r_n_500__44_,r_n_500__43_,r_n_500__42_,r_n_500__41_,r_n_500__40_,
  r_n_500__39_,r_n_500__38_,r_n_500__37_,r_n_500__36_,r_n_500__35_,r_n_500__34_,
  r_n_500__33_,r_n_500__32_,r_n_500__31_,r_n_500__30_,r_n_500__29_,r_n_500__28_,
  r_n_500__27_,r_n_500__26_,r_n_500__25_,r_n_500__24_,r_n_500__23_,r_n_500__22_,
  r_n_500__21_,r_n_500__20_,r_n_500__19_,r_n_500__18_,r_n_500__17_,r_n_500__16_,
  r_n_500__15_,r_n_500__14_,r_n_500__13_,r_n_500__12_,r_n_500__11_,r_n_500__10_,r_n_500__9_,
  r_n_500__8_,r_n_500__7_,r_n_500__6_,r_n_500__5_,r_n_500__4_,r_n_500__3_,
  r_n_500__2_,r_n_500__1_,r_n_500__0_,r_n_499__63_,r_n_499__62_,r_n_499__61_,r_n_499__60_,
  r_n_499__59_,r_n_499__58_,r_n_499__57_,r_n_499__56_,r_n_499__55_,r_n_499__54_,
  r_n_499__53_,r_n_499__52_,r_n_499__51_,r_n_499__50_,r_n_499__49_,r_n_499__48_,
  r_n_499__47_,r_n_499__46_,r_n_499__45_,r_n_499__44_,r_n_499__43_,r_n_499__42_,
  r_n_499__41_,r_n_499__40_,r_n_499__39_,r_n_499__38_,r_n_499__37_,r_n_499__36_,
  r_n_499__35_,r_n_499__34_,r_n_499__33_,r_n_499__32_,r_n_499__31_,r_n_499__30_,
  r_n_499__29_,r_n_499__28_,r_n_499__27_,r_n_499__26_,r_n_499__25_,r_n_499__24_,
  r_n_499__23_,r_n_499__22_,r_n_499__21_,r_n_499__20_,r_n_499__19_,r_n_499__18_,r_n_499__17_,
  r_n_499__16_,r_n_499__15_,r_n_499__14_,r_n_499__13_,r_n_499__12_,r_n_499__11_,
  r_n_499__10_,r_n_499__9_,r_n_499__8_,r_n_499__7_,r_n_499__6_,r_n_499__5_,
  r_n_499__4_,r_n_499__3_,r_n_499__2_,r_n_499__1_,r_n_499__0_,r_n_498__63_,r_n_498__62_,
  r_n_498__61_,r_n_498__60_,r_n_498__59_,r_n_498__58_,r_n_498__57_,r_n_498__56_,
  r_n_498__55_,r_n_498__54_,r_n_498__53_,r_n_498__52_,r_n_498__51_,r_n_498__50_,
  r_n_498__49_,r_n_498__48_,r_n_498__47_,r_n_498__46_,r_n_498__45_,r_n_498__44_,
  r_n_498__43_,r_n_498__42_,r_n_498__41_,r_n_498__40_,r_n_498__39_,r_n_498__38_,
  r_n_498__37_,r_n_498__36_,r_n_498__35_,r_n_498__34_,r_n_498__33_,r_n_498__32_,r_n_498__31_,
  r_n_498__30_,r_n_498__29_,r_n_498__28_,r_n_498__27_,r_n_498__26_,r_n_498__25_,
  r_n_498__24_,r_n_498__23_,r_n_498__22_,r_n_498__21_,r_n_498__20_,r_n_498__19_,
  r_n_498__18_,r_n_498__17_,r_n_498__16_,r_n_498__15_,r_n_498__14_,r_n_498__13_,
  r_n_498__12_,r_n_498__11_,r_n_498__10_,r_n_498__9_,r_n_498__8_,r_n_498__7_,r_n_498__6_,
  r_n_498__5_,r_n_498__4_,r_n_498__3_,r_n_498__2_,r_n_498__1_,r_n_498__0_,
  r_n_497__63_,r_n_497__62_,r_n_497__61_,r_n_497__60_,r_n_497__59_,r_n_497__58_,
  r_n_497__57_,r_n_497__56_,r_n_497__55_,r_n_497__54_,r_n_497__53_,r_n_497__52_,
  r_n_497__51_,r_n_497__50_,r_n_497__49_,r_n_497__48_,r_n_497__47_,r_n_497__46_,r_n_497__45_,
  r_n_497__44_,r_n_497__43_,r_n_497__42_,r_n_497__41_,r_n_497__40_,r_n_497__39_,
  r_n_497__38_,r_n_497__37_,r_n_497__36_,r_n_497__35_,r_n_497__34_,r_n_497__33_,
  r_n_497__32_,r_n_497__31_,r_n_497__30_,r_n_497__29_,r_n_497__28_,r_n_497__27_,
  r_n_497__26_,r_n_497__25_,r_n_497__24_,r_n_497__23_,r_n_497__22_,r_n_497__21_,
  r_n_497__20_,r_n_497__19_,r_n_497__18_,r_n_497__17_,r_n_497__16_,r_n_497__15_,
  r_n_497__14_,r_n_497__13_,r_n_497__12_,r_n_497__11_,r_n_497__10_,r_n_497__9_,r_n_497__8_,
  r_n_497__7_,r_n_497__6_,r_n_497__5_,r_n_497__4_,r_n_497__3_,r_n_497__2_,
  r_n_497__1_,r_n_497__0_,r_n_511__63_,r_n_511__62_,r_n_511__61_,r_n_511__60_,r_n_511__59_,
  r_n_511__58_,r_n_511__57_,r_n_511__56_,r_n_511__55_,r_n_511__54_,r_n_511__53_,
  r_n_511__52_,r_n_511__51_,r_n_511__50_,r_n_511__49_,r_n_511__48_,r_n_511__47_,
  r_n_511__46_,r_n_511__45_,r_n_511__44_,r_n_511__43_,r_n_511__42_,r_n_511__41_,
  r_n_511__40_,r_n_511__39_,r_n_511__38_,r_n_511__37_,r_n_511__36_,r_n_511__35_,
  r_n_511__34_,r_n_511__33_,r_n_511__32_,r_n_511__31_,r_n_511__30_,r_n_511__29_,
  r_n_511__28_,r_n_511__27_,r_n_511__26_,r_n_511__25_,r_n_511__24_,r_n_511__23_,r_n_511__22_,
  r_n_511__21_,r_n_511__20_,r_n_511__19_,r_n_511__18_,r_n_511__17_,r_n_511__16_,
  r_n_511__15_,r_n_511__14_,r_n_511__13_,r_n_511__12_,r_n_511__11_,r_n_511__10_,
  r_n_511__9_,r_n_511__8_,r_n_511__7_,r_n_511__6_,r_n_511__5_,r_n_511__4_,r_n_511__3_,
  r_n_511__2_,r_n_511__1_,r_n_511__0_,r_n_510__63_,r_n_510__62_,r_n_510__61_,
  r_n_510__60_,r_n_510__59_,r_n_510__58_,r_n_510__57_,r_n_510__56_,r_n_510__55_,
  r_n_510__54_,r_n_510__53_,r_n_510__52_,r_n_510__51_,r_n_510__50_,r_n_510__49_,
  r_n_510__48_,r_n_510__47_,r_n_510__46_,r_n_510__45_,r_n_510__44_,r_n_510__43_,
  r_n_510__42_,r_n_510__41_,r_n_510__40_,r_n_510__39_,r_n_510__38_,r_n_510__37_,r_n_510__36_,
  r_n_510__35_,r_n_510__34_,r_n_510__33_,r_n_510__32_,r_n_510__31_,r_n_510__30_,
  r_n_510__29_,r_n_510__28_,r_n_510__27_,r_n_510__26_,r_n_510__25_,r_n_510__24_,
  r_n_510__23_,r_n_510__22_,r_n_510__21_,r_n_510__20_,r_n_510__19_,r_n_510__18_,
  r_n_510__17_,r_n_510__16_,r_n_510__15_,r_n_510__14_,r_n_510__13_,r_n_510__12_,
  r_n_510__11_,r_n_510__10_,r_n_510__9_,r_n_510__8_,r_n_510__7_,r_n_510__6_,r_n_510__5_,
  r_n_510__4_,r_n_510__3_,r_n_510__2_,r_n_510__1_,r_n_510__0_,r_n_509__63_,
  r_n_509__62_,r_n_509__61_,r_n_509__60_,r_n_509__59_,r_n_509__58_,r_n_509__57_,
  r_n_509__56_,r_n_509__55_,r_n_509__54_,r_n_509__53_,r_n_509__52_,r_n_509__51_,r_n_509__50_,
  r_n_509__49_,r_n_509__48_,r_n_509__47_,r_n_509__46_,r_n_509__45_,r_n_509__44_,
  r_n_509__43_,r_n_509__42_,r_n_509__41_,r_n_509__40_,r_n_509__39_,r_n_509__38_,
  r_n_509__37_,r_n_509__36_,r_n_509__35_,r_n_509__34_,r_n_509__33_,r_n_509__32_,
  r_n_509__31_,r_n_509__30_,r_n_509__29_,r_n_509__28_,r_n_509__27_,r_n_509__26_,
  r_n_509__25_,r_n_509__24_,r_n_509__23_,r_n_509__22_,r_n_509__21_,r_n_509__20_,
  r_n_509__19_,r_n_509__18_,r_n_509__17_,r_n_509__16_,r_n_509__15_,r_n_509__14_,
  r_n_509__13_,r_n_509__12_,r_n_509__11_,r_n_509__10_,r_n_509__9_,r_n_509__8_,r_n_509__7_,
  r_n_509__6_,r_n_509__5_,r_n_509__4_,r_n_509__3_,r_n_509__2_,r_n_509__1_,r_n_509__0_,
  r_n_508__63_,r_n_508__62_,r_n_508__61_,r_n_508__60_,r_n_508__59_,r_n_508__58_,
  r_n_508__57_,r_n_508__56_,r_n_508__55_,r_n_508__54_,r_n_508__53_,r_n_508__52_,
  r_n_508__51_,r_n_508__50_,r_n_508__49_,r_n_508__48_,r_n_508__47_,r_n_508__46_,
  r_n_508__45_,r_n_508__44_,r_n_508__43_,r_n_508__42_,r_n_508__41_,r_n_508__40_,
  r_n_508__39_,r_n_508__38_,r_n_508__37_,r_n_508__36_,r_n_508__35_,r_n_508__34_,
  r_n_508__33_,r_n_508__32_,r_n_508__31_,r_n_508__30_,r_n_508__29_,r_n_508__28_,
  r_n_508__27_,r_n_508__26_,r_n_508__25_,r_n_508__24_,r_n_508__23_,r_n_508__22_,r_n_508__21_,
  r_n_508__20_,r_n_508__19_,r_n_508__18_,r_n_508__17_,r_n_508__16_,r_n_508__15_,
  r_n_508__14_,r_n_508__13_,r_n_508__12_,r_n_508__11_,r_n_508__10_,r_n_508__9_,
  r_n_508__8_,r_n_508__7_,r_n_508__6_,r_n_508__5_,r_n_508__4_,r_n_508__3_,r_n_508__2_,
  r_n_508__1_,r_n_508__0_,r_n_507__63_,r_n_507__62_,r_n_507__61_,r_n_507__60_,
  r_n_507__59_,r_n_507__58_,r_n_507__57_,r_n_507__56_,r_n_507__55_,r_n_507__54_,
  r_n_507__53_,r_n_507__52_,r_n_507__51_,r_n_507__50_,r_n_507__49_,r_n_507__48_,
  r_n_507__47_,r_n_507__46_,r_n_507__45_,r_n_507__44_,r_n_507__43_,r_n_507__42_,
  r_n_507__41_,r_n_507__40_,r_n_507__39_,r_n_507__38_,r_n_507__37_,r_n_507__36_,r_n_507__35_,
  r_n_507__34_,r_n_507__33_,r_n_507__32_,r_n_507__31_,r_n_507__30_,r_n_507__29_,
  r_n_507__28_,r_n_507__27_,r_n_507__26_,r_n_507__25_,r_n_507__24_,r_n_507__23_,
  r_n_507__22_,r_n_507__21_,r_n_507__20_,r_n_507__19_,r_n_507__18_,r_n_507__17_,
  r_n_507__16_,r_n_507__15_,r_n_507__14_,r_n_507__13_,r_n_507__12_,r_n_507__11_,
  r_n_507__10_,r_n_507__9_,r_n_507__8_,r_n_507__7_,r_n_507__6_,r_n_507__5_,r_n_507__4_,
  r_n_507__3_,r_n_507__2_,r_n_507__1_,r_n_507__0_,r_n_506__63_,r_n_506__62_,
  r_n_506__61_,r_n_506__60_,r_n_506__59_,r_n_506__58_,r_n_506__57_,r_n_506__56_,
  r_n_506__55_,r_n_506__54_,r_n_506__53_,r_n_506__52_,r_n_506__51_,r_n_506__50_,r_n_506__49_,
  r_n_506__48_,r_n_506__47_,r_n_506__46_,r_n_506__45_,r_n_506__44_,r_n_506__43_,
  r_n_506__42_,r_n_506__41_,r_n_506__40_,r_n_506__39_,r_n_506__38_,r_n_506__37_,
  r_n_506__36_,r_n_506__35_,r_n_506__34_,r_n_506__33_,r_n_506__32_,r_n_506__31_,
  r_n_506__30_,r_n_506__29_,r_n_506__28_,r_n_506__27_,r_n_506__26_,r_n_506__25_,
  r_n_506__24_,r_n_506__23_,r_n_506__22_,r_n_506__21_,r_n_506__20_,r_n_506__19_,
  r_n_506__18_,r_n_506__17_,r_n_506__16_,r_n_506__15_,r_n_506__14_,r_n_506__13_,r_n_506__12_,
  r_n_506__11_,r_n_506__10_,r_n_506__9_,r_n_506__8_,r_n_506__7_,r_n_506__6_,
  r_n_506__5_,r_n_506__4_,r_n_506__3_,r_n_506__2_,r_n_506__1_,r_n_506__0_,r_n_505__63_,
  r_n_505__62_,r_n_505__61_,r_n_505__60_,r_n_505__59_,r_n_505__58_,r_n_505__57_,
  r_n_505__56_,r_n_505__55_,r_n_505__54_,r_n_505__53_,r_n_505__52_,r_n_505__51_,
  r_n_505__50_,r_n_505__49_,r_n_505__48_,r_n_505__47_,r_n_505__46_,r_n_505__45_,
  r_n_505__44_,r_n_505__43_,r_n_505__42_,r_n_505__41_,r_n_505__40_,r_n_505__39_,
  r_n_505__38_,r_n_505__37_,r_n_505__36_,r_n_505__35_,r_n_505__34_,r_n_505__33_,
  r_n_505__32_,r_n_505__31_,r_n_505__30_,r_n_505__29_,r_n_505__28_,r_n_505__27_,r_n_505__26_,
  r_n_505__25_,r_n_505__24_,r_n_505__23_,r_n_505__22_,r_n_505__21_,r_n_505__20_,
  r_n_505__19_,r_n_505__18_,r_n_505__17_,r_n_505__16_,r_n_505__15_,r_n_505__14_,
  r_n_505__13_,r_n_505__12_,r_n_505__11_,r_n_505__10_,r_n_505__9_,r_n_505__8_,
  r_n_505__7_,r_n_505__6_,r_n_505__5_,r_n_505__4_,r_n_505__3_,r_n_505__2_,r_n_505__1_,
  r_n_505__0_,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,
  N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,
  N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,
  N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,
  N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,
  N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,
  N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,
  N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,
  N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,
  N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,
  N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1173,
  N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,
  N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,
  N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,
  N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,
  N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,
  N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,
  N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,
  N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,
  N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,
  N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,
  N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320,
  N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,
  N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,
  N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,
  N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,
  N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,
  N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,
  N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,
  N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,
  N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,
  N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,
  N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,
  N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,
  N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,
  N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,
  N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,
  N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,
  N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,
  N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,
  N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,
  N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,
  N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,
  N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613,
  N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626,
  N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,N1638,N1639,N1640,
  N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,N1651,N1652,N1653,
  N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,N1665,N1666,
  N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680,
  N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693,
  N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,
  N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720,
  N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,N1731,N1732,N1733,
  N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,N1745,N1746,
  N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,N1758,N1759,N1760,
  N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,N1771,N1772,N1773,
  N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,N1785,N1786,
  N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1800,
  N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,N1811,N1812,N1813,
  N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,N1825,N1826,
  N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,N1838,N1839,N1840,
  N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,N1851,N1852,N1853,
  N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,N1865,N1866,
  N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,
  N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,N1891,N1892,N1893,
  N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,N1905,N1906,
  N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918,N1919,N1920,
  N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,
  N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,
  N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,N1958,N1959,N1960,
  N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,
  N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,N1985,N1986,
  N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,N1998,N1999,N2000,
  N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,N2011,N2012,N2013,
  N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,N2025,N2026,
  N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,N2038,N2039,N2040,
  N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,N2051,N2052,N2053,
  N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066,
  N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,N2078,N2079,N2080,
  N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,N2091,N2092,N2093,
  N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,N2105,N2106,
  N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,N2118,N2119,N2120,
  N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,N2131,N2132,N2133,
  N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144,N2145,N2146,
  N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,N2158,N2159,N2160,
  N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,N2170,N2171,N2172,N2173,
  N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,N2184,N2185,N2186,
  N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197,N2198,N2199,N2200,
  N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,N2210,N2211,N2212,N2213,
  N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,N2224,N2225,N2226,
  N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2238,N2239,N2240,
  N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,N2251,N2252,N2253,
  N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,N2264,N2265,N2266,
  N2267,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,N2278,N2279,N2280,
  N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290,N2291,N2292,N2293,
  N2294,N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302,N2303,N2304,N2305,N2306,
  N2307,N2308,N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,N2318,N2319,N2320,
  N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,N2331,N2332,N2333,
  N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,
  N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,N2358,N2359,N2360,
  N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2369,N2370,N2371,N2372,N2373,
  N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382,N2383,N2384,N2385,N2386,
  N2387,N2388,N2389,N2390,N2391,N2392,N2393,N2394,N2395,N2396,N2397,N2398,N2399,N2400,
  N2401,N2402,N2403,N2404,N2405,N2406,N2407,N2408,N2409,N2410,N2411,N2412,N2413,
  N2414,N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422,N2423,N2424,N2425,N2426,
  N2427,N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,N2438,N2439,N2440,
  N2441,N2442,N2443,N2444,N2445,N2446,N2447,N2448,N2449,N2450,N2451,N2452,N2453,
  N2454,N2455,N2456,N2457,N2458,N2459,N2460,N2461,N2462,N2463,N2464,N2465,N2466,
  N2467,N2468,N2469,N2470,N2471,N2472,N2473,N2474,N2475,N2476,N2477,N2478,N2479,N2480,
  N2481,N2482,N2483,N2484,N2485,N2486,N2487,N2488,N2489,N2490,N2491,N2492,N2493,
  N2494,N2495,N2496,N2497,N2498,N2499,N2500,N2501,N2502,N2503,N2504,N2505,N2506,
  N2507,N2508,N2509,N2510,N2511,N2512,N2513,N2514,N2515,N2516,N2517,N2518,N2519,N2520,
  N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528,N2529,N2530,N2531,N2532,N2533,
  N2534,N2535,N2536,N2537,N2538,N2539,N2540,N2541,N2542,N2543,N2544,N2545,N2546,
  N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2554,N2555,N2556,N2557,N2558,N2559,N2560,
  N2561,N2562,N2563,N2564,N2565,N2566,N2567,N2568,N2569,N2570,N2571,N2572,N2573,
  N2574,N2575,N2576,N2577,N2578,N2579,N2580,N2581,N2582,N2583,N2584,N2585,N2586,
  N2587,N2588,N2589,N2590,N2591,N2592,N2593,N2594,N2595,N2596,N2597,N2598,N2599,N2600,
  N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,N2609,N2610,N2611,N2612,N2613,
  N2614,N2615,N2616,N2617,N2618,N2619,N2620,N2621,N2622,N2623,N2624,N2625,N2626,
  N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2637,N2638,N2639,N2640,
  N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,N2649,N2650,N2651,N2652,N2653,
  N2654,N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662,N2663,N2664,N2665,N2666,
  N2667,N2668,N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,N2678,N2679,N2680,
  N2681,N2682,N2683,N2684,N2685,N2686,N2687,N2688,N2689,N2690,N2691,N2692,N2693,
  N2694,N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2704,N2705,N2706,
  N2707,N2708,N2709,N2710,N2711,N2712,N2713,N2714,N2715,N2716,N2717,N2718,N2719,N2720,
  N2721,N2722,N2723,N2724,N2725,N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,
  N2734,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,
  N2747,N2748,N2749,N2750,N2751,N2752,N2753,N2754,N2755,N2756,N2757,N2758,N2759,N2760,
  N2761,N2762,N2763,N2764,N2765,N2766,N2767,N2768,N2769,N2770,N2771,N2772,N2773,
  N2774,N2775,N2776,N2777,N2778,N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,
  N2787,N2788,N2789,N2790,N2791,N2792,N2793,N2794,N2795,N2796,N2797,N2798,N2799,N2800,
  N2801,N2802,N2803,N2804,N2805,N2806,N2807,N2808,N2809,N2810,N2811,N2812,N2813,
  N2814,N2815,N2816,N2817,N2818,N2819,N2820,N2821,N2822,N2823,N2824,N2825,N2826,
  N2827,N2828,N2829,N2830,N2831,N2832,N2833,N2834,N2835,N2836,N2837,N2838,N2839,N2840,
  N2841,N2842,N2843,N2844,N2845,N2846,N2847,N2848,N2849,N2850,N2851,N2852,N2853,
  N2854,N2855,N2856,N2857,N2858,N2859,N2860,N2861,N2862,N2863,N2864,N2865,N2866,
  N2867,N2868,N2869,N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,
  N2881,N2882,N2883,N2884,N2885,N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2893,
  N2894,N2895,N2896,N2897,N2898,N2899,N2900,N2901,N2902,N2903,N2904,N2905,N2906,
  N2907,N2908,N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,N2917,N2918,N2919,N2920,
  N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,N2930,N2931,N2932,N2933,
  N2934,N2935,N2936,N2937,N2938,N2939,N2940,N2941,N2942,N2943,N2944,N2945,N2946,
  N2947,N2948,N2949,N2950,N2951,N2952,N2953,N2954,N2955,N2956,N2957,N2958,N2959,N2960,
  N2961,N2962,N2963,N2964,N2965,N2966,N2967,N2968,N2969,N2970,N2971,N2972,N2973,
  N2974,N2975,N2976,N2977,N2978,N2979,N2980,N2981,N2982,N2983,N2984,N2985,N2986,
  N2987,N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,
  N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,N3010,N3011,N3012,N3013,
  N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022,N3023,N3024,N3025,N3026,
  N3027,N3028,N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,
  N3041,N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,N3050,N3051,N3052,N3053,
  N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3062,N3063,N3064,N3065,N3066,
  N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,N3076,N3077,N3078,N3079,N3080,
  N3081,N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,N3090,N3091,N3092,N3093,
  N3094,N3095,N3096,N3097,N3098,N3099,N3100,N3101,N3102,N3103,N3104,N3105,N3106,
  N3107,N3108,N3109,N3110,N3111,N3112,N3113,N3114,N3115,N3116,N3117,N3118,N3119,N3120,
  N3121,N3122,N3123,N3124,N3125,N3126,N3127,N3128,N3129,N3130,N3131,N3132,N3133,
  N3134,N3135,N3136,N3137,N3138,N3139,N3140,N3141,N3142,N3143,N3144,N3145,N3146,
  N3147,N3148,N3149,N3150,N3151,N3152,N3153,N3154,N3155,N3156,N3157,N3158,N3159,N3160,
  N3161,N3162,N3163,N3164,N3165,N3166,N3167,N3168,N3169,N3170,N3171,N3172,N3173,
  N3174,N3175,N3176,N3177,N3178,N3179,N3180,N3181,N3182,N3183,N3184,N3185,N3186,
  N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194,N3195,N3196,N3197,N3198,N3199,N3200,
  N3201,N3202,N3203,N3204,N3205,N3206,N3207,N3208,N3209,N3210,N3211,N3212,N3213,
  N3214,N3215,N3216,N3217,N3218,N3219,N3220,N3221,N3222,N3223,N3224,N3225,N3226,
  N3227,N3228,N3229,N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,N3238,N3239,N3240,
  N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,N3249,N3250,N3251,N3252,N3253,
  N3254,N3255,N3256,N3257,N3258,N3259,N3260,N3261,N3262,N3263,N3264,N3265,N3266,
  N3267,N3268,N3269,N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,N3278,N3279,N3280,
  N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,N3290,N3291,N3292,N3293,
  N3294,N3295,N3296,N3297,N3298,N3299,N3300,N3301,N3302,N3303,N3304,N3305,N3306,
  N3307,N3308,N3309,N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,N3318,N3319,N3320,
  N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,N3330,N3331,N3332,N3333,
  N3334,N3335,N3336,N3337,N3338,N3339,N3340,N3341,N3342,N3343,N3344,N3345,N3346,
  N3347,N3348,N3349,N3350,N3351,N3352,N3353,N3354,N3355,N3356,N3357,N3358,N3359,N3360,
  N3361,N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,N3370,N3371,N3372,N3373,
  N3374,N3375,N3376,N3377,N3378,N3379,N3380,N3381,N3382,N3383,N3384,N3385,N3386,
  N3387,N3388,N3389,N3390,N3391,N3392,N3393,N3394,N3395,N3396,N3397,N3398,N3399,N3400,
  N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3408,N3409,N3410,N3411,N3412,N3413,
  N3414,N3415,N3416,N3417,N3418,N3419,N3420,N3421,N3422,N3423,N3424,N3425,N3426,
  N3427,N3428,N3429,N3430,N3431,N3432,N3433,N3434,N3435,N3436,N3437,N3438,N3439,N3440,
  N3441,N3442,N3443,N3444,N3445,N3446,N3447,N3448,N3449,N3450,N3451,N3452,N3453,
  N3454,N3455,N3456,N3457,N3458,N3459,N3460,N3461,N3462,N3463,N3464,N3465,N3466,
  N3467,N3468,N3469,N3470,N3471,N3472,N3473,N3474,N3475,N3476,N3477,N3478,N3479,N3480,
  N3481,N3482,N3483,N3484,N3485,N3486,N3487,N3488,N3489,N3490,N3491,N3492,N3493,
  N3494,N3495,N3496,N3497,N3498,N3499,N3500,N3501,N3502,N3503,N3504,N3505,N3506,
  N3507,N3508,N3509,N3510,N3511,N3512,N3513,N3514,N3515,N3516,N3517,N3518,N3519,N3520,
  N3521,N3522,N3523,N3524,N3525,N3526,N3527,N3528,N3529,N3530,N3531,N3532,N3533,
  N3534,N3535,N3536,N3537,N3538,N3539,N3540,N3541,N3542,N3543,N3544,N3545,N3546,
  N3547,N3548,N3549,N3550,N3551,N3552,N3553,N3554,N3555,N3556,N3557,N3558,N3559,N3560,
  N3561,N3562,N3563,N3564,N3565,N3566,N3567,N3568,N3569,N3570,N3571,N3572,N3573,
  N3574,N3575,N3576,N3577,N3578,N3579,N3580,N3581,N3582,N3583,N3584,N3585,N3586,
  N3587,N3588,N3589,N3590,N3591,N3592,N3593,N3594,N3595,N3596,N3597,N3598,N3599,N3600,
  N3601,N3602,N3603,N3604,N3605,N3606,N3607,N3608,N3609,N3610,N3611,N3612,N3613,
  N3614,N3615,N3616,N3617,N3618,N3619,N3620,N3621,N3622,N3623,N3624,N3625,N3626,
  N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3636,N3637,N3638,N3639,N3640,
  N3641,N3642,N3643,N3644,N3645,N3646,N3647,N3648,N3649,N3650,N3651,N3652,N3653,
  N3654,N3655,N3656,N3657,N3658,N3659,N3660,N3661,N3662,N3663,N3664,N3665,N3666,
  N3667,N3668,N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3676,N3677,N3678,N3679,N3680,
  N3681,N3682,N3683,N3684,N3685,N3686,N3687,N3688,N3689,N3690,N3691,N3692,N3693,
  N3694,N3695,N3696,N3697,N3698,N3699,N3700,N3701,N3702,N3703,N3704,N3705,N3706,
  N3707,N3708,N3709,N3710,N3711,N3712,N3713,N3714,N3715,N3716,N3717,N3718,N3719,N3720,
  N3721,N3722,N3723,N3724,N3725,N3726,N3727,N3728,N3729,N3730,N3731,N3732,N3733,
  N3734,N3735,N3736,N3737,N3738,N3739,N3740,N3741,N3742,N3743,N3744,N3745,N3746,
  N3747,N3748,N3749,N3750,N3751,N3752,N3753,N3754,N3755,N3756,N3757,N3758,N3759,N3760,
  N3761,N3762,N3763,N3764,N3765,N3766,N3767,N3768,N3769,N3770,N3771,N3772,N3773,
  N3774,N3775,N3776,N3777,N3778,N3779,N3780,N3781,N3782,N3783,N3784,N3785,N3786,
  N3787,N3788,N3789,N3790,N3791,N3792,N3793,N3794,N3795,N3796,N3797,N3798,N3799,N3800,
  N3801,N3802,N3803,N3804,N3805,N3806,N3807,N3808,N3809,N3810,N3811,N3812,N3813,
  N3814,N3815,N3816,N3817,N3818,N3819,N3820,N3821,N3822,N3823,N3824,N3825,N3826,
  N3827,N3828,N3829,N3830,N3831,N3832,N3833,N3834,N3835,N3836,N3837,N3838,N3839,N3840,
  N3841,N3842,N3843,N3844,N3845,N3846,N3847,N3848,N3849,N3850,N3851,N3852,N3853,
  N3854,N3855,N3856,N3857,N3858,N3859,N3860,N3861,N3862,N3863,N3864,N3865,N3866,
  N3867,N3868,N3869,N3870,N3871,N3872,N3873,N3874,N3875,N3876,N3877,N3878,N3879,N3880,
  N3881,N3882,N3883,N3884,N3885,N3886,N3887,N3888,N3889,N3890,N3891,N3892,N3893,
  N3894,N3895,N3896,N3897,N3898,N3899,N3900,N3901,N3902,N3903,N3904,N3905,N3906,
  N3907,N3908,N3909,N3910,N3911,N3912,N3913,N3914,N3915,N3916,N3917,N3918,N3919,N3920,
  N3921,N3922,N3923,N3924,N3925,N3926,N3927,N3928,N3929,N3930,N3931,N3932,N3933,
  N3934,N3935,N3936,N3937,N3938,N3939,N3940,N3941,N3942,N3943,N3944,N3945,N3946,
  N3947,N3948,N3949,N3950,N3951,N3952,N3953,N3954,N3955,N3956,N3957,N3958,N3959,N3960,
  N3961,N3962,N3963,N3964,N3965,N3966,N3967,N3968,N3969,N3970,N3971,N3972,N3973,
  N3974,N3975,N3976,N3977,N3978,N3979,N3980,N3981,N3982,N3983,N3984,N3985,N3986,
  N3987,N3988,N3989,N3990,N3991,N3992,N3993,N3994,N3995,N3996,N3997,N3998,N3999,N4000,
  N4001,N4002,N4003,N4004,N4005,N4006,N4007,N4008,N4009,N4010,N4011,N4012,N4013,
  N4014,N4015,N4016,N4017,N4018,N4019,N4020,N4021,N4022,N4023,N4024,N4025,N4026,
  N4027,N4028,N4029,N4030,N4031,N4032,N4033,N4034,N4035,N4036,N4037,N4038,N4039,N4040,
  N4041,N4042,N4043,N4044,N4045,N4046,N4047,N4048,N4049,N4050,N4051,N4052,N4053,
  N4054,N4055,N4056,N4057,N4058,N4059,N4060,N4061,N4062,N4063,N4064,N4065,N4066,
  N4067,N4068,N4069,N4070,N4071,N4072,N4073,N4074,N4075,N4076,N4077,N4078,N4079,N4080,
  N4081,N4082,N4083,N4084,N4085,N4086,N4087,N4088,N4089,N4090,N4091,N4092,N4093,
  N4094,N4095;
  reg [63:0] data_o;
  reg r_1__63_,r_1__62_,r_1__61_,r_1__60_,r_1__59_,r_1__58_,r_1__57_,r_1__56_,
  r_1__55_,r_1__54_,r_1__53_,r_1__52_,r_1__51_,r_1__50_,r_1__49_,r_1__48_,r_1__47_,
  r_1__46_,r_1__45_,r_1__44_,r_1__43_,r_1__42_,r_1__41_,r_1__40_,r_1__39_,r_1__38_,
  r_1__37_,r_1__36_,r_1__35_,r_1__34_,r_1__33_,r_1__32_,r_1__31_,r_1__30_,r_1__29_,
  r_1__28_,r_1__27_,r_1__26_,r_1__25_,r_1__24_,r_1__23_,r_1__22_,r_1__21_,r_1__20_,
  r_1__19_,r_1__18_,r_1__17_,r_1__16_,r_1__15_,r_1__14_,r_1__13_,r_1__12_,r_1__11_,
  r_1__10_,r_1__9_,r_1__8_,r_1__7_,r_1__6_,r_1__5_,r_1__4_,r_1__3_,r_1__2_,r_1__1_,
  r_1__0_,r_2__63_,r_2__62_,r_2__61_,r_2__60_,r_2__59_,r_2__58_,r_2__57_,r_2__56_,
  r_2__55_,r_2__54_,r_2__53_,r_2__52_,r_2__51_,r_2__50_,r_2__49_,r_2__48_,r_2__47_,
  r_2__46_,r_2__45_,r_2__44_,r_2__43_,r_2__42_,r_2__41_,r_2__40_,r_2__39_,r_2__38_,
  r_2__37_,r_2__36_,r_2__35_,r_2__34_,r_2__33_,r_2__32_,r_2__31_,r_2__30_,
  r_2__29_,r_2__28_,r_2__27_,r_2__26_,r_2__25_,r_2__24_,r_2__23_,r_2__22_,r_2__21_,
  r_2__20_,r_2__19_,r_2__18_,r_2__17_,r_2__16_,r_2__15_,r_2__14_,r_2__13_,r_2__12_,
  r_2__11_,r_2__10_,r_2__9_,r_2__8_,r_2__7_,r_2__6_,r_2__5_,r_2__4_,r_2__3_,r_2__2_,
  r_2__1_,r_2__0_,r_3__63_,r_3__62_,r_3__61_,r_3__60_,r_3__59_,r_3__58_,r_3__57_,
  r_3__56_,r_3__55_,r_3__54_,r_3__53_,r_3__52_,r_3__51_,r_3__50_,r_3__49_,r_3__48_,
  r_3__47_,r_3__46_,r_3__45_,r_3__44_,r_3__43_,r_3__42_,r_3__41_,r_3__40_,r_3__39_,
  r_3__38_,r_3__37_,r_3__36_,r_3__35_,r_3__34_,r_3__33_,r_3__32_,r_3__31_,r_3__30_,
  r_3__29_,r_3__28_,r_3__27_,r_3__26_,r_3__25_,r_3__24_,r_3__23_,r_3__22_,r_3__21_,
  r_3__20_,r_3__19_,r_3__18_,r_3__17_,r_3__16_,r_3__15_,r_3__14_,r_3__13_,r_3__12_,
  r_3__11_,r_3__10_,r_3__9_,r_3__8_,r_3__7_,r_3__6_,r_3__5_,r_3__4_,r_3__3_,
  r_3__2_,r_3__1_,r_3__0_,r_4__63_,r_4__62_,r_4__61_,r_4__60_,r_4__59_,r_4__58_,
  r_4__57_,r_4__56_,r_4__55_,r_4__54_,r_4__53_,r_4__52_,r_4__51_,r_4__50_,r_4__49_,
  r_4__48_,r_4__47_,r_4__46_,r_4__45_,r_4__44_,r_4__43_,r_4__42_,r_4__41_,r_4__40_,
  r_4__39_,r_4__38_,r_4__37_,r_4__36_,r_4__35_,r_4__34_,r_4__33_,r_4__32_,r_4__31_,
  r_4__30_,r_4__29_,r_4__28_,r_4__27_,r_4__26_,r_4__25_,r_4__24_,r_4__23_,r_4__22_,
  r_4__21_,r_4__20_,r_4__19_,r_4__18_,r_4__17_,r_4__16_,r_4__15_,r_4__14_,r_4__13_,
  r_4__12_,r_4__11_,r_4__10_,r_4__9_,r_4__8_,r_4__7_,r_4__6_,r_4__5_,r_4__4_,r_4__3_,
  r_4__2_,r_4__1_,r_4__0_,r_5__63_,r_5__62_,r_5__61_,r_5__60_,r_5__59_,r_5__58_,
  r_5__57_,r_5__56_,r_5__55_,r_5__54_,r_5__53_,r_5__52_,r_5__51_,r_5__50_,r_5__49_,
  r_5__48_,r_5__47_,r_5__46_,r_5__45_,r_5__44_,r_5__43_,r_5__42_,r_5__41_,r_5__40_,
  r_5__39_,r_5__38_,r_5__37_,r_5__36_,r_5__35_,r_5__34_,r_5__33_,r_5__32_,
  r_5__31_,r_5__30_,r_5__29_,r_5__28_,r_5__27_,r_5__26_,r_5__25_,r_5__24_,r_5__23_,
  r_5__22_,r_5__21_,r_5__20_,r_5__19_,r_5__18_,r_5__17_,r_5__16_,r_5__15_,r_5__14_,
  r_5__13_,r_5__12_,r_5__11_,r_5__10_,r_5__9_,r_5__8_,r_5__7_,r_5__6_,r_5__5_,r_5__4_,
  r_5__3_,r_5__2_,r_5__1_,r_5__0_,r_6__63_,r_6__62_,r_6__61_,r_6__60_,r_6__59_,
  r_6__58_,r_6__57_,r_6__56_,r_6__55_,r_6__54_,r_6__53_,r_6__52_,r_6__51_,r_6__50_,
  r_6__49_,r_6__48_,r_6__47_,r_6__46_,r_6__45_,r_6__44_,r_6__43_,r_6__42_,r_6__41_,
  r_6__40_,r_6__39_,r_6__38_,r_6__37_,r_6__36_,r_6__35_,r_6__34_,r_6__33_,r_6__32_,
  r_6__31_,r_6__30_,r_6__29_,r_6__28_,r_6__27_,r_6__26_,r_6__25_,r_6__24_,r_6__23_,
  r_6__22_,r_6__21_,r_6__20_,r_6__19_,r_6__18_,r_6__17_,r_6__16_,r_6__15_,r_6__14_,
  r_6__13_,r_6__12_,r_6__11_,r_6__10_,r_6__9_,r_6__8_,r_6__7_,r_6__6_,r_6__5_,
  r_6__4_,r_6__3_,r_6__2_,r_6__1_,r_6__0_,r_7__63_,r_7__62_,r_7__61_,r_7__60_,
  r_7__59_,r_7__58_,r_7__57_,r_7__56_,r_7__55_,r_7__54_,r_7__53_,r_7__52_,r_7__51_,
  r_7__50_,r_7__49_,r_7__48_,r_7__47_,r_7__46_,r_7__45_,r_7__44_,r_7__43_,r_7__42_,
  r_7__41_,r_7__40_,r_7__39_,r_7__38_,r_7__37_,r_7__36_,r_7__35_,r_7__34_,r_7__33_,
  r_7__32_,r_7__31_,r_7__30_,r_7__29_,r_7__28_,r_7__27_,r_7__26_,r_7__25_,r_7__24_,
  r_7__23_,r_7__22_,r_7__21_,r_7__20_,r_7__19_,r_7__18_,r_7__17_,r_7__16_,r_7__15_,
  r_7__14_,r_7__13_,r_7__12_,r_7__11_,r_7__10_,r_7__9_,r_7__8_,r_7__7_,r_7__6_,
  r_7__5_,r_7__4_,r_7__3_,r_7__2_,r_7__1_,r_7__0_,r_8__63_,r_8__62_,r_8__61_,r_8__60_,
  r_8__59_,r_8__58_,r_8__57_,r_8__56_,r_8__55_,r_8__54_,r_8__53_,r_8__52_,r_8__51_,
  r_8__50_,r_8__49_,r_8__48_,r_8__47_,r_8__46_,r_8__45_,r_8__44_,r_8__43_,r_8__42_,
  r_8__41_,r_8__40_,r_8__39_,r_8__38_,r_8__37_,r_8__36_,r_8__35_,r_8__34_,
  r_8__33_,r_8__32_,r_8__31_,r_8__30_,r_8__29_,r_8__28_,r_8__27_,r_8__26_,r_8__25_,
  r_8__24_,r_8__23_,r_8__22_,r_8__21_,r_8__20_,r_8__19_,r_8__18_,r_8__17_,r_8__16_,
  r_8__15_,r_8__14_,r_8__13_,r_8__12_,r_8__11_,r_8__10_,r_8__9_,r_8__8_,r_8__7_,r_8__6_,
  r_8__5_,r_8__4_,r_8__3_,r_8__2_,r_8__1_,r_8__0_,r_9__63_,r_9__62_,r_9__61_,
  r_9__60_,r_9__59_,r_9__58_,r_9__57_,r_9__56_,r_9__55_,r_9__54_,r_9__53_,r_9__52_,
  r_9__51_,r_9__50_,r_9__49_,r_9__48_,r_9__47_,r_9__46_,r_9__45_,r_9__44_,r_9__43_,
  r_9__42_,r_9__41_,r_9__40_,r_9__39_,r_9__38_,r_9__37_,r_9__36_,r_9__35_,r_9__34_,
  r_9__33_,r_9__32_,r_9__31_,r_9__30_,r_9__29_,r_9__28_,r_9__27_,r_9__26_,r_9__25_,
  r_9__24_,r_9__23_,r_9__22_,r_9__21_,r_9__20_,r_9__19_,r_9__18_,r_9__17_,r_9__16_,
  r_9__15_,r_9__14_,r_9__13_,r_9__12_,r_9__11_,r_9__10_,r_9__9_,r_9__8_,r_9__7_,
  r_9__6_,r_9__5_,r_9__4_,r_9__3_,r_9__2_,r_9__1_,r_9__0_,r_10__63_,r_10__62_,
  r_10__61_,r_10__60_,r_10__59_,r_10__58_,r_10__57_,r_10__56_,r_10__55_,r_10__54_,
  r_10__53_,r_10__52_,r_10__51_,r_10__50_,r_10__49_,r_10__48_,r_10__47_,r_10__46_,
  r_10__45_,r_10__44_,r_10__43_,r_10__42_,r_10__41_,r_10__40_,r_10__39_,r_10__38_,
  r_10__37_,r_10__36_,r_10__35_,r_10__34_,r_10__33_,r_10__32_,r_10__31_,r_10__30_,
  r_10__29_,r_10__28_,r_10__27_,r_10__26_,r_10__25_,r_10__24_,r_10__23_,r_10__22_,
  r_10__21_,r_10__20_,r_10__19_,r_10__18_,r_10__17_,r_10__16_,r_10__15_,r_10__14_,
  r_10__13_,r_10__12_,r_10__11_,r_10__10_,r_10__9_,r_10__8_,r_10__7_,r_10__6_,r_10__5_,
  r_10__4_,r_10__3_,r_10__2_,r_10__1_,r_10__0_,r_11__63_,r_11__62_,r_11__61_,
  r_11__60_,r_11__59_,r_11__58_,r_11__57_,r_11__56_,r_11__55_,r_11__54_,r_11__53_,
  r_11__52_,r_11__51_,r_11__50_,r_11__49_,r_11__48_,r_11__47_,r_11__46_,r_11__45_,
  r_11__44_,r_11__43_,r_11__42_,r_11__41_,r_11__40_,r_11__39_,r_11__38_,r_11__37_,
  r_11__36_,r_11__35_,r_11__34_,r_11__33_,r_11__32_,r_11__31_,r_11__30_,r_11__29_,
  r_11__28_,r_11__27_,r_11__26_,r_11__25_,r_11__24_,r_11__23_,r_11__22_,r_11__21_,
  r_11__20_,r_11__19_,r_11__18_,r_11__17_,r_11__16_,r_11__15_,r_11__14_,r_11__13_,
  r_11__12_,r_11__11_,r_11__10_,r_11__9_,r_11__8_,r_11__7_,r_11__6_,r_11__5_,r_11__4_,
  r_11__3_,r_11__2_,r_11__1_,r_11__0_,r_12__63_,r_12__62_,r_12__61_,r_12__60_,
  r_12__59_,r_12__58_,r_12__57_,r_12__56_,r_12__55_,r_12__54_,r_12__53_,r_12__52_,
  r_12__51_,r_12__50_,r_12__49_,r_12__48_,r_12__47_,r_12__46_,r_12__45_,r_12__44_,
  r_12__43_,r_12__42_,r_12__41_,r_12__40_,r_12__39_,r_12__38_,r_12__37_,r_12__36_,
  r_12__35_,r_12__34_,r_12__33_,r_12__32_,r_12__31_,r_12__30_,r_12__29_,r_12__28_,
  r_12__27_,r_12__26_,r_12__25_,r_12__24_,r_12__23_,r_12__22_,r_12__21_,r_12__20_,
  r_12__19_,r_12__18_,r_12__17_,r_12__16_,r_12__15_,r_12__14_,r_12__13_,r_12__12_,
  r_12__11_,r_12__10_,r_12__9_,r_12__8_,r_12__7_,r_12__6_,r_12__5_,r_12__4_,r_12__3_,
  r_12__2_,r_12__1_,r_12__0_,r_13__63_,r_13__62_,r_13__61_,r_13__60_,r_13__59_,
  r_13__58_,r_13__57_,r_13__56_,r_13__55_,r_13__54_,r_13__53_,r_13__52_,r_13__51_,
  r_13__50_,r_13__49_,r_13__48_,r_13__47_,r_13__46_,r_13__45_,r_13__44_,r_13__43_,
  r_13__42_,r_13__41_,r_13__40_,r_13__39_,r_13__38_,r_13__37_,r_13__36_,r_13__35_,
  r_13__34_,r_13__33_,r_13__32_,r_13__31_,r_13__30_,r_13__29_,r_13__28_,r_13__27_,
  r_13__26_,r_13__25_,r_13__24_,r_13__23_,r_13__22_,r_13__21_,r_13__20_,r_13__19_,
  r_13__18_,r_13__17_,r_13__16_,r_13__15_,r_13__14_,r_13__13_,r_13__12_,r_13__11_,
  r_13__10_,r_13__9_,r_13__8_,r_13__7_,r_13__6_,r_13__5_,r_13__4_,r_13__3_,r_13__2_,
  r_13__1_,r_13__0_,r_14__63_,r_14__62_,r_14__61_,r_14__60_,r_14__59_,r_14__58_,
  r_14__57_,r_14__56_,r_14__55_,r_14__54_,r_14__53_,r_14__52_,r_14__51_,r_14__50_,
  r_14__49_,r_14__48_,r_14__47_,r_14__46_,r_14__45_,r_14__44_,r_14__43_,r_14__42_,
  r_14__41_,r_14__40_,r_14__39_,r_14__38_,r_14__37_,r_14__36_,r_14__35_,r_14__34_,
  r_14__33_,r_14__32_,r_14__31_,r_14__30_,r_14__29_,r_14__28_,r_14__27_,r_14__26_,
  r_14__25_,r_14__24_,r_14__23_,r_14__22_,r_14__21_,r_14__20_,r_14__19_,r_14__18_,
  r_14__17_,r_14__16_,r_14__15_,r_14__14_,r_14__13_,r_14__12_,r_14__11_,r_14__10_,
  r_14__9_,r_14__8_,r_14__7_,r_14__6_,r_14__5_,r_14__4_,r_14__3_,r_14__2_,r_14__1_,
  r_14__0_,r_15__63_,r_15__62_,r_15__61_,r_15__60_,r_15__59_,r_15__58_,r_15__57_,
  r_15__56_,r_15__55_,r_15__54_,r_15__53_,r_15__52_,r_15__51_,r_15__50_,r_15__49_,
  r_15__48_,r_15__47_,r_15__46_,r_15__45_,r_15__44_,r_15__43_,r_15__42_,r_15__41_,
  r_15__40_,r_15__39_,r_15__38_,r_15__37_,r_15__36_,r_15__35_,r_15__34_,r_15__33_,
  r_15__32_,r_15__31_,r_15__30_,r_15__29_,r_15__28_,r_15__27_,r_15__26_,r_15__25_,
  r_15__24_,r_15__23_,r_15__22_,r_15__21_,r_15__20_,r_15__19_,r_15__18_,r_15__17_,
  r_15__16_,r_15__15_,r_15__14_,r_15__13_,r_15__12_,r_15__11_,r_15__10_,r_15__9_,
  r_15__8_,r_15__7_,r_15__6_,r_15__5_,r_15__4_,r_15__3_,r_15__2_,r_15__1_,r_15__0_,
  r_16__63_,r_16__62_,r_16__61_,r_16__60_,r_16__59_,r_16__58_,r_16__57_,r_16__56_,
  r_16__55_,r_16__54_,r_16__53_,r_16__52_,r_16__51_,r_16__50_,r_16__49_,r_16__48_,
  r_16__47_,r_16__46_,r_16__45_,r_16__44_,r_16__43_,r_16__42_,r_16__41_,r_16__40_,
  r_16__39_,r_16__38_,r_16__37_,r_16__36_,r_16__35_,r_16__34_,r_16__33_,r_16__32_,
  r_16__31_,r_16__30_,r_16__29_,r_16__28_,r_16__27_,r_16__26_,r_16__25_,r_16__24_,
  r_16__23_,r_16__22_,r_16__21_,r_16__20_,r_16__19_,r_16__18_,r_16__17_,r_16__16_,
  r_16__15_,r_16__14_,r_16__13_,r_16__12_,r_16__11_,r_16__10_,r_16__9_,r_16__8_,
  r_16__7_,r_16__6_,r_16__5_,r_16__4_,r_16__3_,r_16__2_,r_16__1_,r_16__0_,r_17__63_,
  r_17__62_,r_17__61_,r_17__60_,r_17__59_,r_17__58_,r_17__57_,r_17__56_,r_17__55_,
  r_17__54_,r_17__53_,r_17__52_,r_17__51_,r_17__50_,r_17__49_,r_17__48_,r_17__47_,
  r_17__46_,r_17__45_,r_17__44_,r_17__43_,r_17__42_,r_17__41_,r_17__40_,r_17__39_,
  r_17__38_,r_17__37_,r_17__36_,r_17__35_,r_17__34_,r_17__33_,r_17__32_,r_17__31_,
  r_17__30_,r_17__29_,r_17__28_,r_17__27_,r_17__26_,r_17__25_,r_17__24_,r_17__23_,
  r_17__22_,r_17__21_,r_17__20_,r_17__19_,r_17__18_,r_17__17_,r_17__16_,r_17__15_,
  r_17__14_,r_17__13_,r_17__12_,r_17__11_,r_17__10_,r_17__9_,r_17__8_,r_17__7_,r_17__6_,
  r_17__5_,r_17__4_,r_17__3_,r_17__2_,r_17__1_,r_17__0_,r_18__63_,r_18__62_,
  r_18__61_,r_18__60_,r_18__59_,r_18__58_,r_18__57_,r_18__56_,r_18__55_,r_18__54_,
  r_18__53_,r_18__52_,r_18__51_,r_18__50_,r_18__49_,r_18__48_,r_18__47_,r_18__46_,
  r_18__45_,r_18__44_,r_18__43_,r_18__42_,r_18__41_,r_18__40_,r_18__39_,r_18__38_,
  r_18__37_,r_18__36_,r_18__35_,r_18__34_,r_18__33_,r_18__32_,r_18__31_,r_18__30_,
  r_18__29_,r_18__28_,r_18__27_,r_18__26_,r_18__25_,r_18__24_,r_18__23_,r_18__22_,
  r_18__21_,r_18__20_,r_18__19_,r_18__18_,r_18__17_,r_18__16_,r_18__15_,r_18__14_,
  r_18__13_,r_18__12_,r_18__11_,r_18__10_,r_18__9_,r_18__8_,r_18__7_,r_18__6_,r_18__5_,
  r_18__4_,r_18__3_,r_18__2_,r_18__1_,r_18__0_,r_19__63_,r_19__62_,r_19__61_,
  r_19__60_,r_19__59_,r_19__58_,r_19__57_,r_19__56_,r_19__55_,r_19__54_,r_19__53_,
  r_19__52_,r_19__51_,r_19__50_,r_19__49_,r_19__48_,r_19__47_,r_19__46_,r_19__45_,
  r_19__44_,r_19__43_,r_19__42_,r_19__41_,r_19__40_,r_19__39_,r_19__38_,r_19__37_,
  r_19__36_,r_19__35_,r_19__34_,r_19__33_,r_19__32_,r_19__31_,r_19__30_,r_19__29_,
  r_19__28_,r_19__27_,r_19__26_,r_19__25_,r_19__24_,r_19__23_,r_19__22_,r_19__21_,
  r_19__20_,r_19__19_,r_19__18_,r_19__17_,r_19__16_,r_19__15_,r_19__14_,r_19__13_,
  r_19__12_,r_19__11_,r_19__10_,r_19__9_,r_19__8_,r_19__7_,r_19__6_,r_19__5_,r_19__4_,
  r_19__3_,r_19__2_,r_19__1_,r_19__0_,r_20__63_,r_20__62_,r_20__61_,r_20__60_,
  r_20__59_,r_20__58_,r_20__57_,r_20__56_,r_20__55_,r_20__54_,r_20__53_,r_20__52_,
  r_20__51_,r_20__50_,r_20__49_,r_20__48_,r_20__47_,r_20__46_,r_20__45_,r_20__44_,
  r_20__43_,r_20__42_,r_20__41_,r_20__40_,r_20__39_,r_20__38_,r_20__37_,r_20__36_,
  r_20__35_,r_20__34_,r_20__33_,r_20__32_,r_20__31_,r_20__30_,r_20__29_,r_20__28_,
  r_20__27_,r_20__26_,r_20__25_,r_20__24_,r_20__23_,r_20__22_,r_20__21_,r_20__20_,
  r_20__19_,r_20__18_,r_20__17_,r_20__16_,r_20__15_,r_20__14_,r_20__13_,r_20__12_,
  r_20__11_,r_20__10_,r_20__9_,r_20__8_,r_20__7_,r_20__6_,r_20__5_,r_20__4_,r_20__3_,
  r_20__2_,r_20__1_,r_20__0_,r_21__63_,r_21__62_,r_21__61_,r_21__60_,r_21__59_,
  r_21__58_,r_21__57_,r_21__56_,r_21__55_,r_21__54_,r_21__53_,r_21__52_,r_21__51_,
  r_21__50_,r_21__49_,r_21__48_,r_21__47_,r_21__46_,r_21__45_,r_21__44_,r_21__43_,
  r_21__42_,r_21__41_,r_21__40_,r_21__39_,r_21__38_,r_21__37_,r_21__36_,r_21__35_,
  r_21__34_,r_21__33_,r_21__32_,r_21__31_,r_21__30_,r_21__29_,r_21__28_,r_21__27_,
  r_21__26_,r_21__25_,r_21__24_,r_21__23_,r_21__22_,r_21__21_,r_21__20_,r_21__19_,
  r_21__18_,r_21__17_,r_21__16_,r_21__15_,r_21__14_,r_21__13_,r_21__12_,r_21__11_,
  r_21__10_,r_21__9_,r_21__8_,r_21__7_,r_21__6_,r_21__5_,r_21__4_,r_21__3_,r_21__2_,
  r_21__1_,r_21__0_,r_22__63_,r_22__62_,r_22__61_,r_22__60_,r_22__59_,r_22__58_,
  r_22__57_,r_22__56_,r_22__55_,r_22__54_,r_22__53_,r_22__52_,r_22__51_,r_22__50_,
  r_22__49_,r_22__48_,r_22__47_,r_22__46_,r_22__45_,r_22__44_,r_22__43_,r_22__42_,
  r_22__41_,r_22__40_,r_22__39_,r_22__38_,r_22__37_,r_22__36_,r_22__35_,r_22__34_,
  r_22__33_,r_22__32_,r_22__31_,r_22__30_,r_22__29_,r_22__28_,r_22__27_,r_22__26_,
  r_22__25_,r_22__24_,r_22__23_,r_22__22_,r_22__21_,r_22__20_,r_22__19_,r_22__18_,
  r_22__17_,r_22__16_,r_22__15_,r_22__14_,r_22__13_,r_22__12_,r_22__11_,r_22__10_,
  r_22__9_,r_22__8_,r_22__7_,r_22__6_,r_22__5_,r_22__4_,r_22__3_,r_22__2_,r_22__1_,
  r_22__0_,r_23__63_,r_23__62_,r_23__61_,r_23__60_,r_23__59_,r_23__58_,r_23__57_,
  r_23__56_,r_23__55_,r_23__54_,r_23__53_,r_23__52_,r_23__51_,r_23__50_,r_23__49_,
  r_23__48_,r_23__47_,r_23__46_,r_23__45_,r_23__44_,r_23__43_,r_23__42_,r_23__41_,
  r_23__40_,r_23__39_,r_23__38_,r_23__37_,r_23__36_,r_23__35_,r_23__34_,r_23__33_,
  r_23__32_,r_23__31_,r_23__30_,r_23__29_,r_23__28_,r_23__27_,r_23__26_,r_23__25_,
  r_23__24_,r_23__23_,r_23__22_,r_23__21_,r_23__20_,r_23__19_,r_23__18_,r_23__17_,
  r_23__16_,r_23__15_,r_23__14_,r_23__13_,r_23__12_,r_23__11_,r_23__10_,r_23__9_,
  r_23__8_,r_23__7_,r_23__6_,r_23__5_,r_23__4_,r_23__3_,r_23__2_,r_23__1_,r_23__0_,
  r_24__63_,r_24__62_,r_24__61_,r_24__60_,r_24__59_,r_24__58_,r_24__57_,r_24__56_,
  r_24__55_,r_24__54_,r_24__53_,r_24__52_,r_24__51_,r_24__50_,r_24__49_,r_24__48_,
  r_24__47_,r_24__46_,r_24__45_,r_24__44_,r_24__43_,r_24__42_,r_24__41_,r_24__40_,
  r_24__39_,r_24__38_,r_24__37_,r_24__36_,r_24__35_,r_24__34_,r_24__33_,r_24__32_,
  r_24__31_,r_24__30_,r_24__29_,r_24__28_,r_24__27_,r_24__26_,r_24__25_,r_24__24_,
  r_24__23_,r_24__22_,r_24__21_,r_24__20_,r_24__19_,r_24__18_,r_24__17_,r_24__16_,
  r_24__15_,r_24__14_,r_24__13_,r_24__12_,r_24__11_,r_24__10_,r_24__9_,r_24__8_,
  r_24__7_,r_24__6_,r_24__5_,r_24__4_,r_24__3_,r_24__2_,r_24__1_,r_24__0_,r_25__63_,
  r_25__62_,r_25__61_,r_25__60_,r_25__59_,r_25__58_,r_25__57_,r_25__56_,r_25__55_,
  r_25__54_,r_25__53_,r_25__52_,r_25__51_,r_25__50_,r_25__49_,r_25__48_,r_25__47_,
  r_25__46_,r_25__45_,r_25__44_,r_25__43_,r_25__42_,r_25__41_,r_25__40_,r_25__39_,
  r_25__38_,r_25__37_,r_25__36_,r_25__35_,r_25__34_,r_25__33_,r_25__32_,r_25__31_,
  r_25__30_,r_25__29_,r_25__28_,r_25__27_,r_25__26_,r_25__25_,r_25__24_,r_25__23_,
  r_25__22_,r_25__21_,r_25__20_,r_25__19_,r_25__18_,r_25__17_,r_25__16_,r_25__15_,
  r_25__14_,r_25__13_,r_25__12_,r_25__11_,r_25__10_,r_25__9_,r_25__8_,r_25__7_,r_25__6_,
  r_25__5_,r_25__4_,r_25__3_,r_25__2_,r_25__1_,r_25__0_,r_26__63_,r_26__62_,
  r_26__61_,r_26__60_,r_26__59_,r_26__58_,r_26__57_,r_26__56_,r_26__55_,r_26__54_,
  r_26__53_,r_26__52_,r_26__51_,r_26__50_,r_26__49_,r_26__48_,r_26__47_,r_26__46_,
  r_26__45_,r_26__44_,r_26__43_,r_26__42_,r_26__41_,r_26__40_,r_26__39_,r_26__38_,
  r_26__37_,r_26__36_,r_26__35_,r_26__34_,r_26__33_,r_26__32_,r_26__31_,r_26__30_,
  r_26__29_,r_26__28_,r_26__27_,r_26__26_,r_26__25_,r_26__24_,r_26__23_,r_26__22_,
  r_26__21_,r_26__20_,r_26__19_,r_26__18_,r_26__17_,r_26__16_,r_26__15_,r_26__14_,
  r_26__13_,r_26__12_,r_26__11_,r_26__10_,r_26__9_,r_26__8_,r_26__7_,r_26__6_,r_26__5_,
  r_26__4_,r_26__3_,r_26__2_,r_26__1_,r_26__0_,r_27__63_,r_27__62_,r_27__61_,
  r_27__60_,r_27__59_,r_27__58_,r_27__57_,r_27__56_,r_27__55_,r_27__54_,r_27__53_,
  r_27__52_,r_27__51_,r_27__50_,r_27__49_,r_27__48_,r_27__47_,r_27__46_,r_27__45_,
  r_27__44_,r_27__43_,r_27__42_,r_27__41_,r_27__40_,r_27__39_,r_27__38_,r_27__37_,
  r_27__36_,r_27__35_,r_27__34_,r_27__33_,r_27__32_,r_27__31_,r_27__30_,r_27__29_,
  r_27__28_,r_27__27_,r_27__26_,r_27__25_,r_27__24_,r_27__23_,r_27__22_,r_27__21_,
  r_27__20_,r_27__19_,r_27__18_,r_27__17_,r_27__16_,r_27__15_,r_27__14_,r_27__13_,
  r_27__12_,r_27__11_,r_27__10_,r_27__9_,r_27__8_,r_27__7_,r_27__6_,r_27__5_,r_27__4_,
  r_27__3_,r_27__2_,r_27__1_,r_27__0_,r_28__63_,r_28__62_,r_28__61_,r_28__60_,
  r_28__59_,r_28__58_,r_28__57_,r_28__56_,r_28__55_,r_28__54_,r_28__53_,r_28__52_,
  r_28__51_,r_28__50_,r_28__49_,r_28__48_,r_28__47_,r_28__46_,r_28__45_,r_28__44_,
  r_28__43_,r_28__42_,r_28__41_,r_28__40_,r_28__39_,r_28__38_,r_28__37_,r_28__36_,
  r_28__35_,r_28__34_,r_28__33_,r_28__32_,r_28__31_,r_28__30_,r_28__29_,r_28__28_,
  r_28__27_,r_28__26_,r_28__25_,r_28__24_,r_28__23_,r_28__22_,r_28__21_,r_28__20_,
  r_28__19_,r_28__18_,r_28__17_,r_28__16_,r_28__15_,r_28__14_,r_28__13_,r_28__12_,
  r_28__11_,r_28__10_,r_28__9_,r_28__8_,r_28__7_,r_28__6_,r_28__5_,r_28__4_,r_28__3_,
  r_28__2_,r_28__1_,r_28__0_,r_29__63_,r_29__62_,r_29__61_,r_29__60_,r_29__59_,
  r_29__58_,r_29__57_,r_29__56_,r_29__55_,r_29__54_,r_29__53_,r_29__52_,r_29__51_,
  r_29__50_,r_29__49_,r_29__48_,r_29__47_,r_29__46_,r_29__45_,r_29__44_,r_29__43_,
  r_29__42_,r_29__41_,r_29__40_,r_29__39_,r_29__38_,r_29__37_,r_29__36_,r_29__35_,
  r_29__34_,r_29__33_,r_29__32_,r_29__31_,r_29__30_,r_29__29_,r_29__28_,r_29__27_,
  r_29__26_,r_29__25_,r_29__24_,r_29__23_,r_29__22_,r_29__21_,r_29__20_,r_29__19_,
  r_29__18_,r_29__17_,r_29__16_,r_29__15_,r_29__14_,r_29__13_,r_29__12_,r_29__11_,
  r_29__10_,r_29__9_,r_29__8_,r_29__7_,r_29__6_,r_29__5_,r_29__4_,r_29__3_,r_29__2_,
  r_29__1_,r_29__0_,r_30__63_,r_30__62_,r_30__61_,r_30__60_,r_30__59_,r_30__58_,
  r_30__57_,r_30__56_,r_30__55_,r_30__54_,r_30__53_,r_30__52_,r_30__51_,r_30__50_,
  r_30__49_,r_30__48_,r_30__47_,r_30__46_,r_30__45_,r_30__44_,r_30__43_,r_30__42_,
  r_30__41_,r_30__40_,r_30__39_,r_30__38_,r_30__37_,r_30__36_,r_30__35_,r_30__34_,
  r_30__33_,r_30__32_,r_30__31_,r_30__30_,r_30__29_,r_30__28_,r_30__27_,r_30__26_,
  r_30__25_,r_30__24_,r_30__23_,r_30__22_,r_30__21_,r_30__20_,r_30__19_,r_30__18_,
  r_30__17_,r_30__16_,r_30__15_,r_30__14_,r_30__13_,r_30__12_,r_30__11_,r_30__10_,
  r_30__9_,r_30__8_,r_30__7_,r_30__6_,r_30__5_,r_30__4_,r_30__3_,r_30__2_,r_30__1_,
  r_30__0_,r_31__63_,r_31__62_,r_31__61_,r_31__60_,r_31__59_,r_31__58_,r_31__57_,
  r_31__56_,r_31__55_,r_31__54_,r_31__53_,r_31__52_,r_31__51_,r_31__50_,r_31__49_,
  r_31__48_,r_31__47_,r_31__46_,r_31__45_,r_31__44_,r_31__43_,r_31__42_,r_31__41_,
  r_31__40_,r_31__39_,r_31__38_,r_31__37_,r_31__36_,r_31__35_,r_31__34_,r_31__33_,
  r_31__32_,r_31__31_,r_31__30_,r_31__29_,r_31__28_,r_31__27_,r_31__26_,r_31__25_,
  r_31__24_,r_31__23_,r_31__22_,r_31__21_,r_31__20_,r_31__19_,r_31__18_,r_31__17_,
  r_31__16_,r_31__15_,r_31__14_,r_31__13_,r_31__12_,r_31__11_,r_31__10_,r_31__9_,
  r_31__8_,r_31__7_,r_31__6_,r_31__5_,r_31__4_,r_31__3_,r_31__2_,r_31__1_,r_31__0_,
  r_32__63_,r_32__62_,r_32__61_,r_32__60_,r_32__59_,r_32__58_,r_32__57_,r_32__56_,
  r_32__55_,r_32__54_,r_32__53_,r_32__52_,r_32__51_,r_32__50_,r_32__49_,r_32__48_,
  r_32__47_,r_32__46_,r_32__45_,r_32__44_,r_32__43_,r_32__42_,r_32__41_,r_32__40_,
  r_32__39_,r_32__38_,r_32__37_,r_32__36_,r_32__35_,r_32__34_,r_32__33_,r_32__32_,
  r_32__31_,r_32__30_,r_32__29_,r_32__28_,r_32__27_,r_32__26_,r_32__25_,r_32__24_,
  r_32__23_,r_32__22_,r_32__21_,r_32__20_,r_32__19_,r_32__18_,r_32__17_,r_32__16_,
  r_32__15_,r_32__14_,r_32__13_,r_32__12_,r_32__11_,r_32__10_,r_32__9_,r_32__8_,
  r_32__7_,r_32__6_,r_32__5_,r_32__4_,r_32__3_,r_32__2_,r_32__1_,r_32__0_,r_33__63_,
  r_33__62_,r_33__61_,r_33__60_,r_33__59_,r_33__58_,r_33__57_,r_33__56_,r_33__55_,
  r_33__54_,r_33__53_,r_33__52_,r_33__51_,r_33__50_,r_33__49_,r_33__48_,r_33__47_,
  r_33__46_,r_33__45_,r_33__44_,r_33__43_,r_33__42_,r_33__41_,r_33__40_,r_33__39_,
  r_33__38_,r_33__37_,r_33__36_,r_33__35_,r_33__34_,r_33__33_,r_33__32_,r_33__31_,
  r_33__30_,r_33__29_,r_33__28_,r_33__27_,r_33__26_,r_33__25_,r_33__24_,r_33__23_,
  r_33__22_,r_33__21_,r_33__20_,r_33__19_,r_33__18_,r_33__17_,r_33__16_,r_33__15_,
  r_33__14_,r_33__13_,r_33__12_,r_33__11_,r_33__10_,r_33__9_,r_33__8_,r_33__7_,r_33__6_,
  r_33__5_,r_33__4_,r_33__3_,r_33__2_,r_33__1_,r_33__0_,r_34__63_,r_34__62_,
  r_34__61_,r_34__60_,r_34__59_,r_34__58_,r_34__57_,r_34__56_,r_34__55_,r_34__54_,
  r_34__53_,r_34__52_,r_34__51_,r_34__50_,r_34__49_,r_34__48_,r_34__47_,r_34__46_,
  r_34__45_,r_34__44_,r_34__43_,r_34__42_,r_34__41_,r_34__40_,r_34__39_,r_34__38_,
  r_34__37_,r_34__36_,r_34__35_,r_34__34_,r_34__33_,r_34__32_,r_34__31_,r_34__30_,
  r_34__29_,r_34__28_,r_34__27_,r_34__26_,r_34__25_,r_34__24_,r_34__23_,r_34__22_,
  r_34__21_,r_34__20_,r_34__19_,r_34__18_,r_34__17_,r_34__16_,r_34__15_,r_34__14_,
  r_34__13_,r_34__12_,r_34__11_,r_34__10_,r_34__9_,r_34__8_,r_34__7_,r_34__6_,r_34__5_,
  r_34__4_,r_34__3_,r_34__2_,r_34__1_,r_34__0_,r_35__63_,r_35__62_,r_35__61_,
  r_35__60_,r_35__59_,r_35__58_,r_35__57_,r_35__56_,r_35__55_,r_35__54_,r_35__53_,
  r_35__52_,r_35__51_,r_35__50_,r_35__49_,r_35__48_,r_35__47_,r_35__46_,r_35__45_,
  r_35__44_,r_35__43_,r_35__42_,r_35__41_,r_35__40_,r_35__39_,r_35__38_,r_35__37_,
  r_35__36_,r_35__35_,r_35__34_,r_35__33_,r_35__32_,r_35__31_,r_35__30_,r_35__29_,
  r_35__28_,r_35__27_,r_35__26_,r_35__25_,r_35__24_,r_35__23_,r_35__22_,r_35__21_,
  r_35__20_,r_35__19_,r_35__18_,r_35__17_,r_35__16_,r_35__15_,r_35__14_,r_35__13_,
  r_35__12_,r_35__11_,r_35__10_,r_35__9_,r_35__8_,r_35__7_,r_35__6_,r_35__5_,r_35__4_,
  r_35__3_,r_35__2_,r_35__1_,r_35__0_,r_36__63_,r_36__62_,r_36__61_,r_36__60_,
  r_36__59_,r_36__58_,r_36__57_,r_36__56_,r_36__55_,r_36__54_,r_36__53_,r_36__52_,
  r_36__51_,r_36__50_,r_36__49_,r_36__48_,r_36__47_,r_36__46_,r_36__45_,r_36__44_,
  r_36__43_,r_36__42_,r_36__41_,r_36__40_,r_36__39_,r_36__38_,r_36__37_,r_36__36_,
  r_36__35_,r_36__34_,r_36__33_,r_36__32_,r_36__31_,r_36__30_,r_36__29_,r_36__28_,
  r_36__27_,r_36__26_,r_36__25_,r_36__24_,r_36__23_,r_36__22_,r_36__21_,r_36__20_,
  r_36__19_,r_36__18_,r_36__17_,r_36__16_,r_36__15_,r_36__14_,r_36__13_,r_36__12_,
  r_36__11_,r_36__10_,r_36__9_,r_36__8_,r_36__7_,r_36__6_,r_36__5_,r_36__4_,r_36__3_,
  r_36__2_,r_36__1_,r_36__0_,r_37__63_,r_37__62_,r_37__61_,r_37__60_,r_37__59_,
  r_37__58_,r_37__57_,r_37__56_,r_37__55_,r_37__54_,r_37__53_,r_37__52_,r_37__51_,
  r_37__50_,r_37__49_,r_37__48_,r_37__47_,r_37__46_,r_37__45_,r_37__44_,r_37__43_,
  r_37__42_,r_37__41_,r_37__40_,r_37__39_,r_37__38_,r_37__37_,r_37__36_,r_37__35_,
  r_37__34_,r_37__33_,r_37__32_,r_37__31_,r_37__30_,r_37__29_,r_37__28_,r_37__27_,
  r_37__26_,r_37__25_,r_37__24_,r_37__23_,r_37__22_,r_37__21_,r_37__20_,r_37__19_,
  r_37__18_,r_37__17_,r_37__16_,r_37__15_,r_37__14_,r_37__13_,r_37__12_,r_37__11_,
  r_37__10_,r_37__9_,r_37__8_,r_37__7_,r_37__6_,r_37__5_,r_37__4_,r_37__3_,r_37__2_,
  r_37__1_,r_37__0_,r_38__63_,r_38__62_,r_38__61_,r_38__60_,r_38__59_,r_38__58_,
  r_38__57_,r_38__56_,r_38__55_,r_38__54_,r_38__53_,r_38__52_,r_38__51_,r_38__50_,
  r_38__49_,r_38__48_,r_38__47_,r_38__46_,r_38__45_,r_38__44_,r_38__43_,r_38__42_,
  r_38__41_,r_38__40_,r_38__39_,r_38__38_,r_38__37_,r_38__36_,r_38__35_,r_38__34_,
  r_38__33_,r_38__32_,r_38__31_,r_38__30_,r_38__29_,r_38__28_,r_38__27_,r_38__26_,
  r_38__25_,r_38__24_,r_38__23_,r_38__22_,r_38__21_,r_38__20_,r_38__19_,r_38__18_,
  r_38__17_,r_38__16_,r_38__15_,r_38__14_,r_38__13_,r_38__12_,r_38__11_,r_38__10_,
  r_38__9_,r_38__8_,r_38__7_,r_38__6_,r_38__5_,r_38__4_,r_38__3_,r_38__2_,r_38__1_,
  r_38__0_,r_39__63_,r_39__62_,r_39__61_,r_39__60_,r_39__59_,r_39__58_,r_39__57_,
  r_39__56_,r_39__55_,r_39__54_,r_39__53_,r_39__52_,r_39__51_,r_39__50_,r_39__49_,
  r_39__48_,r_39__47_,r_39__46_,r_39__45_,r_39__44_,r_39__43_,r_39__42_,r_39__41_,
  r_39__40_,r_39__39_,r_39__38_,r_39__37_,r_39__36_,r_39__35_,r_39__34_,r_39__33_,
  r_39__32_,r_39__31_,r_39__30_,r_39__29_,r_39__28_,r_39__27_,r_39__26_,r_39__25_,
  r_39__24_,r_39__23_,r_39__22_,r_39__21_,r_39__20_,r_39__19_,r_39__18_,r_39__17_,
  r_39__16_,r_39__15_,r_39__14_,r_39__13_,r_39__12_,r_39__11_,r_39__10_,r_39__9_,
  r_39__8_,r_39__7_,r_39__6_,r_39__5_,r_39__4_,r_39__3_,r_39__2_,r_39__1_,r_39__0_,
  r_40__63_,r_40__62_,r_40__61_,r_40__60_,r_40__59_,r_40__58_,r_40__57_,r_40__56_,
  r_40__55_,r_40__54_,r_40__53_,r_40__52_,r_40__51_,r_40__50_,r_40__49_,r_40__48_,
  r_40__47_,r_40__46_,r_40__45_,r_40__44_,r_40__43_,r_40__42_,r_40__41_,r_40__40_,
  r_40__39_,r_40__38_,r_40__37_,r_40__36_,r_40__35_,r_40__34_,r_40__33_,r_40__32_,
  r_40__31_,r_40__30_,r_40__29_,r_40__28_,r_40__27_,r_40__26_,r_40__25_,r_40__24_,
  r_40__23_,r_40__22_,r_40__21_,r_40__20_,r_40__19_,r_40__18_,r_40__17_,r_40__16_,
  r_40__15_,r_40__14_,r_40__13_,r_40__12_,r_40__11_,r_40__10_,r_40__9_,r_40__8_,
  r_40__7_,r_40__6_,r_40__5_,r_40__4_,r_40__3_,r_40__2_,r_40__1_,r_40__0_,r_41__63_,
  r_41__62_,r_41__61_,r_41__60_,r_41__59_,r_41__58_,r_41__57_,r_41__56_,r_41__55_,
  r_41__54_,r_41__53_,r_41__52_,r_41__51_,r_41__50_,r_41__49_,r_41__48_,r_41__47_,
  r_41__46_,r_41__45_,r_41__44_,r_41__43_,r_41__42_,r_41__41_,r_41__40_,r_41__39_,
  r_41__38_,r_41__37_,r_41__36_,r_41__35_,r_41__34_,r_41__33_,r_41__32_,r_41__31_,
  r_41__30_,r_41__29_,r_41__28_,r_41__27_,r_41__26_,r_41__25_,r_41__24_,r_41__23_,
  r_41__22_,r_41__21_,r_41__20_,r_41__19_,r_41__18_,r_41__17_,r_41__16_,r_41__15_,
  r_41__14_,r_41__13_,r_41__12_,r_41__11_,r_41__10_,r_41__9_,r_41__8_,r_41__7_,r_41__6_,
  r_41__5_,r_41__4_,r_41__3_,r_41__2_,r_41__1_,r_41__0_,r_42__63_,r_42__62_,
  r_42__61_,r_42__60_,r_42__59_,r_42__58_,r_42__57_,r_42__56_,r_42__55_,r_42__54_,
  r_42__53_,r_42__52_,r_42__51_,r_42__50_,r_42__49_,r_42__48_,r_42__47_,r_42__46_,
  r_42__45_,r_42__44_,r_42__43_,r_42__42_,r_42__41_,r_42__40_,r_42__39_,r_42__38_,
  r_42__37_,r_42__36_,r_42__35_,r_42__34_,r_42__33_,r_42__32_,r_42__31_,r_42__30_,
  r_42__29_,r_42__28_,r_42__27_,r_42__26_,r_42__25_,r_42__24_,r_42__23_,r_42__22_,
  r_42__21_,r_42__20_,r_42__19_,r_42__18_,r_42__17_,r_42__16_,r_42__15_,r_42__14_,
  r_42__13_,r_42__12_,r_42__11_,r_42__10_,r_42__9_,r_42__8_,r_42__7_,r_42__6_,r_42__5_,
  r_42__4_,r_42__3_,r_42__2_,r_42__1_,r_42__0_,r_43__63_,r_43__62_,r_43__61_,
  r_43__60_,r_43__59_,r_43__58_,r_43__57_,r_43__56_,r_43__55_,r_43__54_,r_43__53_,
  r_43__52_,r_43__51_,r_43__50_,r_43__49_,r_43__48_,r_43__47_,r_43__46_,r_43__45_,
  r_43__44_,r_43__43_,r_43__42_,r_43__41_,r_43__40_,r_43__39_,r_43__38_,r_43__37_,
  r_43__36_,r_43__35_,r_43__34_,r_43__33_,r_43__32_,r_43__31_,r_43__30_,r_43__29_,
  r_43__28_,r_43__27_,r_43__26_,r_43__25_,r_43__24_,r_43__23_,r_43__22_,r_43__21_,
  r_43__20_,r_43__19_,r_43__18_,r_43__17_,r_43__16_,r_43__15_,r_43__14_,r_43__13_,
  r_43__12_,r_43__11_,r_43__10_,r_43__9_,r_43__8_,r_43__7_,r_43__6_,r_43__5_,r_43__4_,
  r_43__3_,r_43__2_,r_43__1_,r_43__0_,r_44__63_,r_44__62_,r_44__61_,r_44__60_,
  r_44__59_,r_44__58_,r_44__57_,r_44__56_,r_44__55_,r_44__54_,r_44__53_,r_44__52_,
  r_44__51_,r_44__50_,r_44__49_,r_44__48_,r_44__47_,r_44__46_,r_44__45_,r_44__44_,
  r_44__43_,r_44__42_,r_44__41_,r_44__40_,r_44__39_,r_44__38_,r_44__37_,r_44__36_,
  r_44__35_,r_44__34_,r_44__33_,r_44__32_,r_44__31_,r_44__30_,r_44__29_,r_44__28_,
  r_44__27_,r_44__26_,r_44__25_,r_44__24_,r_44__23_,r_44__22_,r_44__21_,r_44__20_,
  r_44__19_,r_44__18_,r_44__17_,r_44__16_,r_44__15_,r_44__14_,r_44__13_,r_44__12_,
  r_44__11_,r_44__10_,r_44__9_,r_44__8_,r_44__7_,r_44__6_,r_44__5_,r_44__4_,r_44__3_,
  r_44__2_,r_44__1_,r_44__0_,r_45__63_,r_45__62_,r_45__61_,r_45__60_,r_45__59_,
  r_45__58_,r_45__57_,r_45__56_,r_45__55_,r_45__54_,r_45__53_,r_45__52_,r_45__51_,
  r_45__50_,r_45__49_,r_45__48_,r_45__47_,r_45__46_,r_45__45_,r_45__44_,r_45__43_,
  r_45__42_,r_45__41_,r_45__40_,r_45__39_,r_45__38_,r_45__37_,r_45__36_,r_45__35_,
  r_45__34_,r_45__33_,r_45__32_,r_45__31_,r_45__30_,r_45__29_,r_45__28_,r_45__27_,
  r_45__26_,r_45__25_,r_45__24_,r_45__23_,r_45__22_,r_45__21_,r_45__20_,r_45__19_,
  r_45__18_,r_45__17_,r_45__16_,r_45__15_,r_45__14_,r_45__13_,r_45__12_,r_45__11_,
  r_45__10_,r_45__9_,r_45__8_,r_45__7_,r_45__6_,r_45__5_,r_45__4_,r_45__3_,r_45__2_,
  r_45__1_,r_45__0_,r_46__63_,r_46__62_,r_46__61_,r_46__60_,r_46__59_,r_46__58_,
  r_46__57_,r_46__56_,r_46__55_,r_46__54_,r_46__53_,r_46__52_,r_46__51_,r_46__50_,
  r_46__49_,r_46__48_,r_46__47_,r_46__46_,r_46__45_,r_46__44_,r_46__43_,r_46__42_,
  r_46__41_,r_46__40_,r_46__39_,r_46__38_,r_46__37_,r_46__36_,r_46__35_,r_46__34_,
  r_46__33_,r_46__32_,r_46__31_,r_46__30_,r_46__29_,r_46__28_,r_46__27_,r_46__26_,
  r_46__25_,r_46__24_,r_46__23_,r_46__22_,r_46__21_,r_46__20_,r_46__19_,r_46__18_,
  r_46__17_,r_46__16_,r_46__15_,r_46__14_,r_46__13_,r_46__12_,r_46__11_,r_46__10_,
  r_46__9_,r_46__8_,r_46__7_,r_46__6_,r_46__5_,r_46__4_,r_46__3_,r_46__2_,r_46__1_,
  r_46__0_,r_47__63_,r_47__62_,r_47__61_,r_47__60_,r_47__59_,r_47__58_,r_47__57_,
  r_47__56_,r_47__55_,r_47__54_,r_47__53_,r_47__52_,r_47__51_,r_47__50_,r_47__49_,
  r_47__48_,r_47__47_,r_47__46_,r_47__45_,r_47__44_,r_47__43_,r_47__42_,r_47__41_,
  r_47__40_,r_47__39_,r_47__38_,r_47__37_,r_47__36_,r_47__35_,r_47__34_,r_47__33_,
  r_47__32_,r_47__31_,r_47__30_,r_47__29_,r_47__28_,r_47__27_,r_47__26_,r_47__25_,
  r_47__24_,r_47__23_,r_47__22_,r_47__21_,r_47__20_,r_47__19_,r_47__18_,r_47__17_,
  r_47__16_,r_47__15_,r_47__14_,r_47__13_,r_47__12_,r_47__11_,r_47__10_,r_47__9_,
  r_47__8_,r_47__7_,r_47__6_,r_47__5_,r_47__4_,r_47__3_,r_47__2_,r_47__1_,r_47__0_,
  r_48__63_,r_48__62_,r_48__61_,r_48__60_,r_48__59_,r_48__58_,r_48__57_,r_48__56_,
  r_48__55_,r_48__54_,r_48__53_,r_48__52_,r_48__51_,r_48__50_,r_48__49_,r_48__48_,
  r_48__47_,r_48__46_,r_48__45_,r_48__44_,r_48__43_,r_48__42_,r_48__41_,r_48__40_,
  r_48__39_,r_48__38_,r_48__37_,r_48__36_,r_48__35_,r_48__34_,r_48__33_,r_48__32_,
  r_48__31_,r_48__30_,r_48__29_,r_48__28_,r_48__27_,r_48__26_,r_48__25_,r_48__24_,
  r_48__23_,r_48__22_,r_48__21_,r_48__20_,r_48__19_,r_48__18_,r_48__17_,r_48__16_,
  r_48__15_,r_48__14_,r_48__13_,r_48__12_,r_48__11_,r_48__10_,r_48__9_,r_48__8_,
  r_48__7_,r_48__6_,r_48__5_,r_48__4_,r_48__3_,r_48__2_,r_48__1_,r_48__0_,r_49__63_,
  r_49__62_,r_49__61_,r_49__60_,r_49__59_,r_49__58_,r_49__57_,r_49__56_,r_49__55_,
  r_49__54_,r_49__53_,r_49__52_,r_49__51_,r_49__50_,r_49__49_,r_49__48_,r_49__47_,
  r_49__46_,r_49__45_,r_49__44_,r_49__43_,r_49__42_,r_49__41_,r_49__40_,r_49__39_,
  r_49__38_,r_49__37_,r_49__36_,r_49__35_,r_49__34_,r_49__33_,r_49__32_,r_49__31_,
  r_49__30_,r_49__29_,r_49__28_,r_49__27_,r_49__26_,r_49__25_,r_49__24_,r_49__23_,
  r_49__22_,r_49__21_,r_49__20_,r_49__19_,r_49__18_,r_49__17_,r_49__16_,r_49__15_,
  r_49__14_,r_49__13_,r_49__12_,r_49__11_,r_49__10_,r_49__9_,r_49__8_,r_49__7_,r_49__6_,
  r_49__5_,r_49__4_,r_49__3_,r_49__2_,r_49__1_,r_49__0_,r_50__63_,r_50__62_,
  r_50__61_,r_50__60_,r_50__59_,r_50__58_,r_50__57_,r_50__56_,r_50__55_,r_50__54_,
  r_50__53_,r_50__52_,r_50__51_,r_50__50_,r_50__49_,r_50__48_,r_50__47_,r_50__46_,
  r_50__45_,r_50__44_,r_50__43_,r_50__42_,r_50__41_,r_50__40_,r_50__39_,r_50__38_,
  r_50__37_,r_50__36_,r_50__35_,r_50__34_,r_50__33_,r_50__32_,r_50__31_,r_50__30_,
  r_50__29_,r_50__28_,r_50__27_,r_50__26_,r_50__25_,r_50__24_,r_50__23_,r_50__22_,
  r_50__21_,r_50__20_,r_50__19_,r_50__18_,r_50__17_,r_50__16_,r_50__15_,r_50__14_,
  r_50__13_,r_50__12_,r_50__11_,r_50__10_,r_50__9_,r_50__8_,r_50__7_,r_50__6_,r_50__5_,
  r_50__4_,r_50__3_,r_50__2_,r_50__1_,r_50__0_,r_51__63_,r_51__62_,r_51__61_,
  r_51__60_,r_51__59_,r_51__58_,r_51__57_,r_51__56_,r_51__55_,r_51__54_,r_51__53_,
  r_51__52_,r_51__51_,r_51__50_,r_51__49_,r_51__48_,r_51__47_,r_51__46_,r_51__45_,
  r_51__44_,r_51__43_,r_51__42_,r_51__41_,r_51__40_,r_51__39_,r_51__38_,r_51__37_,
  r_51__36_,r_51__35_,r_51__34_,r_51__33_,r_51__32_,r_51__31_,r_51__30_,r_51__29_,
  r_51__28_,r_51__27_,r_51__26_,r_51__25_,r_51__24_,r_51__23_,r_51__22_,r_51__21_,
  r_51__20_,r_51__19_,r_51__18_,r_51__17_,r_51__16_,r_51__15_,r_51__14_,r_51__13_,
  r_51__12_,r_51__11_,r_51__10_,r_51__9_,r_51__8_,r_51__7_,r_51__6_,r_51__5_,r_51__4_,
  r_51__3_,r_51__2_,r_51__1_,r_51__0_,r_52__63_,r_52__62_,r_52__61_,r_52__60_,
  r_52__59_,r_52__58_,r_52__57_,r_52__56_,r_52__55_,r_52__54_,r_52__53_,r_52__52_,
  r_52__51_,r_52__50_,r_52__49_,r_52__48_,r_52__47_,r_52__46_,r_52__45_,r_52__44_,
  r_52__43_,r_52__42_,r_52__41_,r_52__40_,r_52__39_,r_52__38_,r_52__37_,r_52__36_,
  r_52__35_,r_52__34_,r_52__33_,r_52__32_,r_52__31_,r_52__30_,r_52__29_,r_52__28_,
  r_52__27_,r_52__26_,r_52__25_,r_52__24_,r_52__23_,r_52__22_,r_52__21_,r_52__20_,
  r_52__19_,r_52__18_,r_52__17_,r_52__16_,r_52__15_,r_52__14_,r_52__13_,r_52__12_,
  r_52__11_,r_52__10_,r_52__9_,r_52__8_,r_52__7_,r_52__6_,r_52__5_,r_52__4_,r_52__3_,
  r_52__2_,r_52__1_,r_52__0_,r_53__63_,r_53__62_,r_53__61_,r_53__60_,r_53__59_,
  r_53__58_,r_53__57_,r_53__56_,r_53__55_,r_53__54_,r_53__53_,r_53__52_,r_53__51_,
  r_53__50_,r_53__49_,r_53__48_,r_53__47_,r_53__46_,r_53__45_,r_53__44_,r_53__43_,
  r_53__42_,r_53__41_,r_53__40_,r_53__39_,r_53__38_,r_53__37_,r_53__36_,r_53__35_,
  r_53__34_,r_53__33_,r_53__32_,r_53__31_,r_53__30_,r_53__29_,r_53__28_,r_53__27_,
  r_53__26_,r_53__25_,r_53__24_,r_53__23_,r_53__22_,r_53__21_,r_53__20_,r_53__19_,
  r_53__18_,r_53__17_,r_53__16_,r_53__15_,r_53__14_,r_53__13_,r_53__12_,r_53__11_,
  r_53__10_,r_53__9_,r_53__8_,r_53__7_,r_53__6_,r_53__5_,r_53__4_,r_53__3_,r_53__2_,
  r_53__1_,r_53__0_,r_54__63_,r_54__62_,r_54__61_,r_54__60_,r_54__59_,r_54__58_,
  r_54__57_,r_54__56_,r_54__55_,r_54__54_,r_54__53_,r_54__52_,r_54__51_,r_54__50_,
  r_54__49_,r_54__48_,r_54__47_,r_54__46_,r_54__45_,r_54__44_,r_54__43_,r_54__42_,
  r_54__41_,r_54__40_,r_54__39_,r_54__38_,r_54__37_,r_54__36_,r_54__35_,r_54__34_,
  r_54__33_,r_54__32_,r_54__31_,r_54__30_,r_54__29_,r_54__28_,r_54__27_,r_54__26_,
  r_54__25_,r_54__24_,r_54__23_,r_54__22_,r_54__21_,r_54__20_,r_54__19_,r_54__18_,
  r_54__17_,r_54__16_,r_54__15_,r_54__14_,r_54__13_,r_54__12_,r_54__11_,r_54__10_,
  r_54__9_,r_54__8_,r_54__7_,r_54__6_,r_54__5_,r_54__4_,r_54__3_,r_54__2_,r_54__1_,
  r_54__0_,r_55__63_,r_55__62_,r_55__61_,r_55__60_,r_55__59_,r_55__58_,r_55__57_,
  r_55__56_,r_55__55_,r_55__54_,r_55__53_,r_55__52_,r_55__51_,r_55__50_,r_55__49_,
  r_55__48_,r_55__47_,r_55__46_,r_55__45_,r_55__44_,r_55__43_,r_55__42_,r_55__41_,
  r_55__40_,r_55__39_,r_55__38_,r_55__37_,r_55__36_,r_55__35_,r_55__34_,r_55__33_,
  r_55__32_,r_55__31_,r_55__30_,r_55__29_,r_55__28_,r_55__27_,r_55__26_,r_55__25_,
  r_55__24_,r_55__23_,r_55__22_,r_55__21_,r_55__20_,r_55__19_,r_55__18_,r_55__17_,
  r_55__16_,r_55__15_,r_55__14_,r_55__13_,r_55__12_,r_55__11_,r_55__10_,r_55__9_,
  r_55__8_,r_55__7_,r_55__6_,r_55__5_,r_55__4_,r_55__3_,r_55__2_,r_55__1_,r_55__0_,
  r_56__63_,r_56__62_,r_56__61_,r_56__60_,r_56__59_,r_56__58_,r_56__57_,r_56__56_,
  r_56__55_,r_56__54_,r_56__53_,r_56__52_,r_56__51_,r_56__50_,r_56__49_,r_56__48_,
  r_56__47_,r_56__46_,r_56__45_,r_56__44_,r_56__43_,r_56__42_,r_56__41_,r_56__40_,
  r_56__39_,r_56__38_,r_56__37_,r_56__36_,r_56__35_,r_56__34_,r_56__33_,r_56__32_,
  r_56__31_,r_56__30_,r_56__29_,r_56__28_,r_56__27_,r_56__26_,r_56__25_,r_56__24_,
  r_56__23_,r_56__22_,r_56__21_,r_56__20_,r_56__19_,r_56__18_,r_56__17_,r_56__16_,
  r_56__15_,r_56__14_,r_56__13_,r_56__12_,r_56__11_,r_56__10_,r_56__9_,r_56__8_,
  r_56__7_,r_56__6_,r_56__5_,r_56__4_,r_56__3_,r_56__2_,r_56__1_,r_56__0_,r_57__63_,
  r_57__62_,r_57__61_,r_57__60_,r_57__59_,r_57__58_,r_57__57_,r_57__56_,r_57__55_,
  r_57__54_,r_57__53_,r_57__52_,r_57__51_,r_57__50_,r_57__49_,r_57__48_,r_57__47_,
  r_57__46_,r_57__45_,r_57__44_,r_57__43_,r_57__42_,r_57__41_,r_57__40_,r_57__39_,
  r_57__38_,r_57__37_,r_57__36_,r_57__35_,r_57__34_,r_57__33_,r_57__32_,r_57__31_,
  r_57__30_,r_57__29_,r_57__28_,r_57__27_,r_57__26_,r_57__25_,r_57__24_,r_57__23_,
  r_57__22_,r_57__21_,r_57__20_,r_57__19_,r_57__18_,r_57__17_,r_57__16_,r_57__15_,
  r_57__14_,r_57__13_,r_57__12_,r_57__11_,r_57__10_,r_57__9_,r_57__8_,r_57__7_,r_57__6_,
  r_57__5_,r_57__4_,r_57__3_,r_57__2_,r_57__1_,r_57__0_,r_58__63_,r_58__62_,
  r_58__61_,r_58__60_,r_58__59_,r_58__58_,r_58__57_,r_58__56_,r_58__55_,r_58__54_,
  r_58__53_,r_58__52_,r_58__51_,r_58__50_,r_58__49_,r_58__48_,r_58__47_,r_58__46_,
  r_58__45_,r_58__44_,r_58__43_,r_58__42_,r_58__41_,r_58__40_,r_58__39_,r_58__38_,
  r_58__37_,r_58__36_,r_58__35_,r_58__34_,r_58__33_,r_58__32_,r_58__31_,r_58__30_,
  r_58__29_,r_58__28_,r_58__27_,r_58__26_,r_58__25_,r_58__24_,r_58__23_,r_58__22_,
  r_58__21_,r_58__20_,r_58__19_,r_58__18_,r_58__17_,r_58__16_,r_58__15_,r_58__14_,
  r_58__13_,r_58__12_,r_58__11_,r_58__10_,r_58__9_,r_58__8_,r_58__7_,r_58__6_,r_58__5_,
  r_58__4_,r_58__3_,r_58__2_,r_58__1_,r_58__0_,r_59__63_,r_59__62_,r_59__61_,
  r_59__60_,r_59__59_,r_59__58_,r_59__57_,r_59__56_,r_59__55_,r_59__54_,r_59__53_,
  r_59__52_,r_59__51_,r_59__50_,r_59__49_,r_59__48_,r_59__47_,r_59__46_,r_59__45_,
  r_59__44_,r_59__43_,r_59__42_,r_59__41_,r_59__40_,r_59__39_,r_59__38_,r_59__37_,
  r_59__36_,r_59__35_,r_59__34_,r_59__33_,r_59__32_,r_59__31_,r_59__30_,r_59__29_,
  r_59__28_,r_59__27_,r_59__26_,r_59__25_,r_59__24_,r_59__23_,r_59__22_,r_59__21_,
  r_59__20_,r_59__19_,r_59__18_,r_59__17_,r_59__16_,r_59__15_,r_59__14_,r_59__13_,
  r_59__12_,r_59__11_,r_59__10_,r_59__9_,r_59__8_,r_59__7_,r_59__6_,r_59__5_,r_59__4_,
  r_59__3_,r_59__2_,r_59__1_,r_59__0_,r_60__63_,r_60__62_,r_60__61_,r_60__60_,
  r_60__59_,r_60__58_,r_60__57_,r_60__56_,r_60__55_,r_60__54_,r_60__53_,r_60__52_,
  r_60__51_,r_60__50_,r_60__49_,r_60__48_,r_60__47_,r_60__46_,r_60__45_,r_60__44_,
  r_60__43_,r_60__42_,r_60__41_,r_60__40_,r_60__39_,r_60__38_,r_60__37_,r_60__36_,
  r_60__35_,r_60__34_,r_60__33_,r_60__32_,r_60__31_,r_60__30_,r_60__29_,r_60__28_,
  r_60__27_,r_60__26_,r_60__25_,r_60__24_,r_60__23_,r_60__22_,r_60__21_,r_60__20_,
  r_60__19_,r_60__18_,r_60__17_,r_60__16_,r_60__15_,r_60__14_,r_60__13_,r_60__12_,
  r_60__11_,r_60__10_,r_60__9_,r_60__8_,r_60__7_,r_60__6_,r_60__5_,r_60__4_,r_60__3_,
  r_60__2_,r_60__1_,r_60__0_,r_61__63_,r_61__62_,r_61__61_,r_61__60_,r_61__59_,
  r_61__58_,r_61__57_,r_61__56_,r_61__55_,r_61__54_,r_61__53_,r_61__52_,r_61__51_,
  r_61__50_,r_61__49_,r_61__48_,r_61__47_,r_61__46_,r_61__45_,r_61__44_,r_61__43_,
  r_61__42_,r_61__41_,r_61__40_,r_61__39_,r_61__38_,r_61__37_,r_61__36_,r_61__35_,
  r_61__34_,r_61__33_,r_61__32_,r_61__31_,r_61__30_,r_61__29_,r_61__28_,r_61__27_,
  r_61__26_,r_61__25_,r_61__24_,r_61__23_,r_61__22_,r_61__21_,r_61__20_,r_61__19_,
  r_61__18_,r_61__17_,r_61__16_,r_61__15_,r_61__14_,r_61__13_,r_61__12_,r_61__11_,
  r_61__10_,r_61__9_,r_61__8_,r_61__7_,r_61__6_,r_61__5_,r_61__4_,r_61__3_,r_61__2_,
  r_61__1_,r_61__0_,r_62__63_,r_62__62_,r_62__61_,r_62__60_,r_62__59_,r_62__58_,
  r_62__57_,r_62__56_,r_62__55_,r_62__54_,r_62__53_,r_62__52_,r_62__51_,r_62__50_,
  r_62__49_,r_62__48_,r_62__47_,r_62__46_,r_62__45_,r_62__44_,r_62__43_,r_62__42_,
  r_62__41_,r_62__40_,r_62__39_,r_62__38_,r_62__37_,r_62__36_,r_62__35_,r_62__34_,
  r_62__33_,r_62__32_,r_62__31_,r_62__30_,r_62__29_,r_62__28_,r_62__27_,r_62__26_,
  r_62__25_,r_62__24_,r_62__23_,r_62__22_,r_62__21_,r_62__20_,r_62__19_,r_62__18_,
  r_62__17_,r_62__16_,r_62__15_,r_62__14_,r_62__13_,r_62__12_,r_62__11_,r_62__10_,
  r_62__9_,r_62__8_,r_62__7_,r_62__6_,r_62__5_,r_62__4_,r_62__3_,r_62__2_,r_62__1_,
  r_62__0_,r_63__63_,r_63__62_,r_63__61_,r_63__60_,r_63__59_,r_63__58_,r_63__57_,
  r_63__56_,r_63__55_,r_63__54_,r_63__53_,r_63__52_,r_63__51_,r_63__50_,r_63__49_,
  r_63__48_,r_63__47_,r_63__46_,r_63__45_,r_63__44_,r_63__43_,r_63__42_,r_63__41_,
  r_63__40_,r_63__39_,r_63__38_,r_63__37_,r_63__36_,r_63__35_,r_63__34_,r_63__33_,
  r_63__32_,r_63__31_,r_63__30_,r_63__29_,r_63__28_,r_63__27_,r_63__26_,r_63__25_,
  r_63__24_,r_63__23_,r_63__22_,r_63__21_,r_63__20_,r_63__19_,r_63__18_,r_63__17_,
  r_63__16_,r_63__15_,r_63__14_,r_63__13_,r_63__12_,r_63__11_,r_63__10_,r_63__9_,
  r_63__8_,r_63__7_,r_63__6_,r_63__5_,r_63__4_,r_63__3_,r_63__2_,r_63__1_,r_63__0_,
  r_64__63_,r_64__62_,r_64__61_,r_64__60_,r_64__59_,r_64__58_,r_64__57_,r_64__56_,
  r_64__55_,r_64__54_,r_64__53_,r_64__52_,r_64__51_,r_64__50_,r_64__49_,r_64__48_,
  r_64__47_,r_64__46_,r_64__45_,r_64__44_,r_64__43_,r_64__42_,r_64__41_,r_64__40_,
  r_64__39_,r_64__38_,r_64__37_,r_64__36_,r_64__35_,r_64__34_,r_64__33_,r_64__32_,
  r_64__31_,r_64__30_,r_64__29_,r_64__28_,r_64__27_,r_64__26_,r_64__25_,r_64__24_,
  r_64__23_,r_64__22_,r_64__21_,r_64__20_,r_64__19_,r_64__18_,r_64__17_,r_64__16_,
  r_64__15_,r_64__14_,r_64__13_,r_64__12_,r_64__11_,r_64__10_,r_64__9_,r_64__8_,
  r_64__7_,r_64__6_,r_64__5_,r_64__4_,r_64__3_,r_64__2_,r_64__1_,r_64__0_,r_65__63_,
  r_65__62_,r_65__61_,r_65__60_,r_65__59_,r_65__58_,r_65__57_,r_65__56_,r_65__55_,
  r_65__54_,r_65__53_,r_65__52_,r_65__51_,r_65__50_,r_65__49_,r_65__48_,r_65__47_,
  r_65__46_,r_65__45_,r_65__44_,r_65__43_,r_65__42_,r_65__41_,r_65__40_,r_65__39_,
  r_65__38_,r_65__37_,r_65__36_,r_65__35_,r_65__34_,r_65__33_,r_65__32_,r_65__31_,
  r_65__30_,r_65__29_,r_65__28_,r_65__27_,r_65__26_,r_65__25_,r_65__24_,r_65__23_,
  r_65__22_,r_65__21_,r_65__20_,r_65__19_,r_65__18_,r_65__17_,r_65__16_,r_65__15_,
  r_65__14_,r_65__13_,r_65__12_,r_65__11_,r_65__10_,r_65__9_,r_65__8_,r_65__7_,r_65__6_,
  r_65__5_,r_65__4_,r_65__3_,r_65__2_,r_65__1_,r_65__0_,r_66__63_,r_66__62_,
  r_66__61_,r_66__60_,r_66__59_,r_66__58_,r_66__57_,r_66__56_,r_66__55_,r_66__54_,
  r_66__53_,r_66__52_,r_66__51_,r_66__50_,r_66__49_,r_66__48_,r_66__47_,r_66__46_,
  r_66__45_,r_66__44_,r_66__43_,r_66__42_,r_66__41_,r_66__40_,r_66__39_,r_66__38_,
  r_66__37_,r_66__36_,r_66__35_,r_66__34_,r_66__33_,r_66__32_,r_66__31_,r_66__30_,
  r_66__29_,r_66__28_,r_66__27_,r_66__26_,r_66__25_,r_66__24_,r_66__23_,r_66__22_,
  r_66__21_,r_66__20_,r_66__19_,r_66__18_,r_66__17_,r_66__16_,r_66__15_,r_66__14_,
  r_66__13_,r_66__12_,r_66__11_,r_66__10_,r_66__9_,r_66__8_,r_66__7_,r_66__6_,r_66__5_,
  r_66__4_,r_66__3_,r_66__2_,r_66__1_,r_66__0_,r_67__63_,r_67__62_,r_67__61_,
  r_67__60_,r_67__59_,r_67__58_,r_67__57_,r_67__56_,r_67__55_,r_67__54_,r_67__53_,
  r_67__52_,r_67__51_,r_67__50_,r_67__49_,r_67__48_,r_67__47_,r_67__46_,r_67__45_,
  r_67__44_,r_67__43_,r_67__42_,r_67__41_,r_67__40_,r_67__39_,r_67__38_,r_67__37_,
  r_67__36_,r_67__35_,r_67__34_,r_67__33_,r_67__32_,r_67__31_,r_67__30_,r_67__29_,
  r_67__28_,r_67__27_,r_67__26_,r_67__25_,r_67__24_,r_67__23_,r_67__22_,r_67__21_,
  r_67__20_,r_67__19_,r_67__18_,r_67__17_,r_67__16_,r_67__15_,r_67__14_,r_67__13_,
  r_67__12_,r_67__11_,r_67__10_,r_67__9_,r_67__8_,r_67__7_,r_67__6_,r_67__5_,r_67__4_,
  r_67__3_,r_67__2_,r_67__1_,r_67__0_,r_68__63_,r_68__62_,r_68__61_,r_68__60_,
  r_68__59_,r_68__58_,r_68__57_,r_68__56_,r_68__55_,r_68__54_,r_68__53_,r_68__52_,
  r_68__51_,r_68__50_,r_68__49_,r_68__48_,r_68__47_,r_68__46_,r_68__45_,r_68__44_,
  r_68__43_,r_68__42_,r_68__41_,r_68__40_,r_68__39_,r_68__38_,r_68__37_,r_68__36_,
  r_68__35_,r_68__34_,r_68__33_,r_68__32_,r_68__31_,r_68__30_,r_68__29_,r_68__28_,
  r_68__27_,r_68__26_,r_68__25_,r_68__24_,r_68__23_,r_68__22_,r_68__21_,r_68__20_,
  r_68__19_,r_68__18_,r_68__17_,r_68__16_,r_68__15_,r_68__14_,r_68__13_,r_68__12_,
  r_68__11_,r_68__10_,r_68__9_,r_68__8_,r_68__7_,r_68__6_,r_68__5_,r_68__4_,r_68__3_,
  r_68__2_,r_68__1_,r_68__0_,r_69__63_,r_69__62_,r_69__61_,r_69__60_,r_69__59_,
  r_69__58_,r_69__57_,r_69__56_,r_69__55_,r_69__54_,r_69__53_,r_69__52_,r_69__51_,
  r_69__50_,r_69__49_,r_69__48_,r_69__47_,r_69__46_,r_69__45_,r_69__44_,r_69__43_,
  r_69__42_,r_69__41_,r_69__40_,r_69__39_,r_69__38_,r_69__37_,r_69__36_,r_69__35_,
  r_69__34_,r_69__33_,r_69__32_,r_69__31_,r_69__30_,r_69__29_,r_69__28_,r_69__27_,
  r_69__26_,r_69__25_,r_69__24_,r_69__23_,r_69__22_,r_69__21_,r_69__20_,r_69__19_,
  r_69__18_,r_69__17_,r_69__16_,r_69__15_,r_69__14_,r_69__13_,r_69__12_,r_69__11_,
  r_69__10_,r_69__9_,r_69__8_,r_69__7_,r_69__6_,r_69__5_,r_69__4_,r_69__3_,r_69__2_,
  r_69__1_,r_69__0_,r_70__63_,r_70__62_,r_70__61_,r_70__60_,r_70__59_,r_70__58_,
  r_70__57_,r_70__56_,r_70__55_,r_70__54_,r_70__53_,r_70__52_,r_70__51_,r_70__50_,
  r_70__49_,r_70__48_,r_70__47_,r_70__46_,r_70__45_,r_70__44_,r_70__43_,r_70__42_,
  r_70__41_,r_70__40_,r_70__39_,r_70__38_,r_70__37_,r_70__36_,r_70__35_,r_70__34_,
  r_70__33_,r_70__32_,r_70__31_,r_70__30_,r_70__29_,r_70__28_,r_70__27_,r_70__26_,
  r_70__25_,r_70__24_,r_70__23_,r_70__22_,r_70__21_,r_70__20_,r_70__19_,r_70__18_,
  r_70__17_,r_70__16_,r_70__15_,r_70__14_,r_70__13_,r_70__12_,r_70__11_,r_70__10_,
  r_70__9_,r_70__8_,r_70__7_,r_70__6_,r_70__5_,r_70__4_,r_70__3_,r_70__2_,r_70__1_,
  r_70__0_,r_71__63_,r_71__62_,r_71__61_,r_71__60_,r_71__59_,r_71__58_,r_71__57_,
  r_71__56_,r_71__55_,r_71__54_,r_71__53_,r_71__52_,r_71__51_,r_71__50_,r_71__49_,
  r_71__48_,r_71__47_,r_71__46_,r_71__45_,r_71__44_,r_71__43_,r_71__42_,r_71__41_,
  r_71__40_,r_71__39_,r_71__38_,r_71__37_,r_71__36_,r_71__35_,r_71__34_,r_71__33_,
  r_71__32_,r_71__31_,r_71__30_,r_71__29_,r_71__28_,r_71__27_,r_71__26_,r_71__25_,
  r_71__24_,r_71__23_,r_71__22_,r_71__21_,r_71__20_,r_71__19_,r_71__18_,r_71__17_,
  r_71__16_,r_71__15_,r_71__14_,r_71__13_,r_71__12_,r_71__11_,r_71__10_,r_71__9_,
  r_71__8_,r_71__7_,r_71__6_,r_71__5_,r_71__4_,r_71__3_,r_71__2_,r_71__1_,r_71__0_,
  r_72__63_,r_72__62_,r_72__61_,r_72__60_,r_72__59_,r_72__58_,r_72__57_,r_72__56_,
  r_72__55_,r_72__54_,r_72__53_,r_72__52_,r_72__51_,r_72__50_,r_72__49_,r_72__48_,
  r_72__47_,r_72__46_,r_72__45_,r_72__44_,r_72__43_,r_72__42_,r_72__41_,r_72__40_,
  r_72__39_,r_72__38_,r_72__37_,r_72__36_,r_72__35_,r_72__34_,r_72__33_,r_72__32_,
  r_72__31_,r_72__30_,r_72__29_,r_72__28_,r_72__27_,r_72__26_,r_72__25_,r_72__24_,
  r_72__23_,r_72__22_,r_72__21_,r_72__20_,r_72__19_,r_72__18_,r_72__17_,r_72__16_,
  r_72__15_,r_72__14_,r_72__13_,r_72__12_,r_72__11_,r_72__10_,r_72__9_,r_72__8_,
  r_72__7_,r_72__6_,r_72__5_,r_72__4_,r_72__3_,r_72__2_,r_72__1_,r_72__0_,r_73__63_,
  r_73__62_,r_73__61_,r_73__60_,r_73__59_,r_73__58_,r_73__57_,r_73__56_,r_73__55_,
  r_73__54_,r_73__53_,r_73__52_,r_73__51_,r_73__50_,r_73__49_,r_73__48_,r_73__47_,
  r_73__46_,r_73__45_,r_73__44_,r_73__43_,r_73__42_,r_73__41_,r_73__40_,r_73__39_,
  r_73__38_,r_73__37_,r_73__36_,r_73__35_,r_73__34_,r_73__33_,r_73__32_,r_73__31_,
  r_73__30_,r_73__29_,r_73__28_,r_73__27_,r_73__26_,r_73__25_,r_73__24_,r_73__23_,
  r_73__22_,r_73__21_,r_73__20_,r_73__19_,r_73__18_,r_73__17_,r_73__16_,r_73__15_,
  r_73__14_,r_73__13_,r_73__12_,r_73__11_,r_73__10_,r_73__9_,r_73__8_,r_73__7_,r_73__6_,
  r_73__5_,r_73__4_,r_73__3_,r_73__2_,r_73__1_,r_73__0_,r_74__63_,r_74__62_,
  r_74__61_,r_74__60_,r_74__59_,r_74__58_,r_74__57_,r_74__56_,r_74__55_,r_74__54_,
  r_74__53_,r_74__52_,r_74__51_,r_74__50_,r_74__49_,r_74__48_,r_74__47_,r_74__46_,
  r_74__45_,r_74__44_,r_74__43_,r_74__42_,r_74__41_,r_74__40_,r_74__39_,r_74__38_,
  r_74__37_,r_74__36_,r_74__35_,r_74__34_,r_74__33_,r_74__32_,r_74__31_,r_74__30_,
  r_74__29_,r_74__28_,r_74__27_,r_74__26_,r_74__25_,r_74__24_,r_74__23_,r_74__22_,
  r_74__21_,r_74__20_,r_74__19_,r_74__18_,r_74__17_,r_74__16_,r_74__15_,r_74__14_,
  r_74__13_,r_74__12_,r_74__11_,r_74__10_,r_74__9_,r_74__8_,r_74__7_,r_74__6_,r_74__5_,
  r_74__4_,r_74__3_,r_74__2_,r_74__1_,r_74__0_,r_75__63_,r_75__62_,r_75__61_,
  r_75__60_,r_75__59_,r_75__58_,r_75__57_,r_75__56_,r_75__55_,r_75__54_,r_75__53_,
  r_75__52_,r_75__51_,r_75__50_,r_75__49_,r_75__48_,r_75__47_,r_75__46_,r_75__45_,
  r_75__44_,r_75__43_,r_75__42_,r_75__41_,r_75__40_,r_75__39_,r_75__38_,r_75__37_,
  r_75__36_,r_75__35_,r_75__34_,r_75__33_,r_75__32_,r_75__31_,r_75__30_,r_75__29_,
  r_75__28_,r_75__27_,r_75__26_,r_75__25_,r_75__24_,r_75__23_,r_75__22_,r_75__21_,
  r_75__20_,r_75__19_,r_75__18_,r_75__17_,r_75__16_,r_75__15_,r_75__14_,r_75__13_,
  r_75__12_,r_75__11_,r_75__10_,r_75__9_,r_75__8_,r_75__7_,r_75__6_,r_75__5_,r_75__4_,
  r_75__3_,r_75__2_,r_75__1_,r_75__0_,r_76__63_,r_76__62_,r_76__61_,r_76__60_,
  r_76__59_,r_76__58_,r_76__57_,r_76__56_,r_76__55_,r_76__54_,r_76__53_,r_76__52_,
  r_76__51_,r_76__50_,r_76__49_,r_76__48_,r_76__47_,r_76__46_,r_76__45_,r_76__44_,
  r_76__43_,r_76__42_,r_76__41_,r_76__40_,r_76__39_,r_76__38_,r_76__37_,r_76__36_,
  r_76__35_,r_76__34_,r_76__33_,r_76__32_,r_76__31_,r_76__30_,r_76__29_,r_76__28_,
  r_76__27_,r_76__26_,r_76__25_,r_76__24_,r_76__23_,r_76__22_,r_76__21_,r_76__20_,
  r_76__19_,r_76__18_,r_76__17_,r_76__16_,r_76__15_,r_76__14_,r_76__13_,r_76__12_,
  r_76__11_,r_76__10_,r_76__9_,r_76__8_,r_76__7_,r_76__6_,r_76__5_,r_76__4_,r_76__3_,
  r_76__2_,r_76__1_,r_76__0_,r_77__63_,r_77__62_,r_77__61_,r_77__60_,r_77__59_,
  r_77__58_,r_77__57_,r_77__56_,r_77__55_,r_77__54_,r_77__53_,r_77__52_,r_77__51_,
  r_77__50_,r_77__49_,r_77__48_,r_77__47_,r_77__46_,r_77__45_,r_77__44_,r_77__43_,
  r_77__42_,r_77__41_,r_77__40_,r_77__39_,r_77__38_,r_77__37_,r_77__36_,r_77__35_,
  r_77__34_,r_77__33_,r_77__32_,r_77__31_,r_77__30_,r_77__29_,r_77__28_,r_77__27_,
  r_77__26_,r_77__25_,r_77__24_,r_77__23_,r_77__22_,r_77__21_,r_77__20_,r_77__19_,
  r_77__18_,r_77__17_,r_77__16_,r_77__15_,r_77__14_,r_77__13_,r_77__12_,r_77__11_,
  r_77__10_,r_77__9_,r_77__8_,r_77__7_,r_77__6_,r_77__5_,r_77__4_,r_77__3_,r_77__2_,
  r_77__1_,r_77__0_,r_78__63_,r_78__62_,r_78__61_,r_78__60_,r_78__59_,r_78__58_,
  r_78__57_,r_78__56_,r_78__55_,r_78__54_,r_78__53_,r_78__52_,r_78__51_,r_78__50_,
  r_78__49_,r_78__48_,r_78__47_,r_78__46_,r_78__45_,r_78__44_,r_78__43_,r_78__42_,
  r_78__41_,r_78__40_,r_78__39_,r_78__38_,r_78__37_,r_78__36_,r_78__35_,r_78__34_,
  r_78__33_,r_78__32_,r_78__31_,r_78__30_,r_78__29_,r_78__28_,r_78__27_,r_78__26_,
  r_78__25_,r_78__24_,r_78__23_,r_78__22_,r_78__21_,r_78__20_,r_78__19_,r_78__18_,
  r_78__17_,r_78__16_,r_78__15_,r_78__14_,r_78__13_,r_78__12_,r_78__11_,r_78__10_,
  r_78__9_,r_78__8_,r_78__7_,r_78__6_,r_78__5_,r_78__4_,r_78__3_,r_78__2_,r_78__1_,
  r_78__0_,r_79__63_,r_79__62_,r_79__61_,r_79__60_,r_79__59_,r_79__58_,r_79__57_,
  r_79__56_,r_79__55_,r_79__54_,r_79__53_,r_79__52_,r_79__51_,r_79__50_,r_79__49_,
  r_79__48_,r_79__47_,r_79__46_,r_79__45_,r_79__44_,r_79__43_,r_79__42_,r_79__41_,
  r_79__40_,r_79__39_,r_79__38_,r_79__37_,r_79__36_,r_79__35_,r_79__34_,r_79__33_,
  r_79__32_,r_79__31_,r_79__30_,r_79__29_,r_79__28_,r_79__27_,r_79__26_,r_79__25_,
  r_79__24_,r_79__23_,r_79__22_,r_79__21_,r_79__20_,r_79__19_,r_79__18_,r_79__17_,
  r_79__16_,r_79__15_,r_79__14_,r_79__13_,r_79__12_,r_79__11_,r_79__10_,r_79__9_,
  r_79__8_,r_79__7_,r_79__6_,r_79__5_,r_79__4_,r_79__3_,r_79__2_,r_79__1_,r_79__0_,
  r_80__63_,r_80__62_,r_80__61_,r_80__60_,r_80__59_,r_80__58_,r_80__57_,r_80__56_,
  r_80__55_,r_80__54_,r_80__53_,r_80__52_,r_80__51_,r_80__50_,r_80__49_,r_80__48_,
  r_80__47_,r_80__46_,r_80__45_,r_80__44_,r_80__43_,r_80__42_,r_80__41_,r_80__40_,
  r_80__39_,r_80__38_,r_80__37_,r_80__36_,r_80__35_,r_80__34_,r_80__33_,r_80__32_,
  r_80__31_,r_80__30_,r_80__29_,r_80__28_,r_80__27_,r_80__26_,r_80__25_,r_80__24_,
  r_80__23_,r_80__22_,r_80__21_,r_80__20_,r_80__19_,r_80__18_,r_80__17_,r_80__16_,
  r_80__15_,r_80__14_,r_80__13_,r_80__12_,r_80__11_,r_80__10_,r_80__9_,r_80__8_,
  r_80__7_,r_80__6_,r_80__5_,r_80__4_,r_80__3_,r_80__2_,r_80__1_,r_80__0_,r_81__63_,
  r_81__62_,r_81__61_,r_81__60_,r_81__59_,r_81__58_,r_81__57_,r_81__56_,r_81__55_,
  r_81__54_,r_81__53_,r_81__52_,r_81__51_,r_81__50_,r_81__49_,r_81__48_,r_81__47_,
  r_81__46_,r_81__45_,r_81__44_,r_81__43_,r_81__42_,r_81__41_,r_81__40_,r_81__39_,
  r_81__38_,r_81__37_,r_81__36_,r_81__35_,r_81__34_,r_81__33_,r_81__32_,r_81__31_,
  r_81__30_,r_81__29_,r_81__28_,r_81__27_,r_81__26_,r_81__25_,r_81__24_,r_81__23_,
  r_81__22_,r_81__21_,r_81__20_,r_81__19_,r_81__18_,r_81__17_,r_81__16_,r_81__15_,
  r_81__14_,r_81__13_,r_81__12_,r_81__11_,r_81__10_,r_81__9_,r_81__8_,r_81__7_,r_81__6_,
  r_81__5_,r_81__4_,r_81__3_,r_81__2_,r_81__1_,r_81__0_,r_82__63_,r_82__62_,
  r_82__61_,r_82__60_,r_82__59_,r_82__58_,r_82__57_,r_82__56_,r_82__55_,r_82__54_,
  r_82__53_,r_82__52_,r_82__51_,r_82__50_,r_82__49_,r_82__48_,r_82__47_,r_82__46_,
  r_82__45_,r_82__44_,r_82__43_,r_82__42_,r_82__41_,r_82__40_,r_82__39_,r_82__38_,
  r_82__37_,r_82__36_,r_82__35_,r_82__34_,r_82__33_,r_82__32_,r_82__31_,r_82__30_,
  r_82__29_,r_82__28_,r_82__27_,r_82__26_,r_82__25_,r_82__24_,r_82__23_,r_82__22_,
  r_82__21_,r_82__20_,r_82__19_,r_82__18_,r_82__17_,r_82__16_,r_82__15_,r_82__14_,
  r_82__13_,r_82__12_,r_82__11_,r_82__10_,r_82__9_,r_82__8_,r_82__7_,r_82__6_,r_82__5_,
  r_82__4_,r_82__3_,r_82__2_,r_82__1_,r_82__0_,r_83__63_,r_83__62_,r_83__61_,
  r_83__60_,r_83__59_,r_83__58_,r_83__57_,r_83__56_,r_83__55_,r_83__54_,r_83__53_,
  r_83__52_,r_83__51_,r_83__50_,r_83__49_,r_83__48_,r_83__47_,r_83__46_,r_83__45_,
  r_83__44_,r_83__43_,r_83__42_,r_83__41_,r_83__40_,r_83__39_,r_83__38_,r_83__37_,
  r_83__36_,r_83__35_,r_83__34_,r_83__33_,r_83__32_,r_83__31_,r_83__30_,r_83__29_,
  r_83__28_,r_83__27_,r_83__26_,r_83__25_,r_83__24_,r_83__23_,r_83__22_,r_83__21_,
  r_83__20_,r_83__19_,r_83__18_,r_83__17_,r_83__16_,r_83__15_,r_83__14_,r_83__13_,
  r_83__12_,r_83__11_,r_83__10_,r_83__9_,r_83__8_,r_83__7_,r_83__6_,r_83__5_,r_83__4_,
  r_83__3_,r_83__2_,r_83__1_,r_83__0_,r_84__63_,r_84__62_,r_84__61_,r_84__60_,
  r_84__59_,r_84__58_,r_84__57_,r_84__56_,r_84__55_,r_84__54_,r_84__53_,r_84__52_,
  r_84__51_,r_84__50_,r_84__49_,r_84__48_,r_84__47_,r_84__46_,r_84__45_,r_84__44_,
  r_84__43_,r_84__42_,r_84__41_,r_84__40_,r_84__39_,r_84__38_,r_84__37_,r_84__36_,
  r_84__35_,r_84__34_,r_84__33_,r_84__32_,r_84__31_,r_84__30_,r_84__29_,r_84__28_,
  r_84__27_,r_84__26_,r_84__25_,r_84__24_,r_84__23_,r_84__22_,r_84__21_,r_84__20_,
  r_84__19_,r_84__18_,r_84__17_,r_84__16_,r_84__15_,r_84__14_,r_84__13_,r_84__12_,
  r_84__11_,r_84__10_,r_84__9_,r_84__8_,r_84__7_,r_84__6_,r_84__5_,r_84__4_,r_84__3_,
  r_84__2_,r_84__1_,r_84__0_,r_85__63_,r_85__62_,r_85__61_,r_85__60_,r_85__59_,
  r_85__58_,r_85__57_,r_85__56_,r_85__55_,r_85__54_,r_85__53_,r_85__52_,r_85__51_,
  r_85__50_,r_85__49_,r_85__48_,r_85__47_,r_85__46_,r_85__45_,r_85__44_,r_85__43_,
  r_85__42_,r_85__41_,r_85__40_,r_85__39_,r_85__38_,r_85__37_,r_85__36_,r_85__35_,
  r_85__34_,r_85__33_,r_85__32_,r_85__31_,r_85__30_,r_85__29_,r_85__28_,r_85__27_,
  r_85__26_,r_85__25_,r_85__24_,r_85__23_,r_85__22_,r_85__21_,r_85__20_,r_85__19_,
  r_85__18_,r_85__17_,r_85__16_,r_85__15_,r_85__14_,r_85__13_,r_85__12_,r_85__11_,
  r_85__10_,r_85__9_,r_85__8_,r_85__7_,r_85__6_,r_85__5_,r_85__4_,r_85__3_,r_85__2_,
  r_85__1_,r_85__0_,r_86__63_,r_86__62_,r_86__61_,r_86__60_,r_86__59_,r_86__58_,
  r_86__57_,r_86__56_,r_86__55_,r_86__54_,r_86__53_,r_86__52_,r_86__51_,r_86__50_,
  r_86__49_,r_86__48_,r_86__47_,r_86__46_,r_86__45_,r_86__44_,r_86__43_,r_86__42_,
  r_86__41_,r_86__40_,r_86__39_,r_86__38_,r_86__37_,r_86__36_,r_86__35_,r_86__34_,
  r_86__33_,r_86__32_,r_86__31_,r_86__30_,r_86__29_,r_86__28_,r_86__27_,r_86__26_,
  r_86__25_,r_86__24_,r_86__23_,r_86__22_,r_86__21_,r_86__20_,r_86__19_,r_86__18_,
  r_86__17_,r_86__16_,r_86__15_,r_86__14_,r_86__13_,r_86__12_,r_86__11_,r_86__10_,
  r_86__9_,r_86__8_,r_86__7_,r_86__6_,r_86__5_,r_86__4_,r_86__3_,r_86__2_,r_86__1_,
  r_86__0_,r_87__63_,r_87__62_,r_87__61_,r_87__60_,r_87__59_,r_87__58_,r_87__57_,
  r_87__56_,r_87__55_,r_87__54_,r_87__53_,r_87__52_,r_87__51_,r_87__50_,r_87__49_,
  r_87__48_,r_87__47_,r_87__46_,r_87__45_,r_87__44_,r_87__43_,r_87__42_,r_87__41_,
  r_87__40_,r_87__39_,r_87__38_,r_87__37_,r_87__36_,r_87__35_,r_87__34_,r_87__33_,
  r_87__32_,r_87__31_,r_87__30_,r_87__29_,r_87__28_,r_87__27_,r_87__26_,r_87__25_,
  r_87__24_,r_87__23_,r_87__22_,r_87__21_,r_87__20_,r_87__19_,r_87__18_,r_87__17_,
  r_87__16_,r_87__15_,r_87__14_,r_87__13_,r_87__12_,r_87__11_,r_87__10_,r_87__9_,
  r_87__8_,r_87__7_,r_87__6_,r_87__5_,r_87__4_,r_87__3_,r_87__2_,r_87__1_,r_87__0_,
  r_88__63_,r_88__62_,r_88__61_,r_88__60_,r_88__59_,r_88__58_,r_88__57_,r_88__56_,
  r_88__55_,r_88__54_,r_88__53_,r_88__52_,r_88__51_,r_88__50_,r_88__49_,r_88__48_,
  r_88__47_,r_88__46_,r_88__45_,r_88__44_,r_88__43_,r_88__42_,r_88__41_,r_88__40_,
  r_88__39_,r_88__38_,r_88__37_,r_88__36_,r_88__35_,r_88__34_,r_88__33_,r_88__32_,
  r_88__31_,r_88__30_,r_88__29_,r_88__28_,r_88__27_,r_88__26_,r_88__25_,r_88__24_,
  r_88__23_,r_88__22_,r_88__21_,r_88__20_,r_88__19_,r_88__18_,r_88__17_,r_88__16_,
  r_88__15_,r_88__14_,r_88__13_,r_88__12_,r_88__11_,r_88__10_,r_88__9_,r_88__8_,
  r_88__7_,r_88__6_,r_88__5_,r_88__4_,r_88__3_,r_88__2_,r_88__1_,r_88__0_,r_89__63_,
  r_89__62_,r_89__61_,r_89__60_,r_89__59_,r_89__58_,r_89__57_,r_89__56_,r_89__55_,
  r_89__54_,r_89__53_,r_89__52_,r_89__51_,r_89__50_,r_89__49_,r_89__48_,r_89__47_,
  r_89__46_,r_89__45_,r_89__44_,r_89__43_,r_89__42_,r_89__41_,r_89__40_,r_89__39_,
  r_89__38_,r_89__37_,r_89__36_,r_89__35_,r_89__34_,r_89__33_,r_89__32_,r_89__31_,
  r_89__30_,r_89__29_,r_89__28_,r_89__27_,r_89__26_,r_89__25_,r_89__24_,r_89__23_,
  r_89__22_,r_89__21_,r_89__20_,r_89__19_,r_89__18_,r_89__17_,r_89__16_,r_89__15_,
  r_89__14_,r_89__13_,r_89__12_,r_89__11_,r_89__10_,r_89__9_,r_89__8_,r_89__7_,r_89__6_,
  r_89__5_,r_89__4_,r_89__3_,r_89__2_,r_89__1_,r_89__0_,r_90__63_,r_90__62_,
  r_90__61_,r_90__60_,r_90__59_,r_90__58_,r_90__57_,r_90__56_,r_90__55_,r_90__54_,
  r_90__53_,r_90__52_,r_90__51_,r_90__50_,r_90__49_,r_90__48_,r_90__47_,r_90__46_,
  r_90__45_,r_90__44_,r_90__43_,r_90__42_,r_90__41_,r_90__40_,r_90__39_,r_90__38_,
  r_90__37_,r_90__36_,r_90__35_,r_90__34_,r_90__33_,r_90__32_,r_90__31_,r_90__30_,
  r_90__29_,r_90__28_,r_90__27_,r_90__26_,r_90__25_,r_90__24_,r_90__23_,r_90__22_,
  r_90__21_,r_90__20_,r_90__19_,r_90__18_,r_90__17_,r_90__16_,r_90__15_,r_90__14_,
  r_90__13_,r_90__12_,r_90__11_,r_90__10_,r_90__9_,r_90__8_,r_90__7_,r_90__6_,r_90__5_,
  r_90__4_,r_90__3_,r_90__2_,r_90__1_,r_90__0_,r_91__63_,r_91__62_,r_91__61_,
  r_91__60_,r_91__59_,r_91__58_,r_91__57_,r_91__56_,r_91__55_,r_91__54_,r_91__53_,
  r_91__52_,r_91__51_,r_91__50_,r_91__49_,r_91__48_,r_91__47_,r_91__46_,r_91__45_,
  r_91__44_,r_91__43_,r_91__42_,r_91__41_,r_91__40_,r_91__39_,r_91__38_,r_91__37_,
  r_91__36_,r_91__35_,r_91__34_,r_91__33_,r_91__32_,r_91__31_,r_91__30_,r_91__29_,
  r_91__28_,r_91__27_,r_91__26_,r_91__25_,r_91__24_,r_91__23_,r_91__22_,r_91__21_,
  r_91__20_,r_91__19_,r_91__18_,r_91__17_,r_91__16_,r_91__15_,r_91__14_,r_91__13_,
  r_91__12_,r_91__11_,r_91__10_,r_91__9_,r_91__8_,r_91__7_,r_91__6_,r_91__5_,r_91__4_,
  r_91__3_,r_91__2_,r_91__1_,r_91__0_,r_92__63_,r_92__62_,r_92__61_,r_92__60_,
  r_92__59_,r_92__58_,r_92__57_,r_92__56_,r_92__55_,r_92__54_,r_92__53_,r_92__52_,
  r_92__51_,r_92__50_,r_92__49_,r_92__48_,r_92__47_,r_92__46_,r_92__45_,r_92__44_,
  r_92__43_,r_92__42_,r_92__41_,r_92__40_,r_92__39_,r_92__38_,r_92__37_,r_92__36_,
  r_92__35_,r_92__34_,r_92__33_,r_92__32_,r_92__31_,r_92__30_,r_92__29_,r_92__28_,
  r_92__27_,r_92__26_,r_92__25_,r_92__24_,r_92__23_,r_92__22_,r_92__21_,r_92__20_,
  r_92__19_,r_92__18_,r_92__17_,r_92__16_,r_92__15_,r_92__14_,r_92__13_,r_92__12_,
  r_92__11_,r_92__10_,r_92__9_,r_92__8_,r_92__7_,r_92__6_,r_92__5_,r_92__4_,r_92__3_,
  r_92__2_,r_92__1_,r_92__0_,r_93__63_,r_93__62_,r_93__61_,r_93__60_,r_93__59_,
  r_93__58_,r_93__57_,r_93__56_,r_93__55_,r_93__54_,r_93__53_,r_93__52_,r_93__51_,
  r_93__50_,r_93__49_,r_93__48_,r_93__47_,r_93__46_,r_93__45_,r_93__44_,r_93__43_,
  r_93__42_,r_93__41_,r_93__40_,r_93__39_,r_93__38_,r_93__37_,r_93__36_,r_93__35_,
  r_93__34_,r_93__33_,r_93__32_,r_93__31_,r_93__30_,r_93__29_,r_93__28_,r_93__27_,
  r_93__26_,r_93__25_,r_93__24_,r_93__23_,r_93__22_,r_93__21_,r_93__20_,r_93__19_,
  r_93__18_,r_93__17_,r_93__16_,r_93__15_,r_93__14_,r_93__13_,r_93__12_,r_93__11_,
  r_93__10_,r_93__9_,r_93__8_,r_93__7_,r_93__6_,r_93__5_,r_93__4_,r_93__3_,r_93__2_,
  r_93__1_,r_93__0_,r_94__63_,r_94__62_,r_94__61_,r_94__60_,r_94__59_,r_94__58_,
  r_94__57_,r_94__56_,r_94__55_,r_94__54_,r_94__53_,r_94__52_,r_94__51_,r_94__50_,
  r_94__49_,r_94__48_,r_94__47_,r_94__46_,r_94__45_,r_94__44_,r_94__43_,r_94__42_,
  r_94__41_,r_94__40_,r_94__39_,r_94__38_,r_94__37_,r_94__36_,r_94__35_,r_94__34_,
  r_94__33_,r_94__32_,r_94__31_,r_94__30_,r_94__29_,r_94__28_,r_94__27_,r_94__26_,
  r_94__25_,r_94__24_,r_94__23_,r_94__22_,r_94__21_,r_94__20_,r_94__19_,r_94__18_,
  r_94__17_,r_94__16_,r_94__15_,r_94__14_,r_94__13_,r_94__12_,r_94__11_,r_94__10_,
  r_94__9_,r_94__8_,r_94__7_,r_94__6_,r_94__5_,r_94__4_,r_94__3_,r_94__2_,r_94__1_,
  r_94__0_,r_95__63_,r_95__62_,r_95__61_,r_95__60_,r_95__59_,r_95__58_,r_95__57_,
  r_95__56_,r_95__55_,r_95__54_,r_95__53_,r_95__52_,r_95__51_,r_95__50_,r_95__49_,
  r_95__48_,r_95__47_,r_95__46_,r_95__45_,r_95__44_,r_95__43_,r_95__42_,r_95__41_,
  r_95__40_,r_95__39_,r_95__38_,r_95__37_,r_95__36_,r_95__35_,r_95__34_,r_95__33_,
  r_95__32_,r_95__31_,r_95__30_,r_95__29_,r_95__28_,r_95__27_,r_95__26_,r_95__25_,
  r_95__24_,r_95__23_,r_95__22_,r_95__21_,r_95__20_,r_95__19_,r_95__18_,r_95__17_,
  r_95__16_,r_95__15_,r_95__14_,r_95__13_,r_95__12_,r_95__11_,r_95__10_,r_95__9_,
  r_95__8_,r_95__7_,r_95__6_,r_95__5_,r_95__4_,r_95__3_,r_95__2_,r_95__1_,r_95__0_,
  r_96__63_,r_96__62_,r_96__61_,r_96__60_,r_96__59_,r_96__58_,r_96__57_,r_96__56_,
  r_96__55_,r_96__54_,r_96__53_,r_96__52_,r_96__51_,r_96__50_,r_96__49_,r_96__48_,
  r_96__47_,r_96__46_,r_96__45_,r_96__44_,r_96__43_,r_96__42_,r_96__41_,r_96__40_,
  r_96__39_,r_96__38_,r_96__37_,r_96__36_,r_96__35_,r_96__34_,r_96__33_,r_96__32_,
  r_96__31_,r_96__30_,r_96__29_,r_96__28_,r_96__27_,r_96__26_,r_96__25_,r_96__24_,
  r_96__23_,r_96__22_,r_96__21_,r_96__20_,r_96__19_,r_96__18_,r_96__17_,r_96__16_,
  r_96__15_,r_96__14_,r_96__13_,r_96__12_,r_96__11_,r_96__10_,r_96__9_,r_96__8_,
  r_96__7_,r_96__6_,r_96__5_,r_96__4_,r_96__3_,r_96__2_,r_96__1_,r_96__0_,r_97__63_,
  r_97__62_,r_97__61_,r_97__60_,r_97__59_,r_97__58_,r_97__57_,r_97__56_,r_97__55_,
  r_97__54_,r_97__53_,r_97__52_,r_97__51_,r_97__50_,r_97__49_,r_97__48_,r_97__47_,
  r_97__46_,r_97__45_,r_97__44_,r_97__43_,r_97__42_,r_97__41_,r_97__40_,r_97__39_,
  r_97__38_,r_97__37_,r_97__36_,r_97__35_,r_97__34_,r_97__33_,r_97__32_,r_97__31_,
  r_97__30_,r_97__29_,r_97__28_,r_97__27_,r_97__26_,r_97__25_,r_97__24_,r_97__23_,
  r_97__22_,r_97__21_,r_97__20_,r_97__19_,r_97__18_,r_97__17_,r_97__16_,r_97__15_,
  r_97__14_,r_97__13_,r_97__12_,r_97__11_,r_97__10_,r_97__9_,r_97__8_,r_97__7_,r_97__6_,
  r_97__5_,r_97__4_,r_97__3_,r_97__2_,r_97__1_,r_97__0_,r_98__63_,r_98__62_,
  r_98__61_,r_98__60_,r_98__59_,r_98__58_,r_98__57_,r_98__56_,r_98__55_,r_98__54_,
  r_98__53_,r_98__52_,r_98__51_,r_98__50_,r_98__49_,r_98__48_,r_98__47_,r_98__46_,
  r_98__45_,r_98__44_,r_98__43_,r_98__42_,r_98__41_,r_98__40_,r_98__39_,r_98__38_,
  r_98__37_,r_98__36_,r_98__35_,r_98__34_,r_98__33_,r_98__32_,r_98__31_,r_98__30_,
  r_98__29_,r_98__28_,r_98__27_,r_98__26_,r_98__25_,r_98__24_,r_98__23_,r_98__22_,
  r_98__21_,r_98__20_,r_98__19_,r_98__18_,r_98__17_,r_98__16_,r_98__15_,r_98__14_,
  r_98__13_,r_98__12_,r_98__11_,r_98__10_,r_98__9_,r_98__8_,r_98__7_,r_98__6_,r_98__5_,
  r_98__4_,r_98__3_,r_98__2_,r_98__1_,r_98__0_,r_99__63_,r_99__62_,r_99__61_,
  r_99__60_,r_99__59_,r_99__58_,r_99__57_,r_99__56_,r_99__55_,r_99__54_,r_99__53_,
  r_99__52_,r_99__51_,r_99__50_,r_99__49_,r_99__48_,r_99__47_,r_99__46_,r_99__45_,
  r_99__44_,r_99__43_,r_99__42_,r_99__41_,r_99__40_,r_99__39_,r_99__38_,r_99__37_,
  r_99__36_,r_99__35_,r_99__34_,r_99__33_,r_99__32_,r_99__31_,r_99__30_,r_99__29_,
  r_99__28_,r_99__27_,r_99__26_,r_99__25_,r_99__24_,r_99__23_,r_99__22_,r_99__21_,
  r_99__20_,r_99__19_,r_99__18_,r_99__17_,r_99__16_,r_99__15_,r_99__14_,r_99__13_,
  r_99__12_,r_99__11_,r_99__10_,r_99__9_,r_99__8_,r_99__7_,r_99__6_,r_99__5_,r_99__4_,
  r_99__3_,r_99__2_,r_99__1_,r_99__0_,r_100__63_,r_100__62_,r_100__61_,r_100__60_,
  r_100__59_,r_100__58_,r_100__57_,r_100__56_,r_100__55_,r_100__54_,r_100__53_,
  r_100__52_,r_100__51_,r_100__50_,r_100__49_,r_100__48_,r_100__47_,r_100__46_,
  r_100__45_,r_100__44_,r_100__43_,r_100__42_,r_100__41_,r_100__40_,r_100__39_,r_100__38_,
  r_100__37_,r_100__36_,r_100__35_,r_100__34_,r_100__33_,r_100__32_,r_100__31_,
  r_100__30_,r_100__29_,r_100__28_,r_100__27_,r_100__26_,r_100__25_,r_100__24_,
  r_100__23_,r_100__22_,r_100__21_,r_100__20_,r_100__19_,r_100__18_,r_100__17_,
  r_100__16_,r_100__15_,r_100__14_,r_100__13_,r_100__12_,r_100__11_,r_100__10_,r_100__9_,
  r_100__8_,r_100__7_,r_100__6_,r_100__5_,r_100__4_,r_100__3_,r_100__2_,r_100__1_,
  r_100__0_,r_101__63_,r_101__62_,r_101__61_,r_101__60_,r_101__59_,r_101__58_,
  r_101__57_,r_101__56_,r_101__55_,r_101__54_,r_101__53_,r_101__52_,r_101__51_,
  r_101__50_,r_101__49_,r_101__48_,r_101__47_,r_101__46_,r_101__45_,r_101__44_,r_101__43_,
  r_101__42_,r_101__41_,r_101__40_,r_101__39_,r_101__38_,r_101__37_,r_101__36_,
  r_101__35_,r_101__34_,r_101__33_,r_101__32_,r_101__31_,r_101__30_,r_101__29_,
  r_101__28_,r_101__27_,r_101__26_,r_101__25_,r_101__24_,r_101__23_,r_101__22_,
  r_101__21_,r_101__20_,r_101__19_,r_101__18_,r_101__17_,r_101__16_,r_101__15_,r_101__14_,
  r_101__13_,r_101__12_,r_101__11_,r_101__10_,r_101__9_,r_101__8_,r_101__7_,
  r_101__6_,r_101__5_,r_101__4_,r_101__3_,r_101__2_,r_101__1_,r_101__0_,r_102__63_,
  r_102__62_,r_102__61_,r_102__60_,r_102__59_,r_102__58_,r_102__57_,r_102__56_,
  r_102__55_,r_102__54_,r_102__53_,r_102__52_,r_102__51_,r_102__50_,r_102__49_,r_102__48_,
  r_102__47_,r_102__46_,r_102__45_,r_102__44_,r_102__43_,r_102__42_,r_102__41_,
  r_102__40_,r_102__39_,r_102__38_,r_102__37_,r_102__36_,r_102__35_,r_102__34_,
  r_102__33_,r_102__32_,r_102__31_,r_102__30_,r_102__29_,r_102__28_,r_102__27_,r_102__26_,
  r_102__25_,r_102__24_,r_102__23_,r_102__22_,r_102__21_,r_102__20_,r_102__19_,
  r_102__18_,r_102__17_,r_102__16_,r_102__15_,r_102__14_,r_102__13_,r_102__12_,
  r_102__11_,r_102__10_,r_102__9_,r_102__8_,r_102__7_,r_102__6_,r_102__5_,r_102__4_,
  r_102__3_,r_102__2_,r_102__1_,r_102__0_,r_103__63_,r_103__62_,r_103__61_,r_103__60_,
  r_103__59_,r_103__58_,r_103__57_,r_103__56_,r_103__55_,r_103__54_,r_103__53_,
  r_103__52_,r_103__51_,r_103__50_,r_103__49_,r_103__48_,r_103__47_,r_103__46_,
  r_103__45_,r_103__44_,r_103__43_,r_103__42_,r_103__41_,r_103__40_,r_103__39_,
  r_103__38_,r_103__37_,r_103__36_,r_103__35_,r_103__34_,r_103__33_,r_103__32_,r_103__31_,
  r_103__30_,r_103__29_,r_103__28_,r_103__27_,r_103__26_,r_103__25_,r_103__24_,
  r_103__23_,r_103__22_,r_103__21_,r_103__20_,r_103__19_,r_103__18_,r_103__17_,
  r_103__16_,r_103__15_,r_103__14_,r_103__13_,r_103__12_,r_103__11_,r_103__10_,r_103__9_,
  r_103__8_,r_103__7_,r_103__6_,r_103__5_,r_103__4_,r_103__3_,r_103__2_,r_103__1_,
  r_103__0_,r_104__63_,r_104__62_,r_104__61_,r_104__60_,r_104__59_,r_104__58_,
  r_104__57_,r_104__56_,r_104__55_,r_104__54_,r_104__53_,r_104__52_,r_104__51_,
  r_104__50_,r_104__49_,r_104__48_,r_104__47_,r_104__46_,r_104__45_,r_104__44_,
  r_104__43_,r_104__42_,r_104__41_,r_104__40_,r_104__39_,r_104__38_,r_104__37_,r_104__36_,
  r_104__35_,r_104__34_,r_104__33_,r_104__32_,r_104__31_,r_104__30_,r_104__29_,
  r_104__28_,r_104__27_,r_104__26_,r_104__25_,r_104__24_,r_104__23_,r_104__22_,
  r_104__21_,r_104__20_,r_104__19_,r_104__18_,r_104__17_,r_104__16_,r_104__15_,r_104__14_,
  r_104__13_,r_104__12_,r_104__11_,r_104__10_,r_104__9_,r_104__8_,r_104__7_,
  r_104__6_,r_104__5_,r_104__4_,r_104__3_,r_104__2_,r_104__1_,r_104__0_,r_105__63_,
  r_105__62_,r_105__61_,r_105__60_,r_105__59_,r_105__58_,r_105__57_,r_105__56_,
  r_105__55_,r_105__54_,r_105__53_,r_105__52_,r_105__51_,r_105__50_,r_105__49_,r_105__48_,
  r_105__47_,r_105__46_,r_105__45_,r_105__44_,r_105__43_,r_105__42_,r_105__41_,
  r_105__40_,r_105__39_,r_105__38_,r_105__37_,r_105__36_,r_105__35_,r_105__34_,
  r_105__33_,r_105__32_,r_105__31_,r_105__30_,r_105__29_,r_105__28_,r_105__27_,
  r_105__26_,r_105__25_,r_105__24_,r_105__23_,r_105__22_,r_105__21_,r_105__20_,r_105__19_,
  r_105__18_,r_105__17_,r_105__16_,r_105__15_,r_105__14_,r_105__13_,r_105__12_,
  r_105__11_,r_105__10_,r_105__9_,r_105__8_,r_105__7_,r_105__6_,r_105__5_,r_105__4_,
  r_105__3_,r_105__2_,r_105__1_,r_105__0_,r_106__63_,r_106__62_,r_106__61_,
  r_106__60_,r_106__59_,r_106__58_,r_106__57_,r_106__56_,r_106__55_,r_106__54_,r_106__53_,
  r_106__52_,r_106__51_,r_106__50_,r_106__49_,r_106__48_,r_106__47_,r_106__46_,
  r_106__45_,r_106__44_,r_106__43_,r_106__42_,r_106__41_,r_106__40_,r_106__39_,
  r_106__38_,r_106__37_,r_106__36_,r_106__35_,r_106__34_,r_106__33_,r_106__32_,
  r_106__31_,r_106__30_,r_106__29_,r_106__28_,r_106__27_,r_106__26_,r_106__25_,r_106__24_,
  r_106__23_,r_106__22_,r_106__21_,r_106__20_,r_106__19_,r_106__18_,r_106__17_,
  r_106__16_,r_106__15_,r_106__14_,r_106__13_,r_106__12_,r_106__11_,r_106__10_,
  r_106__9_,r_106__8_,r_106__7_,r_106__6_,r_106__5_,r_106__4_,r_106__3_,r_106__2_,
  r_106__1_,r_106__0_,r_107__63_,r_107__62_,r_107__61_,r_107__60_,r_107__59_,r_107__58_,
  r_107__57_,r_107__56_,r_107__55_,r_107__54_,r_107__53_,r_107__52_,r_107__51_,
  r_107__50_,r_107__49_,r_107__48_,r_107__47_,r_107__46_,r_107__45_,r_107__44_,
  r_107__43_,r_107__42_,r_107__41_,r_107__40_,r_107__39_,r_107__38_,r_107__37_,r_107__36_,
  r_107__35_,r_107__34_,r_107__33_,r_107__32_,r_107__31_,r_107__30_,r_107__29_,
  r_107__28_,r_107__27_,r_107__26_,r_107__25_,r_107__24_,r_107__23_,r_107__22_,
  r_107__21_,r_107__20_,r_107__19_,r_107__18_,r_107__17_,r_107__16_,r_107__15_,
  r_107__14_,r_107__13_,r_107__12_,r_107__11_,r_107__10_,r_107__9_,r_107__8_,r_107__7_,
  r_107__6_,r_107__5_,r_107__4_,r_107__3_,r_107__2_,r_107__1_,r_107__0_,r_108__63_,
  r_108__62_,r_108__61_,r_108__60_,r_108__59_,r_108__58_,r_108__57_,r_108__56_,
  r_108__55_,r_108__54_,r_108__53_,r_108__52_,r_108__51_,r_108__50_,r_108__49_,
  r_108__48_,r_108__47_,r_108__46_,r_108__45_,r_108__44_,r_108__43_,r_108__42_,r_108__41_,
  r_108__40_,r_108__39_,r_108__38_,r_108__37_,r_108__36_,r_108__35_,r_108__34_,
  r_108__33_,r_108__32_,r_108__31_,r_108__30_,r_108__29_,r_108__28_,r_108__27_,
  r_108__26_,r_108__25_,r_108__24_,r_108__23_,r_108__22_,r_108__21_,r_108__20_,
  r_108__19_,r_108__18_,r_108__17_,r_108__16_,r_108__15_,r_108__14_,r_108__13_,r_108__12_,
  r_108__11_,r_108__10_,r_108__9_,r_108__8_,r_108__7_,r_108__6_,r_108__5_,r_108__4_,
  r_108__3_,r_108__2_,r_108__1_,r_108__0_,r_109__63_,r_109__62_,r_109__61_,
  r_109__60_,r_109__59_,r_109__58_,r_109__57_,r_109__56_,r_109__55_,r_109__54_,
  r_109__53_,r_109__52_,r_109__51_,r_109__50_,r_109__49_,r_109__48_,r_109__47_,r_109__46_,
  r_109__45_,r_109__44_,r_109__43_,r_109__42_,r_109__41_,r_109__40_,r_109__39_,
  r_109__38_,r_109__37_,r_109__36_,r_109__35_,r_109__34_,r_109__33_,r_109__32_,
  r_109__31_,r_109__30_,r_109__29_,r_109__28_,r_109__27_,r_109__26_,r_109__25_,r_109__24_,
  r_109__23_,r_109__22_,r_109__21_,r_109__20_,r_109__19_,r_109__18_,r_109__17_,
  r_109__16_,r_109__15_,r_109__14_,r_109__13_,r_109__12_,r_109__11_,r_109__10_,
  r_109__9_,r_109__8_,r_109__7_,r_109__6_,r_109__5_,r_109__4_,r_109__3_,r_109__2_,
  r_109__1_,r_109__0_,r_110__63_,r_110__62_,r_110__61_,r_110__60_,r_110__59_,r_110__58_,
  r_110__57_,r_110__56_,r_110__55_,r_110__54_,r_110__53_,r_110__52_,r_110__51_,
  r_110__50_,r_110__49_,r_110__48_,r_110__47_,r_110__46_,r_110__45_,r_110__44_,
  r_110__43_,r_110__42_,r_110__41_,r_110__40_,r_110__39_,r_110__38_,r_110__37_,
  r_110__36_,r_110__35_,r_110__34_,r_110__33_,r_110__32_,r_110__31_,r_110__30_,r_110__29_,
  r_110__28_,r_110__27_,r_110__26_,r_110__25_,r_110__24_,r_110__23_,r_110__22_,
  r_110__21_,r_110__20_,r_110__19_,r_110__18_,r_110__17_,r_110__16_,r_110__15_,
  r_110__14_,r_110__13_,r_110__12_,r_110__11_,r_110__10_,r_110__9_,r_110__8_,r_110__7_,
  r_110__6_,r_110__5_,r_110__4_,r_110__3_,r_110__2_,r_110__1_,r_110__0_,r_111__63_,
  r_111__62_,r_111__61_,r_111__60_,r_111__59_,r_111__58_,r_111__57_,r_111__56_,
  r_111__55_,r_111__54_,r_111__53_,r_111__52_,r_111__51_,r_111__50_,r_111__49_,
  r_111__48_,r_111__47_,r_111__46_,r_111__45_,r_111__44_,r_111__43_,r_111__42_,
  r_111__41_,r_111__40_,r_111__39_,r_111__38_,r_111__37_,r_111__36_,r_111__35_,r_111__34_,
  r_111__33_,r_111__32_,r_111__31_,r_111__30_,r_111__29_,r_111__28_,r_111__27_,
  r_111__26_,r_111__25_,r_111__24_,r_111__23_,r_111__22_,r_111__21_,r_111__20_,
  r_111__19_,r_111__18_,r_111__17_,r_111__16_,r_111__15_,r_111__14_,r_111__13_,r_111__12_,
  r_111__11_,r_111__10_,r_111__9_,r_111__8_,r_111__7_,r_111__6_,r_111__5_,
  r_111__4_,r_111__3_,r_111__2_,r_111__1_,r_111__0_,r_112__63_,r_112__62_,r_112__61_,
  r_112__60_,r_112__59_,r_112__58_,r_112__57_,r_112__56_,r_112__55_,r_112__54_,
  r_112__53_,r_112__52_,r_112__51_,r_112__50_,r_112__49_,r_112__48_,r_112__47_,r_112__46_,
  r_112__45_,r_112__44_,r_112__43_,r_112__42_,r_112__41_,r_112__40_,r_112__39_,
  r_112__38_,r_112__37_,r_112__36_,r_112__35_,r_112__34_,r_112__33_,r_112__32_,
  r_112__31_,r_112__30_,r_112__29_,r_112__28_,r_112__27_,r_112__26_,r_112__25_,
  r_112__24_,r_112__23_,r_112__22_,r_112__21_,r_112__20_,r_112__19_,r_112__18_,r_112__17_,
  r_112__16_,r_112__15_,r_112__14_,r_112__13_,r_112__12_,r_112__11_,r_112__10_,
  r_112__9_,r_112__8_,r_112__7_,r_112__6_,r_112__5_,r_112__4_,r_112__3_,r_112__2_,
  r_112__1_,r_112__0_,r_113__63_,r_113__62_,r_113__61_,r_113__60_,r_113__59_,
  r_113__58_,r_113__57_,r_113__56_,r_113__55_,r_113__54_,r_113__53_,r_113__52_,r_113__51_,
  r_113__50_,r_113__49_,r_113__48_,r_113__47_,r_113__46_,r_113__45_,r_113__44_,
  r_113__43_,r_113__42_,r_113__41_,r_113__40_,r_113__39_,r_113__38_,r_113__37_,
  r_113__36_,r_113__35_,r_113__34_,r_113__33_,r_113__32_,r_113__31_,r_113__30_,
  r_113__29_,r_113__28_,r_113__27_,r_113__26_,r_113__25_,r_113__24_,r_113__23_,r_113__22_,
  r_113__21_,r_113__20_,r_113__19_,r_113__18_,r_113__17_,r_113__16_,r_113__15_,
  r_113__14_,r_113__13_,r_113__12_,r_113__11_,r_113__10_,r_113__9_,r_113__8_,r_113__7_,
  r_113__6_,r_113__5_,r_113__4_,r_113__3_,r_113__2_,r_113__1_,r_113__0_,
  r_114__63_,r_114__62_,r_114__61_,r_114__60_,r_114__59_,r_114__58_,r_114__57_,r_114__56_,
  r_114__55_,r_114__54_,r_114__53_,r_114__52_,r_114__51_,r_114__50_,r_114__49_,
  r_114__48_,r_114__47_,r_114__46_,r_114__45_,r_114__44_,r_114__43_,r_114__42_,
  r_114__41_,r_114__40_,r_114__39_,r_114__38_,r_114__37_,r_114__36_,r_114__35_,r_114__34_,
  r_114__33_,r_114__32_,r_114__31_,r_114__30_,r_114__29_,r_114__28_,r_114__27_,
  r_114__26_,r_114__25_,r_114__24_,r_114__23_,r_114__22_,r_114__21_,r_114__20_,
  r_114__19_,r_114__18_,r_114__17_,r_114__16_,r_114__15_,r_114__14_,r_114__13_,
  r_114__12_,r_114__11_,r_114__10_,r_114__9_,r_114__8_,r_114__7_,r_114__6_,r_114__5_,
  r_114__4_,r_114__3_,r_114__2_,r_114__1_,r_114__0_,r_115__63_,r_115__62_,r_115__61_,
  r_115__60_,r_115__59_,r_115__58_,r_115__57_,r_115__56_,r_115__55_,r_115__54_,
  r_115__53_,r_115__52_,r_115__51_,r_115__50_,r_115__49_,r_115__48_,r_115__47_,
  r_115__46_,r_115__45_,r_115__44_,r_115__43_,r_115__42_,r_115__41_,r_115__40_,r_115__39_,
  r_115__38_,r_115__37_,r_115__36_,r_115__35_,r_115__34_,r_115__33_,r_115__32_,
  r_115__31_,r_115__30_,r_115__29_,r_115__28_,r_115__27_,r_115__26_,r_115__25_,
  r_115__24_,r_115__23_,r_115__22_,r_115__21_,r_115__20_,r_115__19_,r_115__18_,
  r_115__17_,r_115__16_,r_115__15_,r_115__14_,r_115__13_,r_115__12_,r_115__11_,r_115__10_,
  r_115__9_,r_115__8_,r_115__7_,r_115__6_,r_115__5_,r_115__4_,r_115__3_,r_115__2_,
  r_115__1_,r_115__0_,r_116__63_,r_116__62_,r_116__61_,r_116__60_,r_116__59_,
  r_116__58_,r_116__57_,r_116__56_,r_116__55_,r_116__54_,r_116__53_,r_116__52_,
  r_116__51_,r_116__50_,r_116__49_,r_116__48_,r_116__47_,r_116__46_,r_116__45_,r_116__44_,
  r_116__43_,r_116__42_,r_116__41_,r_116__40_,r_116__39_,r_116__38_,r_116__37_,
  r_116__36_,r_116__35_,r_116__34_,r_116__33_,r_116__32_,r_116__31_,r_116__30_,
  r_116__29_,r_116__28_,r_116__27_,r_116__26_,r_116__25_,r_116__24_,r_116__23_,r_116__22_,
  r_116__21_,r_116__20_,r_116__19_,r_116__18_,r_116__17_,r_116__16_,r_116__15_,
  r_116__14_,r_116__13_,r_116__12_,r_116__11_,r_116__10_,r_116__9_,r_116__8_,
  r_116__7_,r_116__6_,r_116__5_,r_116__4_,r_116__3_,r_116__2_,r_116__1_,r_116__0_,
  r_117__63_,r_117__62_,r_117__61_,r_117__60_,r_117__59_,r_117__58_,r_117__57_,r_117__56_,
  r_117__55_,r_117__54_,r_117__53_,r_117__52_,r_117__51_,r_117__50_,r_117__49_,
  r_117__48_,r_117__47_,r_117__46_,r_117__45_,r_117__44_,r_117__43_,r_117__42_,
  r_117__41_,r_117__40_,r_117__39_,r_117__38_,r_117__37_,r_117__36_,r_117__35_,
  r_117__34_,r_117__33_,r_117__32_,r_117__31_,r_117__30_,r_117__29_,r_117__28_,r_117__27_,
  r_117__26_,r_117__25_,r_117__24_,r_117__23_,r_117__22_,r_117__21_,r_117__20_,
  r_117__19_,r_117__18_,r_117__17_,r_117__16_,r_117__15_,r_117__14_,r_117__13_,
  r_117__12_,r_117__11_,r_117__10_,r_117__9_,r_117__8_,r_117__7_,r_117__6_,r_117__5_,
  r_117__4_,r_117__3_,r_117__2_,r_117__1_,r_117__0_,r_118__63_,r_118__62_,r_118__61_,
  r_118__60_,r_118__59_,r_118__58_,r_118__57_,r_118__56_,r_118__55_,r_118__54_,
  r_118__53_,r_118__52_,r_118__51_,r_118__50_,r_118__49_,r_118__48_,r_118__47_,
  r_118__46_,r_118__45_,r_118__44_,r_118__43_,r_118__42_,r_118__41_,r_118__40_,
  r_118__39_,r_118__38_,r_118__37_,r_118__36_,r_118__35_,r_118__34_,r_118__33_,r_118__32_,
  r_118__31_,r_118__30_,r_118__29_,r_118__28_,r_118__27_,r_118__26_,r_118__25_,
  r_118__24_,r_118__23_,r_118__22_,r_118__21_,r_118__20_,r_118__19_,r_118__18_,
  r_118__17_,r_118__16_,r_118__15_,r_118__14_,r_118__13_,r_118__12_,r_118__11_,r_118__10_,
  r_118__9_,r_118__8_,r_118__7_,r_118__6_,r_118__5_,r_118__4_,r_118__3_,r_118__2_,
  r_118__1_,r_118__0_,r_119__63_,r_119__62_,r_119__61_,r_119__60_,r_119__59_,
  r_119__58_,r_119__57_,r_119__56_,r_119__55_,r_119__54_,r_119__53_,r_119__52_,
  r_119__51_,r_119__50_,r_119__49_,r_119__48_,r_119__47_,r_119__46_,r_119__45_,r_119__44_,
  r_119__43_,r_119__42_,r_119__41_,r_119__40_,r_119__39_,r_119__38_,r_119__37_,
  r_119__36_,r_119__35_,r_119__34_,r_119__33_,r_119__32_,r_119__31_,r_119__30_,
  r_119__29_,r_119__28_,r_119__27_,r_119__26_,r_119__25_,r_119__24_,r_119__23_,
  r_119__22_,r_119__21_,r_119__20_,r_119__19_,r_119__18_,r_119__17_,r_119__16_,r_119__15_,
  r_119__14_,r_119__13_,r_119__12_,r_119__11_,r_119__10_,r_119__9_,r_119__8_,
  r_119__7_,r_119__6_,r_119__5_,r_119__4_,r_119__3_,r_119__2_,r_119__1_,r_119__0_,
  r_120__63_,r_120__62_,r_120__61_,r_120__60_,r_120__59_,r_120__58_,r_120__57_,
  r_120__56_,r_120__55_,r_120__54_,r_120__53_,r_120__52_,r_120__51_,r_120__50_,r_120__49_,
  r_120__48_,r_120__47_,r_120__46_,r_120__45_,r_120__44_,r_120__43_,r_120__42_,
  r_120__41_,r_120__40_,r_120__39_,r_120__38_,r_120__37_,r_120__36_,r_120__35_,
  r_120__34_,r_120__33_,r_120__32_,r_120__31_,r_120__30_,r_120__29_,r_120__28_,
  r_120__27_,r_120__26_,r_120__25_,r_120__24_,r_120__23_,r_120__22_,r_120__21_,r_120__20_,
  r_120__19_,r_120__18_,r_120__17_,r_120__16_,r_120__15_,r_120__14_,r_120__13_,
  r_120__12_,r_120__11_,r_120__10_,r_120__9_,r_120__8_,r_120__7_,r_120__6_,r_120__5_,
  r_120__4_,r_120__3_,r_120__2_,r_120__1_,r_120__0_,r_121__63_,r_121__62_,
  r_121__61_,r_121__60_,r_121__59_,r_121__58_,r_121__57_,r_121__56_,r_121__55_,r_121__54_,
  r_121__53_,r_121__52_,r_121__51_,r_121__50_,r_121__49_,r_121__48_,r_121__47_,
  r_121__46_,r_121__45_,r_121__44_,r_121__43_,r_121__42_,r_121__41_,r_121__40_,
  r_121__39_,r_121__38_,r_121__37_,r_121__36_,r_121__35_,r_121__34_,r_121__33_,r_121__32_,
  r_121__31_,r_121__30_,r_121__29_,r_121__28_,r_121__27_,r_121__26_,r_121__25_,
  r_121__24_,r_121__23_,r_121__22_,r_121__21_,r_121__20_,r_121__19_,r_121__18_,
  r_121__17_,r_121__16_,r_121__15_,r_121__14_,r_121__13_,r_121__12_,r_121__11_,
  r_121__10_,r_121__9_,r_121__8_,r_121__7_,r_121__6_,r_121__5_,r_121__4_,r_121__3_,
  r_121__2_,r_121__1_,r_121__0_,r_122__63_,r_122__62_,r_122__61_,r_122__60_,r_122__59_,
  r_122__58_,r_122__57_,r_122__56_,r_122__55_,r_122__54_,r_122__53_,r_122__52_,
  r_122__51_,r_122__50_,r_122__49_,r_122__48_,r_122__47_,r_122__46_,r_122__45_,
  r_122__44_,r_122__43_,r_122__42_,r_122__41_,r_122__40_,r_122__39_,r_122__38_,r_122__37_,
  r_122__36_,r_122__35_,r_122__34_,r_122__33_,r_122__32_,r_122__31_,r_122__30_,
  r_122__29_,r_122__28_,r_122__27_,r_122__26_,r_122__25_,r_122__24_,r_122__23_,
  r_122__22_,r_122__21_,r_122__20_,r_122__19_,r_122__18_,r_122__17_,r_122__16_,
  r_122__15_,r_122__14_,r_122__13_,r_122__12_,r_122__11_,r_122__10_,r_122__9_,r_122__8_,
  r_122__7_,r_122__6_,r_122__5_,r_122__4_,r_122__3_,r_122__2_,r_122__1_,r_122__0_,
  r_123__63_,r_123__62_,r_123__61_,r_123__60_,r_123__59_,r_123__58_,r_123__57_,
  r_123__56_,r_123__55_,r_123__54_,r_123__53_,r_123__52_,r_123__51_,r_123__50_,
  r_123__49_,r_123__48_,r_123__47_,r_123__46_,r_123__45_,r_123__44_,r_123__43_,r_123__42_,
  r_123__41_,r_123__40_,r_123__39_,r_123__38_,r_123__37_,r_123__36_,r_123__35_,
  r_123__34_,r_123__33_,r_123__32_,r_123__31_,r_123__30_,r_123__29_,r_123__28_,
  r_123__27_,r_123__26_,r_123__25_,r_123__24_,r_123__23_,r_123__22_,r_123__21_,r_123__20_,
  r_123__19_,r_123__18_,r_123__17_,r_123__16_,r_123__15_,r_123__14_,r_123__13_,
  r_123__12_,r_123__11_,r_123__10_,r_123__9_,r_123__8_,r_123__7_,r_123__6_,r_123__5_,
  r_123__4_,r_123__3_,r_123__2_,r_123__1_,r_123__0_,r_124__63_,r_124__62_,
  r_124__61_,r_124__60_,r_124__59_,r_124__58_,r_124__57_,r_124__56_,r_124__55_,r_124__54_,
  r_124__53_,r_124__52_,r_124__51_,r_124__50_,r_124__49_,r_124__48_,r_124__47_,
  r_124__46_,r_124__45_,r_124__44_,r_124__43_,r_124__42_,r_124__41_,r_124__40_,
  r_124__39_,r_124__38_,r_124__37_,r_124__36_,r_124__35_,r_124__34_,r_124__33_,
  r_124__32_,r_124__31_,r_124__30_,r_124__29_,r_124__28_,r_124__27_,r_124__26_,r_124__25_,
  r_124__24_,r_124__23_,r_124__22_,r_124__21_,r_124__20_,r_124__19_,r_124__18_,
  r_124__17_,r_124__16_,r_124__15_,r_124__14_,r_124__13_,r_124__12_,r_124__11_,
  r_124__10_,r_124__9_,r_124__8_,r_124__7_,r_124__6_,r_124__5_,r_124__4_,r_124__3_,
  r_124__2_,r_124__1_,r_124__0_,r_125__63_,r_125__62_,r_125__61_,r_125__60_,r_125__59_,
  r_125__58_,r_125__57_,r_125__56_,r_125__55_,r_125__54_,r_125__53_,r_125__52_,
  r_125__51_,r_125__50_,r_125__49_,r_125__48_,r_125__47_,r_125__46_,r_125__45_,
  r_125__44_,r_125__43_,r_125__42_,r_125__41_,r_125__40_,r_125__39_,r_125__38_,
  r_125__37_,r_125__36_,r_125__35_,r_125__34_,r_125__33_,r_125__32_,r_125__31_,r_125__30_,
  r_125__29_,r_125__28_,r_125__27_,r_125__26_,r_125__25_,r_125__24_,r_125__23_,
  r_125__22_,r_125__21_,r_125__20_,r_125__19_,r_125__18_,r_125__17_,r_125__16_,
  r_125__15_,r_125__14_,r_125__13_,r_125__12_,r_125__11_,r_125__10_,r_125__9_,r_125__8_,
  r_125__7_,r_125__6_,r_125__5_,r_125__4_,r_125__3_,r_125__2_,r_125__1_,r_125__0_,
  r_126__63_,r_126__62_,r_126__61_,r_126__60_,r_126__59_,r_126__58_,r_126__57_,
  r_126__56_,r_126__55_,r_126__54_,r_126__53_,r_126__52_,r_126__51_,r_126__50_,
  r_126__49_,r_126__48_,r_126__47_,r_126__46_,r_126__45_,r_126__44_,r_126__43_,r_126__42_,
  r_126__41_,r_126__40_,r_126__39_,r_126__38_,r_126__37_,r_126__36_,r_126__35_,
  r_126__34_,r_126__33_,r_126__32_,r_126__31_,r_126__30_,r_126__29_,r_126__28_,
  r_126__27_,r_126__26_,r_126__25_,r_126__24_,r_126__23_,r_126__22_,r_126__21_,
  r_126__20_,r_126__19_,r_126__18_,r_126__17_,r_126__16_,r_126__15_,r_126__14_,r_126__13_,
  r_126__12_,r_126__11_,r_126__10_,r_126__9_,r_126__8_,r_126__7_,r_126__6_,
  r_126__5_,r_126__4_,r_126__3_,r_126__2_,r_126__1_,r_126__0_,r_127__63_,r_127__62_,
  r_127__61_,r_127__60_,r_127__59_,r_127__58_,r_127__57_,r_127__56_,r_127__55_,
  r_127__54_,r_127__53_,r_127__52_,r_127__51_,r_127__50_,r_127__49_,r_127__48_,r_127__47_,
  r_127__46_,r_127__45_,r_127__44_,r_127__43_,r_127__42_,r_127__41_,r_127__40_,
  r_127__39_,r_127__38_,r_127__37_,r_127__36_,r_127__35_,r_127__34_,r_127__33_,
  r_127__32_,r_127__31_,r_127__30_,r_127__29_,r_127__28_,r_127__27_,r_127__26_,
  r_127__25_,r_127__24_,r_127__23_,r_127__22_,r_127__21_,r_127__20_,r_127__19_,r_127__18_,
  r_127__17_,r_127__16_,r_127__15_,r_127__14_,r_127__13_,r_127__12_,r_127__11_,
  r_127__10_,r_127__9_,r_127__8_,r_127__7_,r_127__6_,r_127__5_,r_127__4_,r_127__3_,
  r_127__2_,r_127__1_,r_127__0_,r_128__63_,r_128__62_,r_128__61_,r_128__60_,
  r_128__59_,r_128__58_,r_128__57_,r_128__56_,r_128__55_,r_128__54_,r_128__53_,r_128__52_,
  r_128__51_,r_128__50_,r_128__49_,r_128__48_,r_128__47_,r_128__46_,r_128__45_,
  r_128__44_,r_128__43_,r_128__42_,r_128__41_,r_128__40_,r_128__39_,r_128__38_,
  r_128__37_,r_128__36_,r_128__35_,r_128__34_,r_128__33_,r_128__32_,r_128__31_,r_128__30_,
  r_128__29_,r_128__28_,r_128__27_,r_128__26_,r_128__25_,r_128__24_,r_128__23_,
  r_128__22_,r_128__21_,r_128__20_,r_128__19_,r_128__18_,r_128__17_,r_128__16_,
  r_128__15_,r_128__14_,r_128__13_,r_128__12_,r_128__11_,r_128__10_,r_128__9_,r_128__8_,
  r_128__7_,r_128__6_,r_128__5_,r_128__4_,r_128__3_,r_128__2_,r_128__1_,r_128__0_,
  r_129__63_,r_129__62_,r_129__61_,r_129__60_,r_129__59_,r_129__58_,r_129__57_,
  r_129__56_,r_129__55_,r_129__54_,r_129__53_,r_129__52_,r_129__51_,r_129__50_,
  r_129__49_,r_129__48_,r_129__47_,r_129__46_,r_129__45_,r_129__44_,r_129__43_,
  r_129__42_,r_129__41_,r_129__40_,r_129__39_,r_129__38_,r_129__37_,r_129__36_,r_129__35_,
  r_129__34_,r_129__33_,r_129__32_,r_129__31_,r_129__30_,r_129__29_,r_129__28_,
  r_129__27_,r_129__26_,r_129__25_,r_129__24_,r_129__23_,r_129__22_,r_129__21_,
  r_129__20_,r_129__19_,r_129__18_,r_129__17_,r_129__16_,r_129__15_,r_129__14_,
  r_129__13_,r_129__12_,r_129__11_,r_129__10_,r_129__9_,r_129__8_,r_129__7_,r_129__6_,
  r_129__5_,r_129__4_,r_129__3_,r_129__2_,r_129__1_,r_129__0_,r_130__63_,r_130__62_,
  r_130__61_,r_130__60_,r_130__59_,r_130__58_,r_130__57_,r_130__56_,r_130__55_,
  r_130__54_,r_130__53_,r_130__52_,r_130__51_,r_130__50_,r_130__49_,r_130__48_,
  r_130__47_,r_130__46_,r_130__45_,r_130__44_,r_130__43_,r_130__42_,r_130__41_,r_130__40_,
  r_130__39_,r_130__38_,r_130__37_,r_130__36_,r_130__35_,r_130__34_,r_130__33_,
  r_130__32_,r_130__31_,r_130__30_,r_130__29_,r_130__28_,r_130__27_,r_130__26_,
  r_130__25_,r_130__24_,r_130__23_,r_130__22_,r_130__21_,r_130__20_,r_130__19_,r_130__18_,
  r_130__17_,r_130__16_,r_130__15_,r_130__14_,r_130__13_,r_130__12_,r_130__11_,
  r_130__10_,r_130__9_,r_130__8_,r_130__7_,r_130__6_,r_130__5_,r_130__4_,r_130__3_,
  r_130__2_,r_130__1_,r_130__0_,r_131__63_,r_131__62_,r_131__61_,r_131__60_,
  r_131__59_,r_131__58_,r_131__57_,r_131__56_,r_131__55_,r_131__54_,r_131__53_,r_131__52_,
  r_131__51_,r_131__50_,r_131__49_,r_131__48_,r_131__47_,r_131__46_,r_131__45_,
  r_131__44_,r_131__43_,r_131__42_,r_131__41_,r_131__40_,r_131__39_,r_131__38_,
  r_131__37_,r_131__36_,r_131__35_,r_131__34_,r_131__33_,r_131__32_,r_131__31_,
  r_131__30_,r_131__29_,r_131__28_,r_131__27_,r_131__26_,r_131__25_,r_131__24_,r_131__23_,
  r_131__22_,r_131__21_,r_131__20_,r_131__19_,r_131__18_,r_131__17_,r_131__16_,
  r_131__15_,r_131__14_,r_131__13_,r_131__12_,r_131__11_,r_131__10_,r_131__9_,
  r_131__8_,r_131__7_,r_131__6_,r_131__5_,r_131__4_,r_131__3_,r_131__2_,r_131__1_,
  r_131__0_,r_132__63_,r_132__62_,r_132__61_,r_132__60_,r_132__59_,r_132__58_,r_132__57_,
  r_132__56_,r_132__55_,r_132__54_,r_132__53_,r_132__52_,r_132__51_,r_132__50_,
  r_132__49_,r_132__48_,r_132__47_,r_132__46_,r_132__45_,r_132__44_,r_132__43_,
  r_132__42_,r_132__41_,r_132__40_,r_132__39_,r_132__38_,r_132__37_,r_132__36_,
  r_132__35_,r_132__34_,r_132__33_,r_132__32_,r_132__31_,r_132__30_,r_132__29_,r_132__28_,
  r_132__27_,r_132__26_,r_132__25_,r_132__24_,r_132__23_,r_132__22_,r_132__21_,
  r_132__20_,r_132__19_,r_132__18_,r_132__17_,r_132__16_,r_132__15_,r_132__14_,
  r_132__13_,r_132__12_,r_132__11_,r_132__10_,r_132__9_,r_132__8_,r_132__7_,r_132__6_,
  r_132__5_,r_132__4_,r_132__3_,r_132__2_,r_132__1_,r_132__0_,r_133__63_,r_133__62_,
  r_133__61_,r_133__60_,r_133__59_,r_133__58_,r_133__57_,r_133__56_,r_133__55_,
  r_133__54_,r_133__53_,r_133__52_,r_133__51_,r_133__50_,r_133__49_,r_133__48_,
  r_133__47_,r_133__46_,r_133__45_,r_133__44_,r_133__43_,r_133__42_,r_133__41_,r_133__40_,
  r_133__39_,r_133__38_,r_133__37_,r_133__36_,r_133__35_,r_133__34_,r_133__33_,
  r_133__32_,r_133__31_,r_133__30_,r_133__29_,r_133__28_,r_133__27_,r_133__26_,
  r_133__25_,r_133__24_,r_133__23_,r_133__22_,r_133__21_,r_133__20_,r_133__19_,
  r_133__18_,r_133__17_,r_133__16_,r_133__15_,r_133__14_,r_133__13_,r_133__12_,r_133__11_,
  r_133__10_,r_133__9_,r_133__8_,r_133__7_,r_133__6_,r_133__5_,r_133__4_,r_133__3_,
  r_133__2_,r_133__1_,r_133__0_,r_134__63_,r_134__62_,r_134__61_,r_134__60_,
  r_134__59_,r_134__58_,r_134__57_,r_134__56_,r_134__55_,r_134__54_,r_134__53_,
  r_134__52_,r_134__51_,r_134__50_,r_134__49_,r_134__48_,r_134__47_,r_134__46_,r_134__45_,
  r_134__44_,r_134__43_,r_134__42_,r_134__41_,r_134__40_,r_134__39_,r_134__38_,
  r_134__37_,r_134__36_,r_134__35_,r_134__34_,r_134__33_,r_134__32_,r_134__31_,
  r_134__30_,r_134__29_,r_134__28_,r_134__27_,r_134__26_,r_134__25_,r_134__24_,
  r_134__23_,r_134__22_,r_134__21_,r_134__20_,r_134__19_,r_134__18_,r_134__17_,r_134__16_,
  r_134__15_,r_134__14_,r_134__13_,r_134__12_,r_134__11_,r_134__10_,r_134__9_,
  r_134__8_,r_134__7_,r_134__6_,r_134__5_,r_134__4_,r_134__3_,r_134__2_,r_134__1_,
  r_134__0_,r_135__63_,r_135__62_,r_135__61_,r_135__60_,r_135__59_,r_135__58_,
  r_135__57_,r_135__56_,r_135__55_,r_135__54_,r_135__53_,r_135__52_,r_135__51_,r_135__50_,
  r_135__49_,r_135__48_,r_135__47_,r_135__46_,r_135__45_,r_135__44_,r_135__43_,
  r_135__42_,r_135__41_,r_135__40_,r_135__39_,r_135__38_,r_135__37_,r_135__36_,
  r_135__35_,r_135__34_,r_135__33_,r_135__32_,r_135__31_,r_135__30_,r_135__29_,r_135__28_,
  r_135__27_,r_135__26_,r_135__25_,r_135__24_,r_135__23_,r_135__22_,r_135__21_,
  r_135__20_,r_135__19_,r_135__18_,r_135__17_,r_135__16_,r_135__15_,r_135__14_,
  r_135__13_,r_135__12_,r_135__11_,r_135__10_,r_135__9_,r_135__8_,r_135__7_,r_135__6_,
  r_135__5_,r_135__4_,r_135__3_,r_135__2_,r_135__1_,r_135__0_,r_136__63_,r_136__62_,
  r_136__61_,r_136__60_,r_136__59_,r_136__58_,r_136__57_,r_136__56_,r_136__55_,
  r_136__54_,r_136__53_,r_136__52_,r_136__51_,r_136__50_,r_136__49_,r_136__48_,
  r_136__47_,r_136__46_,r_136__45_,r_136__44_,r_136__43_,r_136__42_,r_136__41_,
  r_136__40_,r_136__39_,r_136__38_,r_136__37_,r_136__36_,r_136__35_,r_136__34_,r_136__33_,
  r_136__32_,r_136__31_,r_136__30_,r_136__29_,r_136__28_,r_136__27_,r_136__26_,
  r_136__25_,r_136__24_,r_136__23_,r_136__22_,r_136__21_,r_136__20_,r_136__19_,
  r_136__18_,r_136__17_,r_136__16_,r_136__15_,r_136__14_,r_136__13_,r_136__12_,
  r_136__11_,r_136__10_,r_136__9_,r_136__8_,r_136__7_,r_136__6_,r_136__5_,r_136__4_,
  r_136__3_,r_136__2_,r_136__1_,r_136__0_,r_137__63_,r_137__62_,r_137__61_,r_137__60_,
  r_137__59_,r_137__58_,r_137__57_,r_137__56_,r_137__55_,r_137__54_,r_137__53_,
  r_137__52_,r_137__51_,r_137__50_,r_137__49_,r_137__48_,r_137__47_,r_137__46_,
  r_137__45_,r_137__44_,r_137__43_,r_137__42_,r_137__41_,r_137__40_,r_137__39_,r_137__38_,
  r_137__37_,r_137__36_,r_137__35_,r_137__34_,r_137__33_,r_137__32_,r_137__31_,
  r_137__30_,r_137__29_,r_137__28_,r_137__27_,r_137__26_,r_137__25_,r_137__24_,
  r_137__23_,r_137__22_,r_137__21_,r_137__20_,r_137__19_,r_137__18_,r_137__17_,r_137__16_,
  r_137__15_,r_137__14_,r_137__13_,r_137__12_,r_137__11_,r_137__10_,r_137__9_,
  r_137__8_,r_137__7_,r_137__6_,r_137__5_,r_137__4_,r_137__3_,r_137__2_,r_137__1_,
  r_137__0_,r_138__63_,r_138__62_,r_138__61_,r_138__60_,r_138__59_,r_138__58_,
  r_138__57_,r_138__56_,r_138__55_,r_138__54_,r_138__53_,r_138__52_,r_138__51_,r_138__50_,
  r_138__49_,r_138__48_,r_138__47_,r_138__46_,r_138__45_,r_138__44_,r_138__43_,
  r_138__42_,r_138__41_,r_138__40_,r_138__39_,r_138__38_,r_138__37_,r_138__36_,
  r_138__35_,r_138__34_,r_138__33_,r_138__32_,r_138__31_,r_138__30_,r_138__29_,
  r_138__28_,r_138__27_,r_138__26_,r_138__25_,r_138__24_,r_138__23_,r_138__22_,r_138__21_,
  r_138__20_,r_138__19_,r_138__18_,r_138__17_,r_138__16_,r_138__15_,r_138__14_,
  r_138__13_,r_138__12_,r_138__11_,r_138__10_,r_138__9_,r_138__8_,r_138__7_,r_138__6_,
  r_138__5_,r_138__4_,r_138__3_,r_138__2_,r_138__1_,r_138__0_,r_139__63_,
  r_139__62_,r_139__61_,r_139__60_,r_139__59_,r_139__58_,r_139__57_,r_139__56_,r_139__55_,
  r_139__54_,r_139__53_,r_139__52_,r_139__51_,r_139__50_,r_139__49_,r_139__48_,
  r_139__47_,r_139__46_,r_139__45_,r_139__44_,r_139__43_,r_139__42_,r_139__41_,
  r_139__40_,r_139__39_,r_139__38_,r_139__37_,r_139__36_,r_139__35_,r_139__34_,
  r_139__33_,r_139__32_,r_139__31_,r_139__30_,r_139__29_,r_139__28_,r_139__27_,r_139__26_,
  r_139__25_,r_139__24_,r_139__23_,r_139__22_,r_139__21_,r_139__20_,r_139__19_,
  r_139__18_,r_139__17_,r_139__16_,r_139__15_,r_139__14_,r_139__13_,r_139__12_,
  r_139__11_,r_139__10_,r_139__9_,r_139__8_,r_139__7_,r_139__6_,r_139__5_,r_139__4_,
  r_139__3_,r_139__2_,r_139__1_,r_139__0_,r_140__63_,r_140__62_,r_140__61_,r_140__60_,
  r_140__59_,r_140__58_,r_140__57_,r_140__56_,r_140__55_,r_140__54_,r_140__53_,
  r_140__52_,r_140__51_,r_140__50_,r_140__49_,r_140__48_,r_140__47_,r_140__46_,
  r_140__45_,r_140__44_,r_140__43_,r_140__42_,r_140__41_,r_140__40_,r_140__39_,r_140__38_,
  r_140__37_,r_140__36_,r_140__35_,r_140__34_,r_140__33_,r_140__32_,r_140__31_,
  r_140__30_,r_140__29_,r_140__28_,r_140__27_,r_140__26_,r_140__25_,r_140__24_,
  r_140__23_,r_140__22_,r_140__21_,r_140__20_,r_140__19_,r_140__18_,r_140__17_,
  r_140__16_,r_140__15_,r_140__14_,r_140__13_,r_140__12_,r_140__11_,r_140__10_,r_140__9_,
  r_140__8_,r_140__7_,r_140__6_,r_140__5_,r_140__4_,r_140__3_,r_140__2_,r_140__1_,
  r_140__0_,r_141__63_,r_141__62_,r_141__61_,r_141__60_,r_141__59_,r_141__58_,
  r_141__57_,r_141__56_,r_141__55_,r_141__54_,r_141__53_,r_141__52_,r_141__51_,
  r_141__50_,r_141__49_,r_141__48_,r_141__47_,r_141__46_,r_141__45_,r_141__44_,r_141__43_,
  r_141__42_,r_141__41_,r_141__40_,r_141__39_,r_141__38_,r_141__37_,r_141__36_,
  r_141__35_,r_141__34_,r_141__33_,r_141__32_,r_141__31_,r_141__30_,r_141__29_,
  r_141__28_,r_141__27_,r_141__26_,r_141__25_,r_141__24_,r_141__23_,r_141__22_,
  r_141__21_,r_141__20_,r_141__19_,r_141__18_,r_141__17_,r_141__16_,r_141__15_,r_141__14_,
  r_141__13_,r_141__12_,r_141__11_,r_141__10_,r_141__9_,r_141__8_,r_141__7_,
  r_141__6_,r_141__5_,r_141__4_,r_141__3_,r_141__2_,r_141__1_,r_141__0_,r_142__63_,
  r_142__62_,r_142__61_,r_142__60_,r_142__59_,r_142__58_,r_142__57_,r_142__56_,
  r_142__55_,r_142__54_,r_142__53_,r_142__52_,r_142__51_,r_142__50_,r_142__49_,r_142__48_,
  r_142__47_,r_142__46_,r_142__45_,r_142__44_,r_142__43_,r_142__42_,r_142__41_,
  r_142__40_,r_142__39_,r_142__38_,r_142__37_,r_142__36_,r_142__35_,r_142__34_,
  r_142__33_,r_142__32_,r_142__31_,r_142__30_,r_142__29_,r_142__28_,r_142__27_,r_142__26_,
  r_142__25_,r_142__24_,r_142__23_,r_142__22_,r_142__21_,r_142__20_,r_142__19_,
  r_142__18_,r_142__17_,r_142__16_,r_142__15_,r_142__14_,r_142__13_,r_142__12_,
  r_142__11_,r_142__10_,r_142__9_,r_142__8_,r_142__7_,r_142__6_,r_142__5_,r_142__4_,
  r_142__3_,r_142__2_,r_142__1_,r_142__0_,r_143__63_,r_143__62_,r_143__61_,r_143__60_,
  r_143__59_,r_143__58_,r_143__57_,r_143__56_,r_143__55_,r_143__54_,r_143__53_,
  r_143__52_,r_143__51_,r_143__50_,r_143__49_,r_143__48_,r_143__47_,r_143__46_,
  r_143__45_,r_143__44_,r_143__43_,r_143__42_,r_143__41_,r_143__40_,r_143__39_,
  r_143__38_,r_143__37_,r_143__36_,r_143__35_,r_143__34_,r_143__33_,r_143__32_,r_143__31_,
  r_143__30_,r_143__29_,r_143__28_,r_143__27_,r_143__26_,r_143__25_,r_143__24_,
  r_143__23_,r_143__22_,r_143__21_,r_143__20_,r_143__19_,r_143__18_,r_143__17_,
  r_143__16_,r_143__15_,r_143__14_,r_143__13_,r_143__12_,r_143__11_,r_143__10_,r_143__9_,
  r_143__8_,r_143__7_,r_143__6_,r_143__5_,r_143__4_,r_143__3_,r_143__2_,r_143__1_,
  r_143__0_,r_144__63_,r_144__62_,r_144__61_,r_144__60_,r_144__59_,r_144__58_,
  r_144__57_,r_144__56_,r_144__55_,r_144__54_,r_144__53_,r_144__52_,r_144__51_,
  r_144__50_,r_144__49_,r_144__48_,r_144__47_,r_144__46_,r_144__45_,r_144__44_,
  r_144__43_,r_144__42_,r_144__41_,r_144__40_,r_144__39_,r_144__38_,r_144__37_,r_144__36_,
  r_144__35_,r_144__34_,r_144__33_,r_144__32_,r_144__31_,r_144__30_,r_144__29_,
  r_144__28_,r_144__27_,r_144__26_,r_144__25_,r_144__24_,r_144__23_,r_144__22_,
  r_144__21_,r_144__20_,r_144__19_,r_144__18_,r_144__17_,r_144__16_,r_144__15_,r_144__14_,
  r_144__13_,r_144__12_,r_144__11_,r_144__10_,r_144__9_,r_144__8_,r_144__7_,
  r_144__6_,r_144__5_,r_144__4_,r_144__3_,r_144__2_,r_144__1_,r_144__0_,r_145__63_,
  r_145__62_,r_145__61_,r_145__60_,r_145__59_,r_145__58_,r_145__57_,r_145__56_,
  r_145__55_,r_145__54_,r_145__53_,r_145__52_,r_145__51_,r_145__50_,r_145__49_,r_145__48_,
  r_145__47_,r_145__46_,r_145__45_,r_145__44_,r_145__43_,r_145__42_,r_145__41_,
  r_145__40_,r_145__39_,r_145__38_,r_145__37_,r_145__36_,r_145__35_,r_145__34_,
  r_145__33_,r_145__32_,r_145__31_,r_145__30_,r_145__29_,r_145__28_,r_145__27_,
  r_145__26_,r_145__25_,r_145__24_,r_145__23_,r_145__22_,r_145__21_,r_145__20_,r_145__19_,
  r_145__18_,r_145__17_,r_145__16_,r_145__15_,r_145__14_,r_145__13_,r_145__12_,
  r_145__11_,r_145__10_,r_145__9_,r_145__8_,r_145__7_,r_145__6_,r_145__5_,r_145__4_,
  r_145__3_,r_145__2_,r_145__1_,r_145__0_,r_146__63_,r_146__62_,r_146__61_,
  r_146__60_,r_146__59_,r_146__58_,r_146__57_,r_146__56_,r_146__55_,r_146__54_,r_146__53_,
  r_146__52_,r_146__51_,r_146__50_,r_146__49_,r_146__48_,r_146__47_,r_146__46_,
  r_146__45_,r_146__44_,r_146__43_,r_146__42_,r_146__41_,r_146__40_,r_146__39_,
  r_146__38_,r_146__37_,r_146__36_,r_146__35_,r_146__34_,r_146__33_,r_146__32_,
  r_146__31_,r_146__30_,r_146__29_,r_146__28_,r_146__27_,r_146__26_,r_146__25_,r_146__24_,
  r_146__23_,r_146__22_,r_146__21_,r_146__20_,r_146__19_,r_146__18_,r_146__17_,
  r_146__16_,r_146__15_,r_146__14_,r_146__13_,r_146__12_,r_146__11_,r_146__10_,
  r_146__9_,r_146__8_,r_146__7_,r_146__6_,r_146__5_,r_146__4_,r_146__3_,r_146__2_,
  r_146__1_,r_146__0_,r_147__63_,r_147__62_,r_147__61_,r_147__60_,r_147__59_,r_147__58_,
  r_147__57_,r_147__56_,r_147__55_,r_147__54_,r_147__53_,r_147__52_,r_147__51_,
  r_147__50_,r_147__49_,r_147__48_,r_147__47_,r_147__46_,r_147__45_,r_147__44_,
  r_147__43_,r_147__42_,r_147__41_,r_147__40_,r_147__39_,r_147__38_,r_147__37_,r_147__36_,
  r_147__35_,r_147__34_,r_147__33_,r_147__32_,r_147__31_,r_147__30_,r_147__29_,
  r_147__28_,r_147__27_,r_147__26_,r_147__25_,r_147__24_,r_147__23_,r_147__22_,
  r_147__21_,r_147__20_,r_147__19_,r_147__18_,r_147__17_,r_147__16_,r_147__15_,
  r_147__14_,r_147__13_,r_147__12_,r_147__11_,r_147__10_,r_147__9_,r_147__8_,r_147__7_,
  r_147__6_,r_147__5_,r_147__4_,r_147__3_,r_147__2_,r_147__1_,r_147__0_,r_148__63_,
  r_148__62_,r_148__61_,r_148__60_,r_148__59_,r_148__58_,r_148__57_,r_148__56_,
  r_148__55_,r_148__54_,r_148__53_,r_148__52_,r_148__51_,r_148__50_,r_148__49_,
  r_148__48_,r_148__47_,r_148__46_,r_148__45_,r_148__44_,r_148__43_,r_148__42_,r_148__41_,
  r_148__40_,r_148__39_,r_148__38_,r_148__37_,r_148__36_,r_148__35_,r_148__34_,
  r_148__33_,r_148__32_,r_148__31_,r_148__30_,r_148__29_,r_148__28_,r_148__27_,
  r_148__26_,r_148__25_,r_148__24_,r_148__23_,r_148__22_,r_148__21_,r_148__20_,
  r_148__19_,r_148__18_,r_148__17_,r_148__16_,r_148__15_,r_148__14_,r_148__13_,r_148__12_,
  r_148__11_,r_148__10_,r_148__9_,r_148__8_,r_148__7_,r_148__6_,r_148__5_,r_148__4_,
  r_148__3_,r_148__2_,r_148__1_,r_148__0_,r_149__63_,r_149__62_,r_149__61_,
  r_149__60_,r_149__59_,r_149__58_,r_149__57_,r_149__56_,r_149__55_,r_149__54_,
  r_149__53_,r_149__52_,r_149__51_,r_149__50_,r_149__49_,r_149__48_,r_149__47_,r_149__46_,
  r_149__45_,r_149__44_,r_149__43_,r_149__42_,r_149__41_,r_149__40_,r_149__39_,
  r_149__38_,r_149__37_,r_149__36_,r_149__35_,r_149__34_,r_149__33_,r_149__32_,
  r_149__31_,r_149__30_,r_149__29_,r_149__28_,r_149__27_,r_149__26_,r_149__25_,r_149__24_,
  r_149__23_,r_149__22_,r_149__21_,r_149__20_,r_149__19_,r_149__18_,r_149__17_,
  r_149__16_,r_149__15_,r_149__14_,r_149__13_,r_149__12_,r_149__11_,r_149__10_,
  r_149__9_,r_149__8_,r_149__7_,r_149__6_,r_149__5_,r_149__4_,r_149__3_,r_149__2_,
  r_149__1_,r_149__0_,r_150__63_,r_150__62_,r_150__61_,r_150__60_,r_150__59_,r_150__58_,
  r_150__57_,r_150__56_,r_150__55_,r_150__54_,r_150__53_,r_150__52_,r_150__51_,
  r_150__50_,r_150__49_,r_150__48_,r_150__47_,r_150__46_,r_150__45_,r_150__44_,
  r_150__43_,r_150__42_,r_150__41_,r_150__40_,r_150__39_,r_150__38_,r_150__37_,
  r_150__36_,r_150__35_,r_150__34_,r_150__33_,r_150__32_,r_150__31_,r_150__30_,r_150__29_,
  r_150__28_,r_150__27_,r_150__26_,r_150__25_,r_150__24_,r_150__23_,r_150__22_,
  r_150__21_,r_150__20_,r_150__19_,r_150__18_,r_150__17_,r_150__16_,r_150__15_,
  r_150__14_,r_150__13_,r_150__12_,r_150__11_,r_150__10_,r_150__9_,r_150__8_,r_150__7_,
  r_150__6_,r_150__5_,r_150__4_,r_150__3_,r_150__2_,r_150__1_,r_150__0_,r_151__63_,
  r_151__62_,r_151__61_,r_151__60_,r_151__59_,r_151__58_,r_151__57_,r_151__56_,
  r_151__55_,r_151__54_,r_151__53_,r_151__52_,r_151__51_,r_151__50_,r_151__49_,
  r_151__48_,r_151__47_,r_151__46_,r_151__45_,r_151__44_,r_151__43_,r_151__42_,
  r_151__41_,r_151__40_,r_151__39_,r_151__38_,r_151__37_,r_151__36_,r_151__35_,r_151__34_,
  r_151__33_,r_151__32_,r_151__31_,r_151__30_,r_151__29_,r_151__28_,r_151__27_,
  r_151__26_,r_151__25_,r_151__24_,r_151__23_,r_151__22_,r_151__21_,r_151__20_,
  r_151__19_,r_151__18_,r_151__17_,r_151__16_,r_151__15_,r_151__14_,r_151__13_,r_151__12_,
  r_151__11_,r_151__10_,r_151__9_,r_151__8_,r_151__7_,r_151__6_,r_151__5_,
  r_151__4_,r_151__3_,r_151__2_,r_151__1_,r_151__0_,r_152__63_,r_152__62_,r_152__61_,
  r_152__60_,r_152__59_,r_152__58_,r_152__57_,r_152__56_,r_152__55_,r_152__54_,
  r_152__53_,r_152__52_,r_152__51_,r_152__50_,r_152__49_,r_152__48_,r_152__47_,r_152__46_,
  r_152__45_,r_152__44_,r_152__43_,r_152__42_,r_152__41_,r_152__40_,r_152__39_,
  r_152__38_,r_152__37_,r_152__36_,r_152__35_,r_152__34_,r_152__33_,r_152__32_,
  r_152__31_,r_152__30_,r_152__29_,r_152__28_,r_152__27_,r_152__26_,r_152__25_,
  r_152__24_,r_152__23_,r_152__22_,r_152__21_,r_152__20_,r_152__19_,r_152__18_,r_152__17_,
  r_152__16_,r_152__15_,r_152__14_,r_152__13_,r_152__12_,r_152__11_,r_152__10_,
  r_152__9_,r_152__8_,r_152__7_,r_152__6_,r_152__5_,r_152__4_,r_152__3_,r_152__2_,
  r_152__1_,r_152__0_,r_153__63_,r_153__62_,r_153__61_,r_153__60_,r_153__59_,
  r_153__58_,r_153__57_,r_153__56_,r_153__55_,r_153__54_,r_153__53_,r_153__52_,r_153__51_,
  r_153__50_,r_153__49_,r_153__48_,r_153__47_,r_153__46_,r_153__45_,r_153__44_,
  r_153__43_,r_153__42_,r_153__41_,r_153__40_,r_153__39_,r_153__38_,r_153__37_,
  r_153__36_,r_153__35_,r_153__34_,r_153__33_,r_153__32_,r_153__31_,r_153__30_,
  r_153__29_,r_153__28_,r_153__27_,r_153__26_,r_153__25_,r_153__24_,r_153__23_,r_153__22_,
  r_153__21_,r_153__20_,r_153__19_,r_153__18_,r_153__17_,r_153__16_,r_153__15_,
  r_153__14_,r_153__13_,r_153__12_,r_153__11_,r_153__10_,r_153__9_,r_153__8_,r_153__7_,
  r_153__6_,r_153__5_,r_153__4_,r_153__3_,r_153__2_,r_153__1_,r_153__0_,
  r_154__63_,r_154__62_,r_154__61_,r_154__60_,r_154__59_,r_154__58_,r_154__57_,r_154__56_,
  r_154__55_,r_154__54_,r_154__53_,r_154__52_,r_154__51_,r_154__50_,r_154__49_,
  r_154__48_,r_154__47_,r_154__46_,r_154__45_,r_154__44_,r_154__43_,r_154__42_,
  r_154__41_,r_154__40_,r_154__39_,r_154__38_,r_154__37_,r_154__36_,r_154__35_,r_154__34_,
  r_154__33_,r_154__32_,r_154__31_,r_154__30_,r_154__29_,r_154__28_,r_154__27_,
  r_154__26_,r_154__25_,r_154__24_,r_154__23_,r_154__22_,r_154__21_,r_154__20_,
  r_154__19_,r_154__18_,r_154__17_,r_154__16_,r_154__15_,r_154__14_,r_154__13_,
  r_154__12_,r_154__11_,r_154__10_,r_154__9_,r_154__8_,r_154__7_,r_154__6_,r_154__5_,
  r_154__4_,r_154__3_,r_154__2_,r_154__1_,r_154__0_,r_155__63_,r_155__62_,r_155__61_,
  r_155__60_,r_155__59_,r_155__58_,r_155__57_,r_155__56_,r_155__55_,r_155__54_,
  r_155__53_,r_155__52_,r_155__51_,r_155__50_,r_155__49_,r_155__48_,r_155__47_,
  r_155__46_,r_155__45_,r_155__44_,r_155__43_,r_155__42_,r_155__41_,r_155__40_,r_155__39_,
  r_155__38_,r_155__37_,r_155__36_,r_155__35_,r_155__34_,r_155__33_,r_155__32_,
  r_155__31_,r_155__30_,r_155__29_,r_155__28_,r_155__27_,r_155__26_,r_155__25_,
  r_155__24_,r_155__23_,r_155__22_,r_155__21_,r_155__20_,r_155__19_,r_155__18_,
  r_155__17_,r_155__16_,r_155__15_,r_155__14_,r_155__13_,r_155__12_,r_155__11_,r_155__10_,
  r_155__9_,r_155__8_,r_155__7_,r_155__6_,r_155__5_,r_155__4_,r_155__3_,r_155__2_,
  r_155__1_,r_155__0_,r_156__63_,r_156__62_,r_156__61_,r_156__60_,r_156__59_,
  r_156__58_,r_156__57_,r_156__56_,r_156__55_,r_156__54_,r_156__53_,r_156__52_,
  r_156__51_,r_156__50_,r_156__49_,r_156__48_,r_156__47_,r_156__46_,r_156__45_,r_156__44_,
  r_156__43_,r_156__42_,r_156__41_,r_156__40_,r_156__39_,r_156__38_,r_156__37_,
  r_156__36_,r_156__35_,r_156__34_,r_156__33_,r_156__32_,r_156__31_,r_156__30_,
  r_156__29_,r_156__28_,r_156__27_,r_156__26_,r_156__25_,r_156__24_,r_156__23_,r_156__22_,
  r_156__21_,r_156__20_,r_156__19_,r_156__18_,r_156__17_,r_156__16_,r_156__15_,
  r_156__14_,r_156__13_,r_156__12_,r_156__11_,r_156__10_,r_156__9_,r_156__8_,
  r_156__7_,r_156__6_,r_156__5_,r_156__4_,r_156__3_,r_156__2_,r_156__1_,r_156__0_,
  r_157__63_,r_157__62_,r_157__61_,r_157__60_,r_157__59_,r_157__58_,r_157__57_,r_157__56_,
  r_157__55_,r_157__54_,r_157__53_,r_157__52_,r_157__51_,r_157__50_,r_157__49_,
  r_157__48_,r_157__47_,r_157__46_,r_157__45_,r_157__44_,r_157__43_,r_157__42_,
  r_157__41_,r_157__40_,r_157__39_,r_157__38_,r_157__37_,r_157__36_,r_157__35_,
  r_157__34_,r_157__33_,r_157__32_,r_157__31_,r_157__30_,r_157__29_,r_157__28_,r_157__27_,
  r_157__26_,r_157__25_,r_157__24_,r_157__23_,r_157__22_,r_157__21_,r_157__20_,
  r_157__19_,r_157__18_,r_157__17_,r_157__16_,r_157__15_,r_157__14_,r_157__13_,
  r_157__12_,r_157__11_,r_157__10_,r_157__9_,r_157__8_,r_157__7_,r_157__6_,r_157__5_,
  r_157__4_,r_157__3_,r_157__2_,r_157__1_,r_157__0_,r_158__63_,r_158__62_,r_158__61_,
  r_158__60_,r_158__59_,r_158__58_,r_158__57_,r_158__56_,r_158__55_,r_158__54_,
  r_158__53_,r_158__52_,r_158__51_,r_158__50_,r_158__49_,r_158__48_,r_158__47_,
  r_158__46_,r_158__45_,r_158__44_,r_158__43_,r_158__42_,r_158__41_,r_158__40_,
  r_158__39_,r_158__38_,r_158__37_,r_158__36_,r_158__35_,r_158__34_,r_158__33_,r_158__32_,
  r_158__31_,r_158__30_,r_158__29_,r_158__28_,r_158__27_,r_158__26_,r_158__25_,
  r_158__24_,r_158__23_,r_158__22_,r_158__21_,r_158__20_,r_158__19_,r_158__18_,
  r_158__17_,r_158__16_,r_158__15_,r_158__14_,r_158__13_,r_158__12_,r_158__11_,r_158__10_,
  r_158__9_,r_158__8_,r_158__7_,r_158__6_,r_158__5_,r_158__4_,r_158__3_,r_158__2_,
  r_158__1_,r_158__0_,r_159__63_,r_159__62_,r_159__61_,r_159__60_,r_159__59_,
  r_159__58_,r_159__57_,r_159__56_,r_159__55_,r_159__54_,r_159__53_,r_159__52_,
  r_159__51_,r_159__50_,r_159__49_,r_159__48_,r_159__47_,r_159__46_,r_159__45_,r_159__44_,
  r_159__43_,r_159__42_,r_159__41_,r_159__40_,r_159__39_,r_159__38_,r_159__37_,
  r_159__36_,r_159__35_,r_159__34_,r_159__33_,r_159__32_,r_159__31_,r_159__30_,
  r_159__29_,r_159__28_,r_159__27_,r_159__26_,r_159__25_,r_159__24_,r_159__23_,
  r_159__22_,r_159__21_,r_159__20_,r_159__19_,r_159__18_,r_159__17_,r_159__16_,r_159__15_,
  r_159__14_,r_159__13_,r_159__12_,r_159__11_,r_159__10_,r_159__9_,r_159__8_,
  r_159__7_,r_159__6_,r_159__5_,r_159__4_,r_159__3_,r_159__2_,r_159__1_,r_159__0_,
  r_160__63_,r_160__62_,r_160__61_,r_160__60_,r_160__59_,r_160__58_,r_160__57_,
  r_160__56_,r_160__55_,r_160__54_,r_160__53_,r_160__52_,r_160__51_,r_160__50_,r_160__49_,
  r_160__48_,r_160__47_,r_160__46_,r_160__45_,r_160__44_,r_160__43_,r_160__42_,
  r_160__41_,r_160__40_,r_160__39_,r_160__38_,r_160__37_,r_160__36_,r_160__35_,
  r_160__34_,r_160__33_,r_160__32_,r_160__31_,r_160__30_,r_160__29_,r_160__28_,
  r_160__27_,r_160__26_,r_160__25_,r_160__24_,r_160__23_,r_160__22_,r_160__21_,r_160__20_,
  r_160__19_,r_160__18_,r_160__17_,r_160__16_,r_160__15_,r_160__14_,r_160__13_,
  r_160__12_,r_160__11_,r_160__10_,r_160__9_,r_160__8_,r_160__7_,r_160__6_,r_160__5_,
  r_160__4_,r_160__3_,r_160__2_,r_160__1_,r_160__0_,r_161__63_,r_161__62_,
  r_161__61_,r_161__60_,r_161__59_,r_161__58_,r_161__57_,r_161__56_,r_161__55_,r_161__54_,
  r_161__53_,r_161__52_,r_161__51_,r_161__50_,r_161__49_,r_161__48_,r_161__47_,
  r_161__46_,r_161__45_,r_161__44_,r_161__43_,r_161__42_,r_161__41_,r_161__40_,
  r_161__39_,r_161__38_,r_161__37_,r_161__36_,r_161__35_,r_161__34_,r_161__33_,r_161__32_,
  r_161__31_,r_161__30_,r_161__29_,r_161__28_,r_161__27_,r_161__26_,r_161__25_,
  r_161__24_,r_161__23_,r_161__22_,r_161__21_,r_161__20_,r_161__19_,r_161__18_,
  r_161__17_,r_161__16_,r_161__15_,r_161__14_,r_161__13_,r_161__12_,r_161__11_,
  r_161__10_,r_161__9_,r_161__8_,r_161__7_,r_161__6_,r_161__5_,r_161__4_,r_161__3_,
  r_161__2_,r_161__1_,r_161__0_,r_162__63_,r_162__62_,r_162__61_,r_162__60_,r_162__59_,
  r_162__58_,r_162__57_,r_162__56_,r_162__55_,r_162__54_,r_162__53_,r_162__52_,
  r_162__51_,r_162__50_,r_162__49_,r_162__48_,r_162__47_,r_162__46_,r_162__45_,
  r_162__44_,r_162__43_,r_162__42_,r_162__41_,r_162__40_,r_162__39_,r_162__38_,r_162__37_,
  r_162__36_,r_162__35_,r_162__34_,r_162__33_,r_162__32_,r_162__31_,r_162__30_,
  r_162__29_,r_162__28_,r_162__27_,r_162__26_,r_162__25_,r_162__24_,r_162__23_,
  r_162__22_,r_162__21_,r_162__20_,r_162__19_,r_162__18_,r_162__17_,r_162__16_,
  r_162__15_,r_162__14_,r_162__13_,r_162__12_,r_162__11_,r_162__10_,r_162__9_,r_162__8_,
  r_162__7_,r_162__6_,r_162__5_,r_162__4_,r_162__3_,r_162__2_,r_162__1_,r_162__0_,
  r_163__63_,r_163__62_,r_163__61_,r_163__60_,r_163__59_,r_163__58_,r_163__57_,
  r_163__56_,r_163__55_,r_163__54_,r_163__53_,r_163__52_,r_163__51_,r_163__50_,
  r_163__49_,r_163__48_,r_163__47_,r_163__46_,r_163__45_,r_163__44_,r_163__43_,r_163__42_,
  r_163__41_,r_163__40_,r_163__39_,r_163__38_,r_163__37_,r_163__36_,r_163__35_,
  r_163__34_,r_163__33_,r_163__32_,r_163__31_,r_163__30_,r_163__29_,r_163__28_,
  r_163__27_,r_163__26_,r_163__25_,r_163__24_,r_163__23_,r_163__22_,r_163__21_,r_163__20_,
  r_163__19_,r_163__18_,r_163__17_,r_163__16_,r_163__15_,r_163__14_,r_163__13_,
  r_163__12_,r_163__11_,r_163__10_,r_163__9_,r_163__8_,r_163__7_,r_163__6_,r_163__5_,
  r_163__4_,r_163__3_,r_163__2_,r_163__1_,r_163__0_,r_164__63_,r_164__62_,
  r_164__61_,r_164__60_,r_164__59_,r_164__58_,r_164__57_,r_164__56_,r_164__55_,r_164__54_,
  r_164__53_,r_164__52_,r_164__51_,r_164__50_,r_164__49_,r_164__48_,r_164__47_,
  r_164__46_,r_164__45_,r_164__44_,r_164__43_,r_164__42_,r_164__41_,r_164__40_,
  r_164__39_,r_164__38_,r_164__37_,r_164__36_,r_164__35_,r_164__34_,r_164__33_,
  r_164__32_,r_164__31_,r_164__30_,r_164__29_,r_164__28_,r_164__27_,r_164__26_,r_164__25_,
  r_164__24_,r_164__23_,r_164__22_,r_164__21_,r_164__20_,r_164__19_,r_164__18_,
  r_164__17_,r_164__16_,r_164__15_,r_164__14_,r_164__13_,r_164__12_,r_164__11_,
  r_164__10_,r_164__9_,r_164__8_,r_164__7_,r_164__6_,r_164__5_,r_164__4_,r_164__3_,
  r_164__2_,r_164__1_,r_164__0_,r_165__63_,r_165__62_,r_165__61_,r_165__60_,r_165__59_,
  r_165__58_,r_165__57_,r_165__56_,r_165__55_,r_165__54_,r_165__53_,r_165__52_,
  r_165__51_,r_165__50_,r_165__49_,r_165__48_,r_165__47_,r_165__46_,r_165__45_,
  r_165__44_,r_165__43_,r_165__42_,r_165__41_,r_165__40_,r_165__39_,r_165__38_,
  r_165__37_,r_165__36_,r_165__35_,r_165__34_,r_165__33_,r_165__32_,r_165__31_,r_165__30_,
  r_165__29_,r_165__28_,r_165__27_,r_165__26_,r_165__25_,r_165__24_,r_165__23_,
  r_165__22_,r_165__21_,r_165__20_,r_165__19_,r_165__18_,r_165__17_,r_165__16_,
  r_165__15_,r_165__14_,r_165__13_,r_165__12_,r_165__11_,r_165__10_,r_165__9_,r_165__8_,
  r_165__7_,r_165__6_,r_165__5_,r_165__4_,r_165__3_,r_165__2_,r_165__1_,r_165__0_,
  r_166__63_,r_166__62_,r_166__61_,r_166__60_,r_166__59_,r_166__58_,r_166__57_,
  r_166__56_,r_166__55_,r_166__54_,r_166__53_,r_166__52_,r_166__51_,r_166__50_,
  r_166__49_,r_166__48_,r_166__47_,r_166__46_,r_166__45_,r_166__44_,r_166__43_,r_166__42_,
  r_166__41_,r_166__40_,r_166__39_,r_166__38_,r_166__37_,r_166__36_,r_166__35_,
  r_166__34_,r_166__33_,r_166__32_,r_166__31_,r_166__30_,r_166__29_,r_166__28_,
  r_166__27_,r_166__26_,r_166__25_,r_166__24_,r_166__23_,r_166__22_,r_166__21_,
  r_166__20_,r_166__19_,r_166__18_,r_166__17_,r_166__16_,r_166__15_,r_166__14_,r_166__13_,
  r_166__12_,r_166__11_,r_166__10_,r_166__9_,r_166__8_,r_166__7_,r_166__6_,
  r_166__5_,r_166__4_,r_166__3_,r_166__2_,r_166__1_,r_166__0_,r_167__63_,r_167__62_,
  r_167__61_,r_167__60_,r_167__59_,r_167__58_,r_167__57_,r_167__56_,r_167__55_,
  r_167__54_,r_167__53_,r_167__52_,r_167__51_,r_167__50_,r_167__49_,r_167__48_,r_167__47_,
  r_167__46_,r_167__45_,r_167__44_,r_167__43_,r_167__42_,r_167__41_,r_167__40_,
  r_167__39_,r_167__38_,r_167__37_,r_167__36_,r_167__35_,r_167__34_,r_167__33_,
  r_167__32_,r_167__31_,r_167__30_,r_167__29_,r_167__28_,r_167__27_,r_167__26_,
  r_167__25_,r_167__24_,r_167__23_,r_167__22_,r_167__21_,r_167__20_,r_167__19_,r_167__18_,
  r_167__17_,r_167__16_,r_167__15_,r_167__14_,r_167__13_,r_167__12_,r_167__11_,
  r_167__10_,r_167__9_,r_167__8_,r_167__7_,r_167__6_,r_167__5_,r_167__4_,r_167__3_,
  r_167__2_,r_167__1_,r_167__0_,r_168__63_,r_168__62_,r_168__61_,r_168__60_,
  r_168__59_,r_168__58_,r_168__57_,r_168__56_,r_168__55_,r_168__54_,r_168__53_,r_168__52_,
  r_168__51_,r_168__50_,r_168__49_,r_168__48_,r_168__47_,r_168__46_,r_168__45_,
  r_168__44_,r_168__43_,r_168__42_,r_168__41_,r_168__40_,r_168__39_,r_168__38_,
  r_168__37_,r_168__36_,r_168__35_,r_168__34_,r_168__33_,r_168__32_,r_168__31_,r_168__30_,
  r_168__29_,r_168__28_,r_168__27_,r_168__26_,r_168__25_,r_168__24_,r_168__23_,
  r_168__22_,r_168__21_,r_168__20_,r_168__19_,r_168__18_,r_168__17_,r_168__16_,
  r_168__15_,r_168__14_,r_168__13_,r_168__12_,r_168__11_,r_168__10_,r_168__9_,r_168__8_,
  r_168__7_,r_168__6_,r_168__5_,r_168__4_,r_168__3_,r_168__2_,r_168__1_,r_168__0_,
  r_169__63_,r_169__62_,r_169__61_,r_169__60_,r_169__59_,r_169__58_,r_169__57_,
  r_169__56_,r_169__55_,r_169__54_,r_169__53_,r_169__52_,r_169__51_,r_169__50_,
  r_169__49_,r_169__48_,r_169__47_,r_169__46_,r_169__45_,r_169__44_,r_169__43_,
  r_169__42_,r_169__41_,r_169__40_,r_169__39_,r_169__38_,r_169__37_,r_169__36_,r_169__35_,
  r_169__34_,r_169__33_,r_169__32_,r_169__31_,r_169__30_,r_169__29_,r_169__28_,
  r_169__27_,r_169__26_,r_169__25_,r_169__24_,r_169__23_,r_169__22_,r_169__21_,
  r_169__20_,r_169__19_,r_169__18_,r_169__17_,r_169__16_,r_169__15_,r_169__14_,
  r_169__13_,r_169__12_,r_169__11_,r_169__10_,r_169__9_,r_169__8_,r_169__7_,r_169__6_,
  r_169__5_,r_169__4_,r_169__3_,r_169__2_,r_169__1_,r_169__0_,r_170__63_,r_170__62_,
  r_170__61_,r_170__60_,r_170__59_,r_170__58_,r_170__57_,r_170__56_,r_170__55_,
  r_170__54_,r_170__53_,r_170__52_,r_170__51_,r_170__50_,r_170__49_,r_170__48_,
  r_170__47_,r_170__46_,r_170__45_,r_170__44_,r_170__43_,r_170__42_,r_170__41_,r_170__40_,
  r_170__39_,r_170__38_,r_170__37_,r_170__36_,r_170__35_,r_170__34_,r_170__33_,
  r_170__32_,r_170__31_,r_170__30_,r_170__29_,r_170__28_,r_170__27_,r_170__26_,
  r_170__25_,r_170__24_,r_170__23_,r_170__22_,r_170__21_,r_170__20_,r_170__19_,r_170__18_,
  r_170__17_,r_170__16_,r_170__15_,r_170__14_,r_170__13_,r_170__12_,r_170__11_,
  r_170__10_,r_170__9_,r_170__8_,r_170__7_,r_170__6_,r_170__5_,r_170__4_,r_170__3_,
  r_170__2_,r_170__1_,r_170__0_,r_171__63_,r_171__62_,r_171__61_,r_171__60_,
  r_171__59_,r_171__58_,r_171__57_,r_171__56_,r_171__55_,r_171__54_,r_171__53_,r_171__52_,
  r_171__51_,r_171__50_,r_171__49_,r_171__48_,r_171__47_,r_171__46_,r_171__45_,
  r_171__44_,r_171__43_,r_171__42_,r_171__41_,r_171__40_,r_171__39_,r_171__38_,
  r_171__37_,r_171__36_,r_171__35_,r_171__34_,r_171__33_,r_171__32_,r_171__31_,
  r_171__30_,r_171__29_,r_171__28_,r_171__27_,r_171__26_,r_171__25_,r_171__24_,r_171__23_,
  r_171__22_,r_171__21_,r_171__20_,r_171__19_,r_171__18_,r_171__17_,r_171__16_,
  r_171__15_,r_171__14_,r_171__13_,r_171__12_,r_171__11_,r_171__10_,r_171__9_,
  r_171__8_,r_171__7_,r_171__6_,r_171__5_,r_171__4_,r_171__3_,r_171__2_,r_171__1_,
  r_171__0_,r_172__63_,r_172__62_,r_172__61_,r_172__60_,r_172__59_,r_172__58_,r_172__57_,
  r_172__56_,r_172__55_,r_172__54_,r_172__53_,r_172__52_,r_172__51_,r_172__50_,
  r_172__49_,r_172__48_,r_172__47_,r_172__46_,r_172__45_,r_172__44_,r_172__43_,
  r_172__42_,r_172__41_,r_172__40_,r_172__39_,r_172__38_,r_172__37_,r_172__36_,
  r_172__35_,r_172__34_,r_172__33_,r_172__32_,r_172__31_,r_172__30_,r_172__29_,r_172__28_,
  r_172__27_,r_172__26_,r_172__25_,r_172__24_,r_172__23_,r_172__22_,r_172__21_,
  r_172__20_,r_172__19_,r_172__18_,r_172__17_,r_172__16_,r_172__15_,r_172__14_,
  r_172__13_,r_172__12_,r_172__11_,r_172__10_,r_172__9_,r_172__8_,r_172__7_,r_172__6_,
  r_172__5_,r_172__4_,r_172__3_,r_172__2_,r_172__1_,r_172__0_,r_173__63_,r_173__62_,
  r_173__61_,r_173__60_,r_173__59_,r_173__58_,r_173__57_,r_173__56_,r_173__55_,
  r_173__54_,r_173__53_,r_173__52_,r_173__51_,r_173__50_,r_173__49_,r_173__48_,
  r_173__47_,r_173__46_,r_173__45_,r_173__44_,r_173__43_,r_173__42_,r_173__41_,r_173__40_,
  r_173__39_,r_173__38_,r_173__37_,r_173__36_,r_173__35_,r_173__34_,r_173__33_,
  r_173__32_,r_173__31_,r_173__30_,r_173__29_,r_173__28_,r_173__27_,r_173__26_,
  r_173__25_,r_173__24_,r_173__23_,r_173__22_,r_173__21_,r_173__20_,r_173__19_,
  r_173__18_,r_173__17_,r_173__16_,r_173__15_,r_173__14_,r_173__13_,r_173__12_,r_173__11_,
  r_173__10_,r_173__9_,r_173__8_,r_173__7_,r_173__6_,r_173__5_,r_173__4_,r_173__3_,
  r_173__2_,r_173__1_,r_173__0_,r_174__63_,r_174__62_,r_174__61_,r_174__60_,
  r_174__59_,r_174__58_,r_174__57_,r_174__56_,r_174__55_,r_174__54_,r_174__53_,
  r_174__52_,r_174__51_,r_174__50_,r_174__49_,r_174__48_,r_174__47_,r_174__46_,r_174__45_,
  r_174__44_,r_174__43_,r_174__42_,r_174__41_,r_174__40_,r_174__39_,r_174__38_,
  r_174__37_,r_174__36_,r_174__35_,r_174__34_,r_174__33_,r_174__32_,r_174__31_,
  r_174__30_,r_174__29_,r_174__28_,r_174__27_,r_174__26_,r_174__25_,r_174__24_,
  r_174__23_,r_174__22_,r_174__21_,r_174__20_,r_174__19_,r_174__18_,r_174__17_,r_174__16_,
  r_174__15_,r_174__14_,r_174__13_,r_174__12_,r_174__11_,r_174__10_,r_174__9_,
  r_174__8_,r_174__7_,r_174__6_,r_174__5_,r_174__4_,r_174__3_,r_174__2_,r_174__1_,
  r_174__0_,r_175__63_,r_175__62_,r_175__61_,r_175__60_,r_175__59_,r_175__58_,
  r_175__57_,r_175__56_,r_175__55_,r_175__54_,r_175__53_,r_175__52_,r_175__51_,r_175__50_,
  r_175__49_,r_175__48_,r_175__47_,r_175__46_,r_175__45_,r_175__44_,r_175__43_,
  r_175__42_,r_175__41_,r_175__40_,r_175__39_,r_175__38_,r_175__37_,r_175__36_,
  r_175__35_,r_175__34_,r_175__33_,r_175__32_,r_175__31_,r_175__30_,r_175__29_,r_175__28_,
  r_175__27_,r_175__26_,r_175__25_,r_175__24_,r_175__23_,r_175__22_,r_175__21_,
  r_175__20_,r_175__19_,r_175__18_,r_175__17_,r_175__16_,r_175__15_,r_175__14_,
  r_175__13_,r_175__12_,r_175__11_,r_175__10_,r_175__9_,r_175__8_,r_175__7_,r_175__6_,
  r_175__5_,r_175__4_,r_175__3_,r_175__2_,r_175__1_,r_175__0_,r_176__63_,r_176__62_,
  r_176__61_,r_176__60_,r_176__59_,r_176__58_,r_176__57_,r_176__56_,r_176__55_,
  r_176__54_,r_176__53_,r_176__52_,r_176__51_,r_176__50_,r_176__49_,r_176__48_,
  r_176__47_,r_176__46_,r_176__45_,r_176__44_,r_176__43_,r_176__42_,r_176__41_,
  r_176__40_,r_176__39_,r_176__38_,r_176__37_,r_176__36_,r_176__35_,r_176__34_,r_176__33_,
  r_176__32_,r_176__31_,r_176__30_,r_176__29_,r_176__28_,r_176__27_,r_176__26_,
  r_176__25_,r_176__24_,r_176__23_,r_176__22_,r_176__21_,r_176__20_,r_176__19_,
  r_176__18_,r_176__17_,r_176__16_,r_176__15_,r_176__14_,r_176__13_,r_176__12_,
  r_176__11_,r_176__10_,r_176__9_,r_176__8_,r_176__7_,r_176__6_,r_176__5_,r_176__4_,
  r_176__3_,r_176__2_,r_176__1_,r_176__0_,r_177__63_,r_177__62_,r_177__61_,r_177__60_,
  r_177__59_,r_177__58_,r_177__57_,r_177__56_,r_177__55_,r_177__54_,r_177__53_,
  r_177__52_,r_177__51_,r_177__50_,r_177__49_,r_177__48_,r_177__47_,r_177__46_,
  r_177__45_,r_177__44_,r_177__43_,r_177__42_,r_177__41_,r_177__40_,r_177__39_,r_177__38_,
  r_177__37_,r_177__36_,r_177__35_,r_177__34_,r_177__33_,r_177__32_,r_177__31_,
  r_177__30_,r_177__29_,r_177__28_,r_177__27_,r_177__26_,r_177__25_,r_177__24_,
  r_177__23_,r_177__22_,r_177__21_,r_177__20_,r_177__19_,r_177__18_,r_177__17_,r_177__16_,
  r_177__15_,r_177__14_,r_177__13_,r_177__12_,r_177__11_,r_177__10_,r_177__9_,
  r_177__8_,r_177__7_,r_177__6_,r_177__5_,r_177__4_,r_177__3_,r_177__2_,r_177__1_,
  r_177__0_,r_178__63_,r_178__62_,r_178__61_,r_178__60_,r_178__59_,r_178__58_,
  r_178__57_,r_178__56_,r_178__55_,r_178__54_,r_178__53_,r_178__52_,r_178__51_,r_178__50_,
  r_178__49_,r_178__48_,r_178__47_,r_178__46_,r_178__45_,r_178__44_,r_178__43_,
  r_178__42_,r_178__41_,r_178__40_,r_178__39_,r_178__38_,r_178__37_,r_178__36_,
  r_178__35_,r_178__34_,r_178__33_,r_178__32_,r_178__31_,r_178__30_,r_178__29_,
  r_178__28_,r_178__27_,r_178__26_,r_178__25_,r_178__24_,r_178__23_,r_178__22_,r_178__21_,
  r_178__20_,r_178__19_,r_178__18_,r_178__17_,r_178__16_,r_178__15_,r_178__14_,
  r_178__13_,r_178__12_,r_178__11_,r_178__10_,r_178__9_,r_178__8_,r_178__7_,r_178__6_,
  r_178__5_,r_178__4_,r_178__3_,r_178__2_,r_178__1_,r_178__0_,r_179__63_,
  r_179__62_,r_179__61_,r_179__60_,r_179__59_,r_179__58_,r_179__57_,r_179__56_,r_179__55_,
  r_179__54_,r_179__53_,r_179__52_,r_179__51_,r_179__50_,r_179__49_,r_179__48_,
  r_179__47_,r_179__46_,r_179__45_,r_179__44_,r_179__43_,r_179__42_,r_179__41_,
  r_179__40_,r_179__39_,r_179__38_,r_179__37_,r_179__36_,r_179__35_,r_179__34_,
  r_179__33_,r_179__32_,r_179__31_,r_179__30_,r_179__29_,r_179__28_,r_179__27_,r_179__26_,
  r_179__25_,r_179__24_,r_179__23_,r_179__22_,r_179__21_,r_179__20_,r_179__19_,
  r_179__18_,r_179__17_,r_179__16_,r_179__15_,r_179__14_,r_179__13_,r_179__12_,
  r_179__11_,r_179__10_,r_179__9_,r_179__8_,r_179__7_,r_179__6_,r_179__5_,r_179__4_,
  r_179__3_,r_179__2_,r_179__1_,r_179__0_,r_180__63_,r_180__62_,r_180__61_,r_180__60_,
  r_180__59_,r_180__58_,r_180__57_,r_180__56_,r_180__55_,r_180__54_,r_180__53_,
  r_180__52_,r_180__51_,r_180__50_,r_180__49_,r_180__48_,r_180__47_,r_180__46_,
  r_180__45_,r_180__44_,r_180__43_,r_180__42_,r_180__41_,r_180__40_,r_180__39_,r_180__38_,
  r_180__37_,r_180__36_,r_180__35_,r_180__34_,r_180__33_,r_180__32_,r_180__31_,
  r_180__30_,r_180__29_,r_180__28_,r_180__27_,r_180__26_,r_180__25_,r_180__24_,
  r_180__23_,r_180__22_,r_180__21_,r_180__20_,r_180__19_,r_180__18_,r_180__17_,
  r_180__16_,r_180__15_,r_180__14_,r_180__13_,r_180__12_,r_180__11_,r_180__10_,r_180__9_,
  r_180__8_,r_180__7_,r_180__6_,r_180__5_,r_180__4_,r_180__3_,r_180__2_,r_180__1_,
  r_180__0_,r_181__63_,r_181__62_,r_181__61_,r_181__60_,r_181__59_,r_181__58_,
  r_181__57_,r_181__56_,r_181__55_,r_181__54_,r_181__53_,r_181__52_,r_181__51_,
  r_181__50_,r_181__49_,r_181__48_,r_181__47_,r_181__46_,r_181__45_,r_181__44_,r_181__43_,
  r_181__42_,r_181__41_,r_181__40_,r_181__39_,r_181__38_,r_181__37_,r_181__36_,
  r_181__35_,r_181__34_,r_181__33_,r_181__32_,r_181__31_,r_181__30_,r_181__29_,
  r_181__28_,r_181__27_,r_181__26_,r_181__25_,r_181__24_,r_181__23_,r_181__22_,
  r_181__21_,r_181__20_,r_181__19_,r_181__18_,r_181__17_,r_181__16_,r_181__15_,r_181__14_,
  r_181__13_,r_181__12_,r_181__11_,r_181__10_,r_181__9_,r_181__8_,r_181__7_,
  r_181__6_,r_181__5_,r_181__4_,r_181__3_,r_181__2_,r_181__1_,r_181__0_,r_182__63_,
  r_182__62_,r_182__61_,r_182__60_,r_182__59_,r_182__58_,r_182__57_,r_182__56_,
  r_182__55_,r_182__54_,r_182__53_,r_182__52_,r_182__51_,r_182__50_,r_182__49_,r_182__48_,
  r_182__47_,r_182__46_,r_182__45_,r_182__44_,r_182__43_,r_182__42_,r_182__41_,
  r_182__40_,r_182__39_,r_182__38_,r_182__37_,r_182__36_,r_182__35_,r_182__34_,
  r_182__33_,r_182__32_,r_182__31_,r_182__30_,r_182__29_,r_182__28_,r_182__27_,r_182__26_,
  r_182__25_,r_182__24_,r_182__23_,r_182__22_,r_182__21_,r_182__20_,r_182__19_,
  r_182__18_,r_182__17_,r_182__16_,r_182__15_,r_182__14_,r_182__13_,r_182__12_,
  r_182__11_,r_182__10_,r_182__9_,r_182__8_,r_182__7_,r_182__6_,r_182__5_,r_182__4_,
  r_182__3_,r_182__2_,r_182__1_,r_182__0_,r_183__63_,r_183__62_,r_183__61_,r_183__60_,
  r_183__59_,r_183__58_,r_183__57_,r_183__56_,r_183__55_,r_183__54_,r_183__53_,
  r_183__52_,r_183__51_,r_183__50_,r_183__49_,r_183__48_,r_183__47_,r_183__46_,
  r_183__45_,r_183__44_,r_183__43_,r_183__42_,r_183__41_,r_183__40_,r_183__39_,
  r_183__38_,r_183__37_,r_183__36_,r_183__35_,r_183__34_,r_183__33_,r_183__32_,r_183__31_,
  r_183__30_,r_183__29_,r_183__28_,r_183__27_,r_183__26_,r_183__25_,r_183__24_,
  r_183__23_,r_183__22_,r_183__21_,r_183__20_,r_183__19_,r_183__18_,r_183__17_,
  r_183__16_,r_183__15_,r_183__14_,r_183__13_,r_183__12_,r_183__11_,r_183__10_,r_183__9_,
  r_183__8_,r_183__7_,r_183__6_,r_183__5_,r_183__4_,r_183__3_,r_183__2_,r_183__1_,
  r_183__0_,r_184__63_,r_184__62_,r_184__61_,r_184__60_,r_184__59_,r_184__58_,
  r_184__57_,r_184__56_,r_184__55_,r_184__54_,r_184__53_,r_184__52_,r_184__51_,
  r_184__50_,r_184__49_,r_184__48_,r_184__47_,r_184__46_,r_184__45_,r_184__44_,
  r_184__43_,r_184__42_,r_184__41_,r_184__40_,r_184__39_,r_184__38_,r_184__37_,r_184__36_,
  r_184__35_,r_184__34_,r_184__33_,r_184__32_,r_184__31_,r_184__30_,r_184__29_,
  r_184__28_,r_184__27_,r_184__26_,r_184__25_,r_184__24_,r_184__23_,r_184__22_,
  r_184__21_,r_184__20_,r_184__19_,r_184__18_,r_184__17_,r_184__16_,r_184__15_,r_184__14_,
  r_184__13_,r_184__12_,r_184__11_,r_184__10_,r_184__9_,r_184__8_,r_184__7_,
  r_184__6_,r_184__5_,r_184__4_,r_184__3_,r_184__2_,r_184__1_,r_184__0_,r_185__63_,
  r_185__62_,r_185__61_,r_185__60_,r_185__59_,r_185__58_,r_185__57_,r_185__56_,
  r_185__55_,r_185__54_,r_185__53_,r_185__52_,r_185__51_,r_185__50_,r_185__49_,r_185__48_,
  r_185__47_,r_185__46_,r_185__45_,r_185__44_,r_185__43_,r_185__42_,r_185__41_,
  r_185__40_,r_185__39_,r_185__38_,r_185__37_,r_185__36_,r_185__35_,r_185__34_,
  r_185__33_,r_185__32_,r_185__31_,r_185__30_,r_185__29_,r_185__28_,r_185__27_,
  r_185__26_,r_185__25_,r_185__24_,r_185__23_,r_185__22_,r_185__21_,r_185__20_,r_185__19_,
  r_185__18_,r_185__17_,r_185__16_,r_185__15_,r_185__14_,r_185__13_,r_185__12_,
  r_185__11_,r_185__10_,r_185__9_,r_185__8_,r_185__7_,r_185__6_,r_185__5_,r_185__4_,
  r_185__3_,r_185__2_,r_185__1_,r_185__0_,r_186__63_,r_186__62_,r_186__61_,
  r_186__60_,r_186__59_,r_186__58_,r_186__57_,r_186__56_,r_186__55_,r_186__54_,r_186__53_,
  r_186__52_,r_186__51_,r_186__50_,r_186__49_,r_186__48_,r_186__47_,r_186__46_,
  r_186__45_,r_186__44_,r_186__43_,r_186__42_,r_186__41_,r_186__40_,r_186__39_,
  r_186__38_,r_186__37_,r_186__36_,r_186__35_,r_186__34_,r_186__33_,r_186__32_,
  r_186__31_,r_186__30_,r_186__29_,r_186__28_,r_186__27_,r_186__26_,r_186__25_,r_186__24_,
  r_186__23_,r_186__22_,r_186__21_,r_186__20_,r_186__19_,r_186__18_,r_186__17_,
  r_186__16_,r_186__15_,r_186__14_,r_186__13_,r_186__12_,r_186__11_,r_186__10_,
  r_186__9_,r_186__8_,r_186__7_,r_186__6_,r_186__5_,r_186__4_,r_186__3_,r_186__2_,
  r_186__1_,r_186__0_,r_187__63_,r_187__62_,r_187__61_,r_187__60_,r_187__59_,r_187__58_,
  r_187__57_,r_187__56_,r_187__55_,r_187__54_,r_187__53_,r_187__52_,r_187__51_,
  r_187__50_,r_187__49_,r_187__48_,r_187__47_,r_187__46_,r_187__45_,r_187__44_,
  r_187__43_,r_187__42_,r_187__41_,r_187__40_,r_187__39_,r_187__38_,r_187__37_,r_187__36_,
  r_187__35_,r_187__34_,r_187__33_,r_187__32_,r_187__31_,r_187__30_,r_187__29_,
  r_187__28_,r_187__27_,r_187__26_,r_187__25_,r_187__24_,r_187__23_,r_187__22_,
  r_187__21_,r_187__20_,r_187__19_,r_187__18_,r_187__17_,r_187__16_,r_187__15_,
  r_187__14_,r_187__13_,r_187__12_,r_187__11_,r_187__10_,r_187__9_,r_187__8_,r_187__7_,
  r_187__6_,r_187__5_,r_187__4_,r_187__3_,r_187__2_,r_187__1_,r_187__0_,r_188__63_,
  r_188__62_,r_188__61_,r_188__60_,r_188__59_,r_188__58_,r_188__57_,r_188__56_,
  r_188__55_,r_188__54_,r_188__53_,r_188__52_,r_188__51_,r_188__50_,r_188__49_,
  r_188__48_,r_188__47_,r_188__46_,r_188__45_,r_188__44_,r_188__43_,r_188__42_,r_188__41_,
  r_188__40_,r_188__39_,r_188__38_,r_188__37_,r_188__36_,r_188__35_,r_188__34_,
  r_188__33_,r_188__32_,r_188__31_,r_188__30_,r_188__29_,r_188__28_,r_188__27_,
  r_188__26_,r_188__25_,r_188__24_,r_188__23_,r_188__22_,r_188__21_,r_188__20_,
  r_188__19_,r_188__18_,r_188__17_,r_188__16_,r_188__15_,r_188__14_,r_188__13_,r_188__12_,
  r_188__11_,r_188__10_,r_188__9_,r_188__8_,r_188__7_,r_188__6_,r_188__5_,r_188__4_,
  r_188__3_,r_188__2_,r_188__1_,r_188__0_,r_189__63_,r_189__62_,r_189__61_,
  r_189__60_,r_189__59_,r_189__58_,r_189__57_,r_189__56_,r_189__55_,r_189__54_,
  r_189__53_,r_189__52_,r_189__51_,r_189__50_,r_189__49_,r_189__48_,r_189__47_,r_189__46_,
  r_189__45_,r_189__44_,r_189__43_,r_189__42_,r_189__41_,r_189__40_,r_189__39_,
  r_189__38_,r_189__37_,r_189__36_,r_189__35_,r_189__34_,r_189__33_,r_189__32_,
  r_189__31_,r_189__30_,r_189__29_,r_189__28_,r_189__27_,r_189__26_,r_189__25_,r_189__24_,
  r_189__23_,r_189__22_,r_189__21_,r_189__20_,r_189__19_,r_189__18_,r_189__17_,
  r_189__16_,r_189__15_,r_189__14_,r_189__13_,r_189__12_,r_189__11_,r_189__10_,
  r_189__9_,r_189__8_,r_189__7_,r_189__6_,r_189__5_,r_189__4_,r_189__3_,r_189__2_,
  r_189__1_,r_189__0_,r_190__63_,r_190__62_,r_190__61_,r_190__60_,r_190__59_,r_190__58_,
  r_190__57_,r_190__56_,r_190__55_,r_190__54_,r_190__53_,r_190__52_,r_190__51_,
  r_190__50_,r_190__49_,r_190__48_,r_190__47_,r_190__46_,r_190__45_,r_190__44_,
  r_190__43_,r_190__42_,r_190__41_,r_190__40_,r_190__39_,r_190__38_,r_190__37_,
  r_190__36_,r_190__35_,r_190__34_,r_190__33_,r_190__32_,r_190__31_,r_190__30_,r_190__29_,
  r_190__28_,r_190__27_,r_190__26_,r_190__25_,r_190__24_,r_190__23_,r_190__22_,
  r_190__21_,r_190__20_,r_190__19_,r_190__18_,r_190__17_,r_190__16_,r_190__15_,
  r_190__14_,r_190__13_,r_190__12_,r_190__11_,r_190__10_,r_190__9_,r_190__8_,r_190__7_,
  r_190__6_,r_190__5_,r_190__4_,r_190__3_,r_190__2_,r_190__1_,r_190__0_,r_191__63_,
  r_191__62_,r_191__61_,r_191__60_,r_191__59_,r_191__58_,r_191__57_,r_191__56_,
  r_191__55_,r_191__54_,r_191__53_,r_191__52_,r_191__51_,r_191__50_,r_191__49_,
  r_191__48_,r_191__47_,r_191__46_,r_191__45_,r_191__44_,r_191__43_,r_191__42_,
  r_191__41_,r_191__40_,r_191__39_,r_191__38_,r_191__37_,r_191__36_,r_191__35_,r_191__34_,
  r_191__33_,r_191__32_,r_191__31_,r_191__30_,r_191__29_,r_191__28_,r_191__27_,
  r_191__26_,r_191__25_,r_191__24_,r_191__23_,r_191__22_,r_191__21_,r_191__20_,
  r_191__19_,r_191__18_,r_191__17_,r_191__16_,r_191__15_,r_191__14_,r_191__13_,r_191__12_,
  r_191__11_,r_191__10_,r_191__9_,r_191__8_,r_191__7_,r_191__6_,r_191__5_,
  r_191__4_,r_191__3_,r_191__2_,r_191__1_,r_191__0_,r_192__63_,r_192__62_,r_192__61_,
  r_192__60_,r_192__59_,r_192__58_,r_192__57_,r_192__56_,r_192__55_,r_192__54_,
  r_192__53_,r_192__52_,r_192__51_,r_192__50_,r_192__49_,r_192__48_,r_192__47_,r_192__46_,
  r_192__45_,r_192__44_,r_192__43_,r_192__42_,r_192__41_,r_192__40_,r_192__39_,
  r_192__38_,r_192__37_,r_192__36_,r_192__35_,r_192__34_,r_192__33_,r_192__32_,
  r_192__31_,r_192__30_,r_192__29_,r_192__28_,r_192__27_,r_192__26_,r_192__25_,
  r_192__24_,r_192__23_,r_192__22_,r_192__21_,r_192__20_,r_192__19_,r_192__18_,r_192__17_,
  r_192__16_,r_192__15_,r_192__14_,r_192__13_,r_192__12_,r_192__11_,r_192__10_,
  r_192__9_,r_192__8_,r_192__7_,r_192__6_,r_192__5_,r_192__4_,r_192__3_,r_192__2_,
  r_192__1_,r_192__0_,r_193__63_,r_193__62_,r_193__61_,r_193__60_,r_193__59_,
  r_193__58_,r_193__57_,r_193__56_,r_193__55_,r_193__54_,r_193__53_,r_193__52_,r_193__51_,
  r_193__50_,r_193__49_,r_193__48_,r_193__47_,r_193__46_,r_193__45_,r_193__44_,
  r_193__43_,r_193__42_,r_193__41_,r_193__40_,r_193__39_,r_193__38_,r_193__37_,
  r_193__36_,r_193__35_,r_193__34_,r_193__33_,r_193__32_,r_193__31_,r_193__30_,
  r_193__29_,r_193__28_,r_193__27_,r_193__26_,r_193__25_,r_193__24_,r_193__23_,r_193__22_,
  r_193__21_,r_193__20_,r_193__19_,r_193__18_,r_193__17_,r_193__16_,r_193__15_,
  r_193__14_,r_193__13_,r_193__12_,r_193__11_,r_193__10_,r_193__9_,r_193__8_,r_193__7_,
  r_193__6_,r_193__5_,r_193__4_,r_193__3_,r_193__2_,r_193__1_,r_193__0_,
  r_194__63_,r_194__62_,r_194__61_,r_194__60_,r_194__59_,r_194__58_,r_194__57_,r_194__56_,
  r_194__55_,r_194__54_,r_194__53_,r_194__52_,r_194__51_,r_194__50_,r_194__49_,
  r_194__48_,r_194__47_,r_194__46_,r_194__45_,r_194__44_,r_194__43_,r_194__42_,
  r_194__41_,r_194__40_,r_194__39_,r_194__38_,r_194__37_,r_194__36_,r_194__35_,r_194__34_,
  r_194__33_,r_194__32_,r_194__31_,r_194__30_,r_194__29_,r_194__28_,r_194__27_,
  r_194__26_,r_194__25_,r_194__24_,r_194__23_,r_194__22_,r_194__21_,r_194__20_,
  r_194__19_,r_194__18_,r_194__17_,r_194__16_,r_194__15_,r_194__14_,r_194__13_,
  r_194__12_,r_194__11_,r_194__10_,r_194__9_,r_194__8_,r_194__7_,r_194__6_,r_194__5_,
  r_194__4_,r_194__3_,r_194__2_,r_194__1_,r_194__0_,r_195__63_,r_195__62_,r_195__61_,
  r_195__60_,r_195__59_,r_195__58_,r_195__57_,r_195__56_,r_195__55_,r_195__54_,
  r_195__53_,r_195__52_,r_195__51_,r_195__50_,r_195__49_,r_195__48_,r_195__47_,
  r_195__46_,r_195__45_,r_195__44_,r_195__43_,r_195__42_,r_195__41_,r_195__40_,r_195__39_,
  r_195__38_,r_195__37_,r_195__36_,r_195__35_,r_195__34_,r_195__33_,r_195__32_,
  r_195__31_,r_195__30_,r_195__29_,r_195__28_,r_195__27_,r_195__26_,r_195__25_,
  r_195__24_,r_195__23_,r_195__22_,r_195__21_,r_195__20_,r_195__19_,r_195__18_,
  r_195__17_,r_195__16_,r_195__15_,r_195__14_,r_195__13_,r_195__12_,r_195__11_,r_195__10_,
  r_195__9_,r_195__8_,r_195__7_,r_195__6_,r_195__5_,r_195__4_,r_195__3_,r_195__2_,
  r_195__1_,r_195__0_,r_196__63_,r_196__62_,r_196__61_,r_196__60_,r_196__59_,
  r_196__58_,r_196__57_,r_196__56_,r_196__55_,r_196__54_,r_196__53_,r_196__52_,
  r_196__51_,r_196__50_,r_196__49_,r_196__48_,r_196__47_,r_196__46_,r_196__45_,r_196__44_,
  r_196__43_,r_196__42_,r_196__41_,r_196__40_,r_196__39_,r_196__38_,r_196__37_,
  r_196__36_,r_196__35_,r_196__34_,r_196__33_,r_196__32_,r_196__31_,r_196__30_,
  r_196__29_,r_196__28_,r_196__27_,r_196__26_,r_196__25_,r_196__24_,r_196__23_,r_196__22_,
  r_196__21_,r_196__20_,r_196__19_,r_196__18_,r_196__17_,r_196__16_,r_196__15_,
  r_196__14_,r_196__13_,r_196__12_,r_196__11_,r_196__10_,r_196__9_,r_196__8_,
  r_196__7_,r_196__6_,r_196__5_,r_196__4_,r_196__3_,r_196__2_,r_196__1_,r_196__0_,
  r_197__63_,r_197__62_,r_197__61_,r_197__60_,r_197__59_,r_197__58_,r_197__57_,r_197__56_,
  r_197__55_,r_197__54_,r_197__53_,r_197__52_,r_197__51_,r_197__50_,r_197__49_,
  r_197__48_,r_197__47_,r_197__46_,r_197__45_,r_197__44_,r_197__43_,r_197__42_,
  r_197__41_,r_197__40_,r_197__39_,r_197__38_,r_197__37_,r_197__36_,r_197__35_,
  r_197__34_,r_197__33_,r_197__32_,r_197__31_,r_197__30_,r_197__29_,r_197__28_,r_197__27_,
  r_197__26_,r_197__25_,r_197__24_,r_197__23_,r_197__22_,r_197__21_,r_197__20_,
  r_197__19_,r_197__18_,r_197__17_,r_197__16_,r_197__15_,r_197__14_,r_197__13_,
  r_197__12_,r_197__11_,r_197__10_,r_197__9_,r_197__8_,r_197__7_,r_197__6_,r_197__5_,
  r_197__4_,r_197__3_,r_197__2_,r_197__1_,r_197__0_,r_198__63_,r_198__62_,r_198__61_,
  r_198__60_,r_198__59_,r_198__58_,r_198__57_,r_198__56_,r_198__55_,r_198__54_,
  r_198__53_,r_198__52_,r_198__51_,r_198__50_,r_198__49_,r_198__48_,r_198__47_,
  r_198__46_,r_198__45_,r_198__44_,r_198__43_,r_198__42_,r_198__41_,r_198__40_,
  r_198__39_,r_198__38_,r_198__37_,r_198__36_,r_198__35_,r_198__34_,r_198__33_,r_198__32_,
  r_198__31_,r_198__30_,r_198__29_,r_198__28_,r_198__27_,r_198__26_,r_198__25_,
  r_198__24_,r_198__23_,r_198__22_,r_198__21_,r_198__20_,r_198__19_,r_198__18_,
  r_198__17_,r_198__16_,r_198__15_,r_198__14_,r_198__13_,r_198__12_,r_198__11_,r_198__10_,
  r_198__9_,r_198__8_,r_198__7_,r_198__6_,r_198__5_,r_198__4_,r_198__3_,r_198__2_,
  r_198__1_,r_198__0_,r_199__63_,r_199__62_,r_199__61_,r_199__60_,r_199__59_,
  r_199__58_,r_199__57_,r_199__56_,r_199__55_,r_199__54_,r_199__53_,r_199__52_,
  r_199__51_,r_199__50_,r_199__49_,r_199__48_,r_199__47_,r_199__46_,r_199__45_,r_199__44_,
  r_199__43_,r_199__42_,r_199__41_,r_199__40_,r_199__39_,r_199__38_,r_199__37_,
  r_199__36_,r_199__35_,r_199__34_,r_199__33_,r_199__32_,r_199__31_,r_199__30_,
  r_199__29_,r_199__28_,r_199__27_,r_199__26_,r_199__25_,r_199__24_,r_199__23_,
  r_199__22_,r_199__21_,r_199__20_,r_199__19_,r_199__18_,r_199__17_,r_199__16_,r_199__15_,
  r_199__14_,r_199__13_,r_199__12_,r_199__11_,r_199__10_,r_199__9_,r_199__8_,
  r_199__7_,r_199__6_,r_199__5_,r_199__4_,r_199__3_,r_199__2_,r_199__1_,r_199__0_,
  r_200__63_,r_200__62_,r_200__61_,r_200__60_,r_200__59_,r_200__58_,r_200__57_,
  r_200__56_,r_200__55_,r_200__54_,r_200__53_,r_200__52_,r_200__51_,r_200__50_,r_200__49_,
  r_200__48_,r_200__47_,r_200__46_,r_200__45_,r_200__44_,r_200__43_,r_200__42_,
  r_200__41_,r_200__40_,r_200__39_,r_200__38_,r_200__37_,r_200__36_,r_200__35_,
  r_200__34_,r_200__33_,r_200__32_,r_200__31_,r_200__30_,r_200__29_,r_200__28_,
  r_200__27_,r_200__26_,r_200__25_,r_200__24_,r_200__23_,r_200__22_,r_200__21_,r_200__20_,
  r_200__19_,r_200__18_,r_200__17_,r_200__16_,r_200__15_,r_200__14_,r_200__13_,
  r_200__12_,r_200__11_,r_200__10_,r_200__9_,r_200__8_,r_200__7_,r_200__6_,r_200__5_,
  r_200__4_,r_200__3_,r_200__2_,r_200__1_,r_200__0_,r_201__63_,r_201__62_,
  r_201__61_,r_201__60_,r_201__59_,r_201__58_,r_201__57_,r_201__56_,r_201__55_,r_201__54_,
  r_201__53_,r_201__52_,r_201__51_,r_201__50_,r_201__49_,r_201__48_,r_201__47_,
  r_201__46_,r_201__45_,r_201__44_,r_201__43_,r_201__42_,r_201__41_,r_201__40_,
  r_201__39_,r_201__38_,r_201__37_,r_201__36_,r_201__35_,r_201__34_,r_201__33_,r_201__32_,
  r_201__31_,r_201__30_,r_201__29_,r_201__28_,r_201__27_,r_201__26_,r_201__25_,
  r_201__24_,r_201__23_,r_201__22_,r_201__21_,r_201__20_,r_201__19_,r_201__18_,
  r_201__17_,r_201__16_,r_201__15_,r_201__14_,r_201__13_,r_201__12_,r_201__11_,
  r_201__10_,r_201__9_,r_201__8_,r_201__7_,r_201__6_,r_201__5_,r_201__4_,r_201__3_,
  r_201__2_,r_201__1_,r_201__0_,r_202__63_,r_202__62_,r_202__61_,r_202__60_,r_202__59_,
  r_202__58_,r_202__57_,r_202__56_,r_202__55_,r_202__54_,r_202__53_,r_202__52_,
  r_202__51_,r_202__50_,r_202__49_,r_202__48_,r_202__47_,r_202__46_,r_202__45_,
  r_202__44_,r_202__43_,r_202__42_,r_202__41_,r_202__40_,r_202__39_,r_202__38_,r_202__37_,
  r_202__36_,r_202__35_,r_202__34_,r_202__33_,r_202__32_,r_202__31_,r_202__30_,
  r_202__29_,r_202__28_,r_202__27_,r_202__26_,r_202__25_,r_202__24_,r_202__23_,
  r_202__22_,r_202__21_,r_202__20_,r_202__19_,r_202__18_,r_202__17_,r_202__16_,
  r_202__15_,r_202__14_,r_202__13_,r_202__12_,r_202__11_,r_202__10_,r_202__9_,r_202__8_,
  r_202__7_,r_202__6_,r_202__5_,r_202__4_,r_202__3_,r_202__2_,r_202__1_,r_202__0_,
  r_203__63_,r_203__62_,r_203__61_,r_203__60_,r_203__59_,r_203__58_,r_203__57_,
  r_203__56_,r_203__55_,r_203__54_,r_203__53_,r_203__52_,r_203__51_,r_203__50_,
  r_203__49_,r_203__48_,r_203__47_,r_203__46_,r_203__45_,r_203__44_,r_203__43_,r_203__42_,
  r_203__41_,r_203__40_,r_203__39_,r_203__38_,r_203__37_,r_203__36_,r_203__35_,
  r_203__34_,r_203__33_,r_203__32_,r_203__31_,r_203__30_,r_203__29_,r_203__28_,
  r_203__27_,r_203__26_,r_203__25_,r_203__24_,r_203__23_,r_203__22_,r_203__21_,r_203__20_,
  r_203__19_,r_203__18_,r_203__17_,r_203__16_,r_203__15_,r_203__14_,r_203__13_,
  r_203__12_,r_203__11_,r_203__10_,r_203__9_,r_203__8_,r_203__7_,r_203__6_,r_203__5_,
  r_203__4_,r_203__3_,r_203__2_,r_203__1_,r_203__0_,r_204__63_,r_204__62_,
  r_204__61_,r_204__60_,r_204__59_,r_204__58_,r_204__57_,r_204__56_,r_204__55_,r_204__54_,
  r_204__53_,r_204__52_,r_204__51_,r_204__50_,r_204__49_,r_204__48_,r_204__47_,
  r_204__46_,r_204__45_,r_204__44_,r_204__43_,r_204__42_,r_204__41_,r_204__40_,
  r_204__39_,r_204__38_,r_204__37_,r_204__36_,r_204__35_,r_204__34_,r_204__33_,
  r_204__32_,r_204__31_,r_204__30_,r_204__29_,r_204__28_,r_204__27_,r_204__26_,r_204__25_,
  r_204__24_,r_204__23_,r_204__22_,r_204__21_,r_204__20_,r_204__19_,r_204__18_,
  r_204__17_,r_204__16_,r_204__15_,r_204__14_,r_204__13_,r_204__12_,r_204__11_,
  r_204__10_,r_204__9_,r_204__8_,r_204__7_,r_204__6_,r_204__5_,r_204__4_,r_204__3_,
  r_204__2_,r_204__1_,r_204__0_,r_205__63_,r_205__62_,r_205__61_,r_205__60_,r_205__59_,
  r_205__58_,r_205__57_,r_205__56_,r_205__55_,r_205__54_,r_205__53_,r_205__52_,
  r_205__51_,r_205__50_,r_205__49_,r_205__48_,r_205__47_,r_205__46_,r_205__45_,
  r_205__44_,r_205__43_,r_205__42_,r_205__41_,r_205__40_,r_205__39_,r_205__38_,
  r_205__37_,r_205__36_,r_205__35_,r_205__34_,r_205__33_,r_205__32_,r_205__31_,r_205__30_,
  r_205__29_,r_205__28_,r_205__27_,r_205__26_,r_205__25_,r_205__24_,r_205__23_,
  r_205__22_,r_205__21_,r_205__20_,r_205__19_,r_205__18_,r_205__17_,r_205__16_,
  r_205__15_,r_205__14_,r_205__13_,r_205__12_,r_205__11_,r_205__10_,r_205__9_,r_205__8_,
  r_205__7_,r_205__6_,r_205__5_,r_205__4_,r_205__3_,r_205__2_,r_205__1_,r_205__0_,
  r_206__63_,r_206__62_,r_206__61_,r_206__60_,r_206__59_,r_206__58_,r_206__57_,
  r_206__56_,r_206__55_,r_206__54_,r_206__53_,r_206__52_,r_206__51_,r_206__50_,
  r_206__49_,r_206__48_,r_206__47_,r_206__46_,r_206__45_,r_206__44_,r_206__43_,r_206__42_,
  r_206__41_,r_206__40_,r_206__39_,r_206__38_,r_206__37_,r_206__36_,r_206__35_,
  r_206__34_,r_206__33_,r_206__32_,r_206__31_,r_206__30_,r_206__29_,r_206__28_,
  r_206__27_,r_206__26_,r_206__25_,r_206__24_,r_206__23_,r_206__22_,r_206__21_,
  r_206__20_,r_206__19_,r_206__18_,r_206__17_,r_206__16_,r_206__15_,r_206__14_,r_206__13_,
  r_206__12_,r_206__11_,r_206__10_,r_206__9_,r_206__8_,r_206__7_,r_206__6_,
  r_206__5_,r_206__4_,r_206__3_,r_206__2_,r_206__1_,r_206__0_,r_207__63_,r_207__62_,
  r_207__61_,r_207__60_,r_207__59_,r_207__58_,r_207__57_,r_207__56_,r_207__55_,
  r_207__54_,r_207__53_,r_207__52_,r_207__51_,r_207__50_,r_207__49_,r_207__48_,r_207__47_,
  r_207__46_,r_207__45_,r_207__44_,r_207__43_,r_207__42_,r_207__41_,r_207__40_,
  r_207__39_,r_207__38_,r_207__37_,r_207__36_,r_207__35_,r_207__34_,r_207__33_,
  r_207__32_,r_207__31_,r_207__30_,r_207__29_,r_207__28_,r_207__27_,r_207__26_,
  r_207__25_,r_207__24_,r_207__23_,r_207__22_,r_207__21_,r_207__20_,r_207__19_,r_207__18_,
  r_207__17_,r_207__16_,r_207__15_,r_207__14_,r_207__13_,r_207__12_,r_207__11_,
  r_207__10_,r_207__9_,r_207__8_,r_207__7_,r_207__6_,r_207__5_,r_207__4_,r_207__3_,
  r_207__2_,r_207__1_,r_207__0_,r_208__63_,r_208__62_,r_208__61_,r_208__60_,
  r_208__59_,r_208__58_,r_208__57_,r_208__56_,r_208__55_,r_208__54_,r_208__53_,r_208__52_,
  r_208__51_,r_208__50_,r_208__49_,r_208__48_,r_208__47_,r_208__46_,r_208__45_,
  r_208__44_,r_208__43_,r_208__42_,r_208__41_,r_208__40_,r_208__39_,r_208__38_,
  r_208__37_,r_208__36_,r_208__35_,r_208__34_,r_208__33_,r_208__32_,r_208__31_,r_208__30_,
  r_208__29_,r_208__28_,r_208__27_,r_208__26_,r_208__25_,r_208__24_,r_208__23_,
  r_208__22_,r_208__21_,r_208__20_,r_208__19_,r_208__18_,r_208__17_,r_208__16_,
  r_208__15_,r_208__14_,r_208__13_,r_208__12_,r_208__11_,r_208__10_,r_208__9_,r_208__8_,
  r_208__7_,r_208__6_,r_208__5_,r_208__4_,r_208__3_,r_208__2_,r_208__1_,r_208__0_,
  r_209__63_,r_209__62_,r_209__61_,r_209__60_,r_209__59_,r_209__58_,r_209__57_,
  r_209__56_,r_209__55_,r_209__54_,r_209__53_,r_209__52_,r_209__51_,r_209__50_,
  r_209__49_,r_209__48_,r_209__47_,r_209__46_,r_209__45_,r_209__44_,r_209__43_,
  r_209__42_,r_209__41_,r_209__40_,r_209__39_,r_209__38_,r_209__37_,r_209__36_,r_209__35_,
  r_209__34_,r_209__33_,r_209__32_,r_209__31_,r_209__30_,r_209__29_,r_209__28_,
  r_209__27_,r_209__26_,r_209__25_,r_209__24_,r_209__23_,r_209__22_,r_209__21_,
  r_209__20_,r_209__19_,r_209__18_,r_209__17_,r_209__16_,r_209__15_,r_209__14_,
  r_209__13_,r_209__12_,r_209__11_,r_209__10_,r_209__9_,r_209__8_,r_209__7_,r_209__6_,
  r_209__5_,r_209__4_,r_209__3_,r_209__2_,r_209__1_,r_209__0_,r_210__63_,r_210__62_,
  r_210__61_,r_210__60_,r_210__59_,r_210__58_,r_210__57_,r_210__56_,r_210__55_,
  r_210__54_,r_210__53_,r_210__52_,r_210__51_,r_210__50_,r_210__49_,r_210__48_,
  r_210__47_,r_210__46_,r_210__45_,r_210__44_,r_210__43_,r_210__42_,r_210__41_,r_210__40_,
  r_210__39_,r_210__38_,r_210__37_,r_210__36_,r_210__35_,r_210__34_,r_210__33_,
  r_210__32_,r_210__31_,r_210__30_,r_210__29_,r_210__28_,r_210__27_,r_210__26_,
  r_210__25_,r_210__24_,r_210__23_,r_210__22_,r_210__21_,r_210__20_,r_210__19_,r_210__18_,
  r_210__17_,r_210__16_,r_210__15_,r_210__14_,r_210__13_,r_210__12_,r_210__11_,
  r_210__10_,r_210__9_,r_210__8_,r_210__7_,r_210__6_,r_210__5_,r_210__4_,r_210__3_,
  r_210__2_,r_210__1_,r_210__0_,r_211__63_,r_211__62_,r_211__61_,r_211__60_,
  r_211__59_,r_211__58_,r_211__57_,r_211__56_,r_211__55_,r_211__54_,r_211__53_,r_211__52_,
  r_211__51_,r_211__50_,r_211__49_,r_211__48_,r_211__47_,r_211__46_,r_211__45_,
  r_211__44_,r_211__43_,r_211__42_,r_211__41_,r_211__40_,r_211__39_,r_211__38_,
  r_211__37_,r_211__36_,r_211__35_,r_211__34_,r_211__33_,r_211__32_,r_211__31_,
  r_211__30_,r_211__29_,r_211__28_,r_211__27_,r_211__26_,r_211__25_,r_211__24_,r_211__23_,
  r_211__22_,r_211__21_,r_211__20_,r_211__19_,r_211__18_,r_211__17_,r_211__16_,
  r_211__15_,r_211__14_,r_211__13_,r_211__12_,r_211__11_,r_211__10_,r_211__9_,
  r_211__8_,r_211__7_,r_211__6_,r_211__5_,r_211__4_,r_211__3_,r_211__2_,r_211__1_,
  r_211__0_,r_212__63_,r_212__62_,r_212__61_,r_212__60_,r_212__59_,r_212__58_,r_212__57_,
  r_212__56_,r_212__55_,r_212__54_,r_212__53_,r_212__52_,r_212__51_,r_212__50_,
  r_212__49_,r_212__48_,r_212__47_,r_212__46_,r_212__45_,r_212__44_,r_212__43_,
  r_212__42_,r_212__41_,r_212__40_,r_212__39_,r_212__38_,r_212__37_,r_212__36_,
  r_212__35_,r_212__34_,r_212__33_,r_212__32_,r_212__31_,r_212__30_,r_212__29_,r_212__28_,
  r_212__27_,r_212__26_,r_212__25_,r_212__24_,r_212__23_,r_212__22_,r_212__21_,
  r_212__20_,r_212__19_,r_212__18_,r_212__17_,r_212__16_,r_212__15_,r_212__14_,
  r_212__13_,r_212__12_,r_212__11_,r_212__10_,r_212__9_,r_212__8_,r_212__7_,r_212__6_,
  r_212__5_,r_212__4_,r_212__3_,r_212__2_,r_212__1_,r_212__0_,r_213__63_,r_213__62_,
  r_213__61_,r_213__60_,r_213__59_,r_213__58_,r_213__57_,r_213__56_,r_213__55_,
  r_213__54_,r_213__53_,r_213__52_,r_213__51_,r_213__50_,r_213__49_,r_213__48_,
  r_213__47_,r_213__46_,r_213__45_,r_213__44_,r_213__43_,r_213__42_,r_213__41_,r_213__40_,
  r_213__39_,r_213__38_,r_213__37_,r_213__36_,r_213__35_,r_213__34_,r_213__33_,
  r_213__32_,r_213__31_,r_213__30_,r_213__29_,r_213__28_,r_213__27_,r_213__26_,
  r_213__25_,r_213__24_,r_213__23_,r_213__22_,r_213__21_,r_213__20_,r_213__19_,
  r_213__18_,r_213__17_,r_213__16_,r_213__15_,r_213__14_,r_213__13_,r_213__12_,r_213__11_,
  r_213__10_,r_213__9_,r_213__8_,r_213__7_,r_213__6_,r_213__5_,r_213__4_,r_213__3_,
  r_213__2_,r_213__1_,r_213__0_,r_214__63_,r_214__62_,r_214__61_,r_214__60_,
  r_214__59_,r_214__58_,r_214__57_,r_214__56_,r_214__55_,r_214__54_,r_214__53_,
  r_214__52_,r_214__51_,r_214__50_,r_214__49_,r_214__48_,r_214__47_,r_214__46_,r_214__45_,
  r_214__44_,r_214__43_,r_214__42_,r_214__41_,r_214__40_,r_214__39_,r_214__38_,
  r_214__37_,r_214__36_,r_214__35_,r_214__34_,r_214__33_,r_214__32_,r_214__31_,
  r_214__30_,r_214__29_,r_214__28_,r_214__27_,r_214__26_,r_214__25_,r_214__24_,
  r_214__23_,r_214__22_,r_214__21_,r_214__20_,r_214__19_,r_214__18_,r_214__17_,r_214__16_,
  r_214__15_,r_214__14_,r_214__13_,r_214__12_,r_214__11_,r_214__10_,r_214__9_,
  r_214__8_,r_214__7_,r_214__6_,r_214__5_,r_214__4_,r_214__3_,r_214__2_,r_214__1_,
  r_214__0_,r_215__63_,r_215__62_,r_215__61_,r_215__60_,r_215__59_,r_215__58_,
  r_215__57_,r_215__56_,r_215__55_,r_215__54_,r_215__53_,r_215__52_,r_215__51_,r_215__50_,
  r_215__49_,r_215__48_,r_215__47_,r_215__46_,r_215__45_,r_215__44_,r_215__43_,
  r_215__42_,r_215__41_,r_215__40_,r_215__39_,r_215__38_,r_215__37_,r_215__36_,
  r_215__35_,r_215__34_,r_215__33_,r_215__32_,r_215__31_,r_215__30_,r_215__29_,r_215__28_,
  r_215__27_,r_215__26_,r_215__25_,r_215__24_,r_215__23_,r_215__22_,r_215__21_,
  r_215__20_,r_215__19_,r_215__18_,r_215__17_,r_215__16_,r_215__15_,r_215__14_,
  r_215__13_,r_215__12_,r_215__11_,r_215__10_,r_215__9_,r_215__8_,r_215__7_,r_215__6_,
  r_215__5_,r_215__4_,r_215__3_,r_215__2_,r_215__1_,r_215__0_,r_216__63_,r_216__62_,
  r_216__61_,r_216__60_,r_216__59_,r_216__58_,r_216__57_,r_216__56_,r_216__55_,
  r_216__54_,r_216__53_,r_216__52_,r_216__51_,r_216__50_,r_216__49_,r_216__48_,
  r_216__47_,r_216__46_,r_216__45_,r_216__44_,r_216__43_,r_216__42_,r_216__41_,
  r_216__40_,r_216__39_,r_216__38_,r_216__37_,r_216__36_,r_216__35_,r_216__34_,r_216__33_,
  r_216__32_,r_216__31_,r_216__30_,r_216__29_,r_216__28_,r_216__27_,r_216__26_,
  r_216__25_,r_216__24_,r_216__23_,r_216__22_,r_216__21_,r_216__20_,r_216__19_,
  r_216__18_,r_216__17_,r_216__16_,r_216__15_,r_216__14_,r_216__13_,r_216__12_,
  r_216__11_,r_216__10_,r_216__9_,r_216__8_,r_216__7_,r_216__6_,r_216__5_,r_216__4_,
  r_216__3_,r_216__2_,r_216__1_,r_216__0_,r_217__63_,r_217__62_,r_217__61_,r_217__60_,
  r_217__59_,r_217__58_,r_217__57_,r_217__56_,r_217__55_,r_217__54_,r_217__53_,
  r_217__52_,r_217__51_,r_217__50_,r_217__49_,r_217__48_,r_217__47_,r_217__46_,
  r_217__45_,r_217__44_,r_217__43_,r_217__42_,r_217__41_,r_217__40_,r_217__39_,r_217__38_,
  r_217__37_,r_217__36_,r_217__35_,r_217__34_,r_217__33_,r_217__32_,r_217__31_,
  r_217__30_,r_217__29_,r_217__28_,r_217__27_,r_217__26_,r_217__25_,r_217__24_,
  r_217__23_,r_217__22_,r_217__21_,r_217__20_,r_217__19_,r_217__18_,r_217__17_,r_217__16_,
  r_217__15_,r_217__14_,r_217__13_,r_217__12_,r_217__11_,r_217__10_,r_217__9_,
  r_217__8_,r_217__7_,r_217__6_,r_217__5_,r_217__4_,r_217__3_,r_217__2_,r_217__1_,
  r_217__0_,r_218__63_,r_218__62_,r_218__61_,r_218__60_,r_218__59_,r_218__58_,
  r_218__57_,r_218__56_,r_218__55_,r_218__54_,r_218__53_,r_218__52_,r_218__51_,r_218__50_,
  r_218__49_,r_218__48_,r_218__47_,r_218__46_,r_218__45_,r_218__44_,r_218__43_,
  r_218__42_,r_218__41_,r_218__40_,r_218__39_,r_218__38_,r_218__37_,r_218__36_,
  r_218__35_,r_218__34_,r_218__33_,r_218__32_,r_218__31_,r_218__30_,r_218__29_,
  r_218__28_,r_218__27_,r_218__26_,r_218__25_,r_218__24_,r_218__23_,r_218__22_,r_218__21_,
  r_218__20_,r_218__19_,r_218__18_,r_218__17_,r_218__16_,r_218__15_,r_218__14_,
  r_218__13_,r_218__12_,r_218__11_,r_218__10_,r_218__9_,r_218__8_,r_218__7_,r_218__6_,
  r_218__5_,r_218__4_,r_218__3_,r_218__2_,r_218__1_,r_218__0_,r_219__63_,
  r_219__62_,r_219__61_,r_219__60_,r_219__59_,r_219__58_,r_219__57_,r_219__56_,r_219__55_,
  r_219__54_,r_219__53_,r_219__52_,r_219__51_,r_219__50_,r_219__49_,r_219__48_,
  r_219__47_,r_219__46_,r_219__45_,r_219__44_,r_219__43_,r_219__42_,r_219__41_,
  r_219__40_,r_219__39_,r_219__38_,r_219__37_,r_219__36_,r_219__35_,r_219__34_,
  r_219__33_,r_219__32_,r_219__31_,r_219__30_,r_219__29_,r_219__28_,r_219__27_,r_219__26_,
  r_219__25_,r_219__24_,r_219__23_,r_219__22_,r_219__21_,r_219__20_,r_219__19_,
  r_219__18_,r_219__17_,r_219__16_,r_219__15_,r_219__14_,r_219__13_,r_219__12_,
  r_219__11_,r_219__10_,r_219__9_,r_219__8_,r_219__7_,r_219__6_,r_219__5_,r_219__4_,
  r_219__3_,r_219__2_,r_219__1_,r_219__0_,r_220__63_,r_220__62_,r_220__61_,r_220__60_,
  r_220__59_,r_220__58_,r_220__57_,r_220__56_,r_220__55_,r_220__54_,r_220__53_,
  r_220__52_,r_220__51_,r_220__50_,r_220__49_,r_220__48_,r_220__47_,r_220__46_,
  r_220__45_,r_220__44_,r_220__43_,r_220__42_,r_220__41_,r_220__40_,r_220__39_,r_220__38_,
  r_220__37_,r_220__36_,r_220__35_,r_220__34_,r_220__33_,r_220__32_,r_220__31_,
  r_220__30_,r_220__29_,r_220__28_,r_220__27_,r_220__26_,r_220__25_,r_220__24_,
  r_220__23_,r_220__22_,r_220__21_,r_220__20_,r_220__19_,r_220__18_,r_220__17_,
  r_220__16_,r_220__15_,r_220__14_,r_220__13_,r_220__12_,r_220__11_,r_220__10_,r_220__9_,
  r_220__8_,r_220__7_,r_220__6_,r_220__5_,r_220__4_,r_220__3_,r_220__2_,r_220__1_,
  r_220__0_,r_221__63_,r_221__62_,r_221__61_,r_221__60_,r_221__59_,r_221__58_,
  r_221__57_,r_221__56_,r_221__55_,r_221__54_,r_221__53_,r_221__52_,r_221__51_,
  r_221__50_,r_221__49_,r_221__48_,r_221__47_,r_221__46_,r_221__45_,r_221__44_,r_221__43_,
  r_221__42_,r_221__41_,r_221__40_,r_221__39_,r_221__38_,r_221__37_,r_221__36_,
  r_221__35_,r_221__34_,r_221__33_,r_221__32_,r_221__31_,r_221__30_,r_221__29_,
  r_221__28_,r_221__27_,r_221__26_,r_221__25_,r_221__24_,r_221__23_,r_221__22_,
  r_221__21_,r_221__20_,r_221__19_,r_221__18_,r_221__17_,r_221__16_,r_221__15_,r_221__14_,
  r_221__13_,r_221__12_,r_221__11_,r_221__10_,r_221__9_,r_221__8_,r_221__7_,
  r_221__6_,r_221__5_,r_221__4_,r_221__3_,r_221__2_,r_221__1_,r_221__0_,r_222__63_,
  r_222__62_,r_222__61_,r_222__60_,r_222__59_,r_222__58_,r_222__57_,r_222__56_,
  r_222__55_,r_222__54_,r_222__53_,r_222__52_,r_222__51_,r_222__50_,r_222__49_,r_222__48_,
  r_222__47_,r_222__46_,r_222__45_,r_222__44_,r_222__43_,r_222__42_,r_222__41_,
  r_222__40_,r_222__39_,r_222__38_,r_222__37_,r_222__36_,r_222__35_,r_222__34_,
  r_222__33_,r_222__32_,r_222__31_,r_222__30_,r_222__29_,r_222__28_,r_222__27_,r_222__26_,
  r_222__25_,r_222__24_,r_222__23_,r_222__22_,r_222__21_,r_222__20_,r_222__19_,
  r_222__18_,r_222__17_,r_222__16_,r_222__15_,r_222__14_,r_222__13_,r_222__12_,
  r_222__11_,r_222__10_,r_222__9_,r_222__8_,r_222__7_,r_222__6_,r_222__5_,r_222__4_,
  r_222__3_,r_222__2_,r_222__1_,r_222__0_,r_223__63_,r_223__62_,r_223__61_,r_223__60_,
  r_223__59_,r_223__58_,r_223__57_,r_223__56_,r_223__55_,r_223__54_,r_223__53_,
  r_223__52_,r_223__51_,r_223__50_,r_223__49_,r_223__48_,r_223__47_,r_223__46_,
  r_223__45_,r_223__44_,r_223__43_,r_223__42_,r_223__41_,r_223__40_,r_223__39_,
  r_223__38_,r_223__37_,r_223__36_,r_223__35_,r_223__34_,r_223__33_,r_223__32_,r_223__31_,
  r_223__30_,r_223__29_,r_223__28_,r_223__27_,r_223__26_,r_223__25_,r_223__24_,
  r_223__23_,r_223__22_,r_223__21_,r_223__20_,r_223__19_,r_223__18_,r_223__17_,
  r_223__16_,r_223__15_,r_223__14_,r_223__13_,r_223__12_,r_223__11_,r_223__10_,r_223__9_,
  r_223__8_,r_223__7_,r_223__6_,r_223__5_,r_223__4_,r_223__3_,r_223__2_,r_223__1_,
  r_223__0_,r_224__63_,r_224__62_,r_224__61_,r_224__60_,r_224__59_,r_224__58_,
  r_224__57_,r_224__56_,r_224__55_,r_224__54_,r_224__53_,r_224__52_,r_224__51_,
  r_224__50_,r_224__49_,r_224__48_,r_224__47_,r_224__46_,r_224__45_,r_224__44_,
  r_224__43_,r_224__42_,r_224__41_,r_224__40_,r_224__39_,r_224__38_,r_224__37_,r_224__36_,
  r_224__35_,r_224__34_,r_224__33_,r_224__32_,r_224__31_,r_224__30_,r_224__29_,
  r_224__28_,r_224__27_,r_224__26_,r_224__25_,r_224__24_,r_224__23_,r_224__22_,
  r_224__21_,r_224__20_,r_224__19_,r_224__18_,r_224__17_,r_224__16_,r_224__15_,r_224__14_,
  r_224__13_,r_224__12_,r_224__11_,r_224__10_,r_224__9_,r_224__8_,r_224__7_,
  r_224__6_,r_224__5_,r_224__4_,r_224__3_,r_224__2_,r_224__1_,r_224__0_,r_225__63_,
  r_225__62_,r_225__61_,r_225__60_,r_225__59_,r_225__58_,r_225__57_,r_225__56_,
  r_225__55_,r_225__54_,r_225__53_,r_225__52_,r_225__51_,r_225__50_,r_225__49_,r_225__48_,
  r_225__47_,r_225__46_,r_225__45_,r_225__44_,r_225__43_,r_225__42_,r_225__41_,
  r_225__40_,r_225__39_,r_225__38_,r_225__37_,r_225__36_,r_225__35_,r_225__34_,
  r_225__33_,r_225__32_,r_225__31_,r_225__30_,r_225__29_,r_225__28_,r_225__27_,
  r_225__26_,r_225__25_,r_225__24_,r_225__23_,r_225__22_,r_225__21_,r_225__20_,r_225__19_,
  r_225__18_,r_225__17_,r_225__16_,r_225__15_,r_225__14_,r_225__13_,r_225__12_,
  r_225__11_,r_225__10_,r_225__9_,r_225__8_,r_225__7_,r_225__6_,r_225__5_,r_225__4_,
  r_225__3_,r_225__2_,r_225__1_,r_225__0_,r_226__63_,r_226__62_,r_226__61_,
  r_226__60_,r_226__59_,r_226__58_,r_226__57_,r_226__56_,r_226__55_,r_226__54_,r_226__53_,
  r_226__52_,r_226__51_,r_226__50_,r_226__49_,r_226__48_,r_226__47_,r_226__46_,
  r_226__45_,r_226__44_,r_226__43_,r_226__42_,r_226__41_,r_226__40_,r_226__39_,
  r_226__38_,r_226__37_,r_226__36_,r_226__35_,r_226__34_,r_226__33_,r_226__32_,
  r_226__31_,r_226__30_,r_226__29_,r_226__28_,r_226__27_,r_226__26_,r_226__25_,r_226__24_,
  r_226__23_,r_226__22_,r_226__21_,r_226__20_,r_226__19_,r_226__18_,r_226__17_,
  r_226__16_,r_226__15_,r_226__14_,r_226__13_,r_226__12_,r_226__11_,r_226__10_,
  r_226__9_,r_226__8_,r_226__7_,r_226__6_,r_226__5_,r_226__4_,r_226__3_,r_226__2_,
  r_226__1_,r_226__0_,r_227__63_,r_227__62_,r_227__61_,r_227__60_,r_227__59_,r_227__58_,
  r_227__57_,r_227__56_,r_227__55_,r_227__54_,r_227__53_,r_227__52_,r_227__51_,
  r_227__50_,r_227__49_,r_227__48_,r_227__47_,r_227__46_,r_227__45_,r_227__44_,
  r_227__43_,r_227__42_,r_227__41_,r_227__40_,r_227__39_,r_227__38_,r_227__37_,r_227__36_,
  r_227__35_,r_227__34_,r_227__33_,r_227__32_,r_227__31_,r_227__30_,r_227__29_,
  r_227__28_,r_227__27_,r_227__26_,r_227__25_,r_227__24_,r_227__23_,r_227__22_,
  r_227__21_,r_227__20_,r_227__19_,r_227__18_,r_227__17_,r_227__16_,r_227__15_,
  r_227__14_,r_227__13_,r_227__12_,r_227__11_,r_227__10_,r_227__9_,r_227__8_,r_227__7_,
  r_227__6_,r_227__5_,r_227__4_,r_227__3_,r_227__2_,r_227__1_,r_227__0_,r_228__63_,
  r_228__62_,r_228__61_,r_228__60_,r_228__59_,r_228__58_,r_228__57_,r_228__56_,
  r_228__55_,r_228__54_,r_228__53_,r_228__52_,r_228__51_,r_228__50_,r_228__49_,
  r_228__48_,r_228__47_,r_228__46_,r_228__45_,r_228__44_,r_228__43_,r_228__42_,r_228__41_,
  r_228__40_,r_228__39_,r_228__38_,r_228__37_,r_228__36_,r_228__35_,r_228__34_,
  r_228__33_,r_228__32_,r_228__31_,r_228__30_,r_228__29_,r_228__28_,r_228__27_,
  r_228__26_,r_228__25_,r_228__24_,r_228__23_,r_228__22_,r_228__21_,r_228__20_,
  r_228__19_,r_228__18_,r_228__17_,r_228__16_,r_228__15_,r_228__14_,r_228__13_,r_228__12_,
  r_228__11_,r_228__10_,r_228__9_,r_228__8_,r_228__7_,r_228__6_,r_228__5_,r_228__4_,
  r_228__3_,r_228__2_,r_228__1_,r_228__0_,r_229__63_,r_229__62_,r_229__61_,
  r_229__60_,r_229__59_,r_229__58_,r_229__57_,r_229__56_,r_229__55_,r_229__54_,
  r_229__53_,r_229__52_,r_229__51_,r_229__50_,r_229__49_,r_229__48_,r_229__47_,r_229__46_,
  r_229__45_,r_229__44_,r_229__43_,r_229__42_,r_229__41_,r_229__40_,r_229__39_,
  r_229__38_,r_229__37_,r_229__36_,r_229__35_,r_229__34_,r_229__33_,r_229__32_,
  r_229__31_,r_229__30_,r_229__29_,r_229__28_,r_229__27_,r_229__26_,r_229__25_,r_229__24_,
  r_229__23_,r_229__22_,r_229__21_,r_229__20_,r_229__19_,r_229__18_,r_229__17_,
  r_229__16_,r_229__15_,r_229__14_,r_229__13_,r_229__12_,r_229__11_,r_229__10_,
  r_229__9_,r_229__8_,r_229__7_,r_229__6_,r_229__5_,r_229__4_,r_229__3_,r_229__2_,
  r_229__1_,r_229__0_,r_230__63_,r_230__62_,r_230__61_,r_230__60_,r_230__59_,r_230__58_,
  r_230__57_,r_230__56_,r_230__55_,r_230__54_,r_230__53_,r_230__52_,r_230__51_,
  r_230__50_,r_230__49_,r_230__48_,r_230__47_,r_230__46_,r_230__45_,r_230__44_,
  r_230__43_,r_230__42_,r_230__41_,r_230__40_,r_230__39_,r_230__38_,r_230__37_,
  r_230__36_,r_230__35_,r_230__34_,r_230__33_,r_230__32_,r_230__31_,r_230__30_,r_230__29_,
  r_230__28_,r_230__27_,r_230__26_,r_230__25_,r_230__24_,r_230__23_,r_230__22_,
  r_230__21_,r_230__20_,r_230__19_,r_230__18_,r_230__17_,r_230__16_,r_230__15_,
  r_230__14_,r_230__13_,r_230__12_,r_230__11_,r_230__10_,r_230__9_,r_230__8_,r_230__7_,
  r_230__6_,r_230__5_,r_230__4_,r_230__3_,r_230__2_,r_230__1_,r_230__0_,r_231__63_,
  r_231__62_,r_231__61_,r_231__60_,r_231__59_,r_231__58_,r_231__57_,r_231__56_,
  r_231__55_,r_231__54_,r_231__53_,r_231__52_,r_231__51_,r_231__50_,r_231__49_,
  r_231__48_,r_231__47_,r_231__46_,r_231__45_,r_231__44_,r_231__43_,r_231__42_,
  r_231__41_,r_231__40_,r_231__39_,r_231__38_,r_231__37_,r_231__36_,r_231__35_,r_231__34_,
  r_231__33_,r_231__32_,r_231__31_,r_231__30_,r_231__29_,r_231__28_,r_231__27_,
  r_231__26_,r_231__25_,r_231__24_,r_231__23_,r_231__22_,r_231__21_,r_231__20_,
  r_231__19_,r_231__18_,r_231__17_,r_231__16_,r_231__15_,r_231__14_,r_231__13_,r_231__12_,
  r_231__11_,r_231__10_,r_231__9_,r_231__8_,r_231__7_,r_231__6_,r_231__5_,
  r_231__4_,r_231__3_,r_231__2_,r_231__1_,r_231__0_,r_232__63_,r_232__62_,r_232__61_,
  r_232__60_,r_232__59_,r_232__58_,r_232__57_,r_232__56_,r_232__55_,r_232__54_,
  r_232__53_,r_232__52_,r_232__51_,r_232__50_,r_232__49_,r_232__48_,r_232__47_,r_232__46_,
  r_232__45_,r_232__44_,r_232__43_,r_232__42_,r_232__41_,r_232__40_,r_232__39_,
  r_232__38_,r_232__37_,r_232__36_,r_232__35_,r_232__34_,r_232__33_,r_232__32_,
  r_232__31_,r_232__30_,r_232__29_,r_232__28_,r_232__27_,r_232__26_,r_232__25_,
  r_232__24_,r_232__23_,r_232__22_,r_232__21_,r_232__20_,r_232__19_,r_232__18_,r_232__17_,
  r_232__16_,r_232__15_,r_232__14_,r_232__13_,r_232__12_,r_232__11_,r_232__10_,
  r_232__9_,r_232__8_,r_232__7_,r_232__6_,r_232__5_,r_232__4_,r_232__3_,r_232__2_,
  r_232__1_,r_232__0_,r_233__63_,r_233__62_,r_233__61_,r_233__60_,r_233__59_,
  r_233__58_,r_233__57_,r_233__56_,r_233__55_,r_233__54_,r_233__53_,r_233__52_,r_233__51_,
  r_233__50_,r_233__49_,r_233__48_,r_233__47_,r_233__46_,r_233__45_,r_233__44_,
  r_233__43_,r_233__42_,r_233__41_,r_233__40_,r_233__39_,r_233__38_,r_233__37_,
  r_233__36_,r_233__35_,r_233__34_,r_233__33_,r_233__32_,r_233__31_,r_233__30_,
  r_233__29_,r_233__28_,r_233__27_,r_233__26_,r_233__25_,r_233__24_,r_233__23_,r_233__22_,
  r_233__21_,r_233__20_,r_233__19_,r_233__18_,r_233__17_,r_233__16_,r_233__15_,
  r_233__14_,r_233__13_,r_233__12_,r_233__11_,r_233__10_,r_233__9_,r_233__8_,r_233__7_,
  r_233__6_,r_233__5_,r_233__4_,r_233__3_,r_233__2_,r_233__1_,r_233__0_,
  r_234__63_,r_234__62_,r_234__61_,r_234__60_,r_234__59_,r_234__58_,r_234__57_,r_234__56_,
  r_234__55_,r_234__54_,r_234__53_,r_234__52_,r_234__51_,r_234__50_,r_234__49_,
  r_234__48_,r_234__47_,r_234__46_,r_234__45_,r_234__44_,r_234__43_,r_234__42_,
  r_234__41_,r_234__40_,r_234__39_,r_234__38_,r_234__37_,r_234__36_,r_234__35_,r_234__34_,
  r_234__33_,r_234__32_,r_234__31_,r_234__30_,r_234__29_,r_234__28_,r_234__27_,
  r_234__26_,r_234__25_,r_234__24_,r_234__23_,r_234__22_,r_234__21_,r_234__20_,
  r_234__19_,r_234__18_,r_234__17_,r_234__16_,r_234__15_,r_234__14_,r_234__13_,
  r_234__12_,r_234__11_,r_234__10_,r_234__9_,r_234__8_,r_234__7_,r_234__6_,r_234__5_,
  r_234__4_,r_234__3_,r_234__2_,r_234__1_,r_234__0_,r_235__63_,r_235__62_,r_235__61_,
  r_235__60_,r_235__59_,r_235__58_,r_235__57_,r_235__56_,r_235__55_,r_235__54_,
  r_235__53_,r_235__52_,r_235__51_,r_235__50_,r_235__49_,r_235__48_,r_235__47_,
  r_235__46_,r_235__45_,r_235__44_,r_235__43_,r_235__42_,r_235__41_,r_235__40_,r_235__39_,
  r_235__38_,r_235__37_,r_235__36_,r_235__35_,r_235__34_,r_235__33_,r_235__32_,
  r_235__31_,r_235__30_,r_235__29_,r_235__28_,r_235__27_,r_235__26_,r_235__25_,
  r_235__24_,r_235__23_,r_235__22_,r_235__21_,r_235__20_,r_235__19_,r_235__18_,
  r_235__17_,r_235__16_,r_235__15_,r_235__14_,r_235__13_,r_235__12_,r_235__11_,r_235__10_,
  r_235__9_,r_235__8_,r_235__7_,r_235__6_,r_235__5_,r_235__4_,r_235__3_,r_235__2_,
  r_235__1_,r_235__0_,r_236__63_,r_236__62_,r_236__61_,r_236__60_,r_236__59_,
  r_236__58_,r_236__57_,r_236__56_,r_236__55_,r_236__54_,r_236__53_,r_236__52_,
  r_236__51_,r_236__50_,r_236__49_,r_236__48_,r_236__47_,r_236__46_,r_236__45_,r_236__44_,
  r_236__43_,r_236__42_,r_236__41_,r_236__40_,r_236__39_,r_236__38_,r_236__37_,
  r_236__36_,r_236__35_,r_236__34_,r_236__33_,r_236__32_,r_236__31_,r_236__30_,
  r_236__29_,r_236__28_,r_236__27_,r_236__26_,r_236__25_,r_236__24_,r_236__23_,r_236__22_,
  r_236__21_,r_236__20_,r_236__19_,r_236__18_,r_236__17_,r_236__16_,r_236__15_,
  r_236__14_,r_236__13_,r_236__12_,r_236__11_,r_236__10_,r_236__9_,r_236__8_,
  r_236__7_,r_236__6_,r_236__5_,r_236__4_,r_236__3_,r_236__2_,r_236__1_,r_236__0_,
  r_237__63_,r_237__62_,r_237__61_,r_237__60_,r_237__59_,r_237__58_,r_237__57_,r_237__56_,
  r_237__55_,r_237__54_,r_237__53_,r_237__52_,r_237__51_,r_237__50_,r_237__49_,
  r_237__48_,r_237__47_,r_237__46_,r_237__45_,r_237__44_,r_237__43_,r_237__42_,
  r_237__41_,r_237__40_,r_237__39_,r_237__38_,r_237__37_,r_237__36_,r_237__35_,
  r_237__34_,r_237__33_,r_237__32_,r_237__31_,r_237__30_,r_237__29_,r_237__28_,r_237__27_,
  r_237__26_,r_237__25_,r_237__24_,r_237__23_,r_237__22_,r_237__21_,r_237__20_,
  r_237__19_,r_237__18_,r_237__17_,r_237__16_,r_237__15_,r_237__14_,r_237__13_,
  r_237__12_,r_237__11_,r_237__10_,r_237__9_,r_237__8_,r_237__7_,r_237__6_,r_237__5_,
  r_237__4_,r_237__3_,r_237__2_,r_237__1_,r_237__0_,r_238__63_,r_238__62_,r_238__61_,
  r_238__60_,r_238__59_,r_238__58_,r_238__57_,r_238__56_,r_238__55_,r_238__54_,
  r_238__53_,r_238__52_,r_238__51_,r_238__50_,r_238__49_,r_238__48_,r_238__47_,
  r_238__46_,r_238__45_,r_238__44_,r_238__43_,r_238__42_,r_238__41_,r_238__40_,
  r_238__39_,r_238__38_,r_238__37_,r_238__36_,r_238__35_,r_238__34_,r_238__33_,r_238__32_,
  r_238__31_,r_238__30_,r_238__29_,r_238__28_,r_238__27_,r_238__26_,r_238__25_,
  r_238__24_,r_238__23_,r_238__22_,r_238__21_,r_238__20_,r_238__19_,r_238__18_,
  r_238__17_,r_238__16_,r_238__15_,r_238__14_,r_238__13_,r_238__12_,r_238__11_,r_238__10_,
  r_238__9_,r_238__8_,r_238__7_,r_238__6_,r_238__5_,r_238__4_,r_238__3_,r_238__2_,
  r_238__1_,r_238__0_,r_239__63_,r_239__62_,r_239__61_,r_239__60_,r_239__59_,
  r_239__58_,r_239__57_,r_239__56_,r_239__55_,r_239__54_,r_239__53_,r_239__52_,
  r_239__51_,r_239__50_,r_239__49_,r_239__48_,r_239__47_,r_239__46_,r_239__45_,r_239__44_,
  r_239__43_,r_239__42_,r_239__41_,r_239__40_,r_239__39_,r_239__38_,r_239__37_,
  r_239__36_,r_239__35_,r_239__34_,r_239__33_,r_239__32_,r_239__31_,r_239__30_,
  r_239__29_,r_239__28_,r_239__27_,r_239__26_,r_239__25_,r_239__24_,r_239__23_,
  r_239__22_,r_239__21_,r_239__20_,r_239__19_,r_239__18_,r_239__17_,r_239__16_,r_239__15_,
  r_239__14_,r_239__13_,r_239__12_,r_239__11_,r_239__10_,r_239__9_,r_239__8_,
  r_239__7_,r_239__6_,r_239__5_,r_239__4_,r_239__3_,r_239__2_,r_239__1_,r_239__0_,
  r_240__63_,r_240__62_,r_240__61_,r_240__60_,r_240__59_,r_240__58_,r_240__57_,
  r_240__56_,r_240__55_,r_240__54_,r_240__53_,r_240__52_,r_240__51_,r_240__50_,r_240__49_,
  r_240__48_,r_240__47_,r_240__46_,r_240__45_,r_240__44_,r_240__43_,r_240__42_,
  r_240__41_,r_240__40_,r_240__39_,r_240__38_,r_240__37_,r_240__36_,r_240__35_,
  r_240__34_,r_240__33_,r_240__32_,r_240__31_,r_240__30_,r_240__29_,r_240__28_,
  r_240__27_,r_240__26_,r_240__25_,r_240__24_,r_240__23_,r_240__22_,r_240__21_,r_240__20_,
  r_240__19_,r_240__18_,r_240__17_,r_240__16_,r_240__15_,r_240__14_,r_240__13_,
  r_240__12_,r_240__11_,r_240__10_,r_240__9_,r_240__8_,r_240__7_,r_240__6_,r_240__5_,
  r_240__4_,r_240__3_,r_240__2_,r_240__1_,r_240__0_,r_241__63_,r_241__62_,
  r_241__61_,r_241__60_,r_241__59_,r_241__58_,r_241__57_,r_241__56_,r_241__55_,r_241__54_,
  r_241__53_,r_241__52_,r_241__51_,r_241__50_,r_241__49_,r_241__48_,r_241__47_,
  r_241__46_,r_241__45_,r_241__44_,r_241__43_,r_241__42_,r_241__41_,r_241__40_,
  r_241__39_,r_241__38_,r_241__37_,r_241__36_,r_241__35_,r_241__34_,r_241__33_,r_241__32_,
  r_241__31_,r_241__30_,r_241__29_,r_241__28_,r_241__27_,r_241__26_,r_241__25_,
  r_241__24_,r_241__23_,r_241__22_,r_241__21_,r_241__20_,r_241__19_,r_241__18_,
  r_241__17_,r_241__16_,r_241__15_,r_241__14_,r_241__13_,r_241__12_,r_241__11_,
  r_241__10_,r_241__9_,r_241__8_,r_241__7_,r_241__6_,r_241__5_,r_241__4_,r_241__3_,
  r_241__2_,r_241__1_,r_241__0_,r_242__63_,r_242__62_,r_242__61_,r_242__60_,r_242__59_,
  r_242__58_,r_242__57_,r_242__56_,r_242__55_,r_242__54_,r_242__53_,r_242__52_,
  r_242__51_,r_242__50_,r_242__49_,r_242__48_,r_242__47_,r_242__46_,r_242__45_,
  r_242__44_,r_242__43_,r_242__42_,r_242__41_,r_242__40_,r_242__39_,r_242__38_,r_242__37_,
  r_242__36_,r_242__35_,r_242__34_,r_242__33_,r_242__32_,r_242__31_,r_242__30_,
  r_242__29_,r_242__28_,r_242__27_,r_242__26_,r_242__25_,r_242__24_,r_242__23_,
  r_242__22_,r_242__21_,r_242__20_,r_242__19_,r_242__18_,r_242__17_,r_242__16_,
  r_242__15_,r_242__14_,r_242__13_,r_242__12_,r_242__11_,r_242__10_,r_242__9_,r_242__8_,
  r_242__7_,r_242__6_,r_242__5_,r_242__4_,r_242__3_,r_242__2_,r_242__1_,r_242__0_,
  r_243__63_,r_243__62_,r_243__61_,r_243__60_,r_243__59_,r_243__58_,r_243__57_,
  r_243__56_,r_243__55_,r_243__54_,r_243__53_,r_243__52_,r_243__51_,r_243__50_,
  r_243__49_,r_243__48_,r_243__47_,r_243__46_,r_243__45_,r_243__44_,r_243__43_,r_243__42_,
  r_243__41_,r_243__40_,r_243__39_,r_243__38_,r_243__37_,r_243__36_,r_243__35_,
  r_243__34_,r_243__33_,r_243__32_,r_243__31_,r_243__30_,r_243__29_,r_243__28_,
  r_243__27_,r_243__26_,r_243__25_,r_243__24_,r_243__23_,r_243__22_,r_243__21_,r_243__20_,
  r_243__19_,r_243__18_,r_243__17_,r_243__16_,r_243__15_,r_243__14_,r_243__13_,
  r_243__12_,r_243__11_,r_243__10_,r_243__9_,r_243__8_,r_243__7_,r_243__6_,r_243__5_,
  r_243__4_,r_243__3_,r_243__2_,r_243__1_,r_243__0_,r_244__63_,r_244__62_,
  r_244__61_,r_244__60_,r_244__59_,r_244__58_,r_244__57_,r_244__56_,r_244__55_,r_244__54_,
  r_244__53_,r_244__52_,r_244__51_,r_244__50_,r_244__49_,r_244__48_,r_244__47_,
  r_244__46_,r_244__45_,r_244__44_,r_244__43_,r_244__42_,r_244__41_,r_244__40_,
  r_244__39_,r_244__38_,r_244__37_,r_244__36_,r_244__35_,r_244__34_,r_244__33_,
  r_244__32_,r_244__31_,r_244__30_,r_244__29_,r_244__28_,r_244__27_,r_244__26_,r_244__25_,
  r_244__24_,r_244__23_,r_244__22_,r_244__21_,r_244__20_,r_244__19_,r_244__18_,
  r_244__17_,r_244__16_,r_244__15_,r_244__14_,r_244__13_,r_244__12_,r_244__11_,
  r_244__10_,r_244__9_,r_244__8_,r_244__7_,r_244__6_,r_244__5_,r_244__4_,r_244__3_,
  r_244__2_,r_244__1_,r_244__0_,r_245__63_,r_245__62_,r_245__61_,r_245__60_,r_245__59_,
  r_245__58_,r_245__57_,r_245__56_,r_245__55_,r_245__54_,r_245__53_,r_245__52_,
  r_245__51_,r_245__50_,r_245__49_,r_245__48_,r_245__47_,r_245__46_,r_245__45_,
  r_245__44_,r_245__43_,r_245__42_,r_245__41_,r_245__40_,r_245__39_,r_245__38_,
  r_245__37_,r_245__36_,r_245__35_,r_245__34_,r_245__33_,r_245__32_,r_245__31_,r_245__30_,
  r_245__29_,r_245__28_,r_245__27_,r_245__26_,r_245__25_,r_245__24_,r_245__23_,
  r_245__22_,r_245__21_,r_245__20_,r_245__19_,r_245__18_,r_245__17_,r_245__16_,
  r_245__15_,r_245__14_,r_245__13_,r_245__12_,r_245__11_,r_245__10_,r_245__9_,r_245__8_,
  r_245__7_,r_245__6_,r_245__5_,r_245__4_,r_245__3_,r_245__2_,r_245__1_,r_245__0_,
  r_246__63_,r_246__62_,r_246__61_,r_246__60_,r_246__59_,r_246__58_,r_246__57_,
  r_246__56_,r_246__55_,r_246__54_,r_246__53_,r_246__52_,r_246__51_,r_246__50_,
  r_246__49_,r_246__48_,r_246__47_,r_246__46_,r_246__45_,r_246__44_,r_246__43_,r_246__42_,
  r_246__41_,r_246__40_,r_246__39_,r_246__38_,r_246__37_,r_246__36_,r_246__35_,
  r_246__34_,r_246__33_,r_246__32_,r_246__31_,r_246__30_,r_246__29_,r_246__28_,
  r_246__27_,r_246__26_,r_246__25_,r_246__24_,r_246__23_,r_246__22_,r_246__21_,
  r_246__20_,r_246__19_,r_246__18_,r_246__17_,r_246__16_,r_246__15_,r_246__14_,r_246__13_,
  r_246__12_,r_246__11_,r_246__10_,r_246__9_,r_246__8_,r_246__7_,r_246__6_,
  r_246__5_,r_246__4_,r_246__3_,r_246__2_,r_246__1_,r_246__0_,r_247__63_,r_247__62_,
  r_247__61_,r_247__60_,r_247__59_,r_247__58_,r_247__57_,r_247__56_,r_247__55_,
  r_247__54_,r_247__53_,r_247__52_,r_247__51_,r_247__50_,r_247__49_,r_247__48_,r_247__47_,
  r_247__46_,r_247__45_,r_247__44_,r_247__43_,r_247__42_,r_247__41_,r_247__40_,
  r_247__39_,r_247__38_,r_247__37_,r_247__36_,r_247__35_,r_247__34_,r_247__33_,
  r_247__32_,r_247__31_,r_247__30_,r_247__29_,r_247__28_,r_247__27_,r_247__26_,
  r_247__25_,r_247__24_,r_247__23_,r_247__22_,r_247__21_,r_247__20_,r_247__19_,r_247__18_,
  r_247__17_,r_247__16_,r_247__15_,r_247__14_,r_247__13_,r_247__12_,r_247__11_,
  r_247__10_,r_247__9_,r_247__8_,r_247__7_,r_247__6_,r_247__5_,r_247__4_,r_247__3_,
  r_247__2_,r_247__1_,r_247__0_,r_248__63_,r_248__62_,r_248__61_,r_248__60_,
  r_248__59_,r_248__58_,r_248__57_,r_248__56_,r_248__55_,r_248__54_,r_248__53_,r_248__52_,
  r_248__51_,r_248__50_,r_248__49_,r_248__48_,r_248__47_,r_248__46_,r_248__45_,
  r_248__44_,r_248__43_,r_248__42_,r_248__41_,r_248__40_,r_248__39_,r_248__38_,
  r_248__37_,r_248__36_,r_248__35_,r_248__34_,r_248__33_,r_248__32_,r_248__31_,r_248__30_,
  r_248__29_,r_248__28_,r_248__27_,r_248__26_,r_248__25_,r_248__24_,r_248__23_,
  r_248__22_,r_248__21_,r_248__20_,r_248__19_,r_248__18_,r_248__17_,r_248__16_,
  r_248__15_,r_248__14_,r_248__13_,r_248__12_,r_248__11_,r_248__10_,r_248__9_,r_248__8_,
  r_248__7_,r_248__6_,r_248__5_,r_248__4_,r_248__3_,r_248__2_,r_248__1_,r_248__0_,
  r_249__63_,r_249__62_,r_249__61_,r_249__60_,r_249__59_,r_249__58_,r_249__57_,
  r_249__56_,r_249__55_,r_249__54_,r_249__53_,r_249__52_,r_249__51_,r_249__50_,
  r_249__49_,r_249__48_,r_249__47_,r_249__46_,r_249__45_,r_249__44_,r_249__43_,
  r_249__42_,r_249__41_,r_249__40_,r_249__39_,r_249__38_,r_249__37_,r_249__36_,r_249__35_,
  r_249__34_,r_249__33_,r_249__32_,r_249__31_,r_249__30_,r_249__29_,r_249__28_,
  r_249__27_,r_249__26_,r_249__25_,r_249__24_,r_249__23_,r_249__22_,r_249__21_,
  r_249__20_,r_249__19_,r_249__18_,r_249__17_,r_249__16_,r_249__15_,r_249__14_,
  r_249__13_,r_249__12_,r_249__11_,r_249__10_,r_249__9_,r_249__8_,r_249__7_,r_249__6_,
  r_249__5_,r_249__4_,r_249__3_,r_249__2_,r_249__1_,r_249__0_,r_250__63_,r_250__62_,
  r_250__61_,r_250__60_,r_250__59_,r_250__58_,r_250__57_,r_250__56_,r_250__55_,
  r_250__54_,r_250__53_,r_250__52_,r_250__51_,r_250__50_,r_250__49_,r_250__48_,
  r_250__47_,r_250__46_,r_250__45_,r_250__44_,r_250__43_,r_250__42_,r_250__41_,r_250__40_,
  r_250__39_,r_250__38_,r_250__37_,r_250__36_,r_250__35_,r_250__34_,r_250__33_,
  r_250__32_,r_250__31_,r_250__30_,r_250__29_,r_250__28_,r_250__27_,r_250__26_,
  r_250__25_,r_250__24_,r_250__23_,r_250__22_,r_250__21_,r_250__20_,r_250__19_,r_250__18_,
  r_250__17_,r_250__16_,r_250__15_,r_250__14_,r_250__13_,r_250__12_,r_250__11_,
  r_250__10_,r_250__9_,r_250__8_,r_250__7_,r_250__6_,r_250__5_,r_250__4_,r_250__3_,
  r_250__2_,r_250__1_,r_250__0_,r_251__63_,r_251__62_,r_251__61_,r_251__60_,
  r_251__59_,r_251__58_,r_251__57_,r_251__56_,r_251__55_,r_251__54_,r_251__53_,r_251__52_,
  r_251__51_,r_251__50_,r_251__49_,r_251__48_,r_251__47_,r_251__46_,r_251__45_,
  r_251__44_,r_251__43_,r_251__42_,r_251__41_,r_251__40_,r_251__39_,r_251__38_,
  r_251__37_,r_251__36_,r_251__35_,r_251__34_,r_251__33_,r_251__32_,r_251__31_,
  r_251__30_,r_251__29_,r_251__28_,r_251__27_,r_251__26_,r_251__25_,r_251__24_,r_251__23_,
  r_251__22_,r_251__21_,r_251__20_,r_251__19_,r_251__18_,r_251__17_,r_251__16_,
  r_251__15_,r_251__14_,r_251__13_,r_251__12_,r_251__11_,r_251__10_,r_251__9_,
  r_251__8_,r_251__7_,r_251__6_,r_251__5_,r_251__4_,r_251__3_,r_251__2_,r_251__1_,
  r_251__0_,r_252__63_,r_252__62_,r_252__61_,r_252__60_,r_252__59_,r_252__58_,r_252__57_,
  r_252__56_,r_252__55_,r_252__54_,r_252__53_,r_252__52_,r_252__51_,r_252__50_,
  r_252__49_,r_252__48_,r_252__47_,r_252__46_,r_252__45_,r_252__44_,r_252__43_,
  r_252__42_,r_252__41_,r_252__40_,r_252__39_,r_252__38_,r_252__37_,r_252__36_,
  r_252__35_,r_252__34_,r_252__33_,r_252__32_,r_252__31_,r_252__30_,r_252__29_,r_252__28_,
  r_252__27_,r_252__26_,r_252__25_,r_252__24_,r_252__23_,r_252__22_,r_252__21_,
  r_252__20_,r_252__19_,r_252__18_,r_252__17_,r_252__16_,r_252__15_,r_252__14_,
  r_252__13_,r_252__12_,r_252__11_,r_252__10_,r_252__9_,r_252__8_,r_252__7_,r_252__6_,
  r_252__5_,r_252__4_,r_252__3_,r_252__2_,r_252__1_,r_252__0_,r_253__63_,r_253__62_,
  r_253__61_,r_253__60_,r_253__59_,r_253__58_,r_253__57_,r_253__56_,r_253__55_,
  r_253__54_,r_253__53_,r_253__52_,r_253__51_,r_253__50_,r_253__49_,r_253__48_,
  r_253__47_,r_253__46_,r_253__45_,r_253__44_,r_253__43_,r_253__42_,r_253__41_,r_253__40_,
  r_253__39_,r_253__38_,r_253__37_,r_253__36_,r_253__35_,r_253__34_,r_253__33_,
  r_253__32_,r_253__31_,r_253__30_,r_253__29_,r_253__28_,r_253__27_,r_253__26_,
  r_253__25_,r_253__24_,r_253__23_,r_253__22_,r_253__21_,r_253__20_,r_253__19_,
  r_253__18_,r_253__17_,r_253__16_,r_253__15_,r_253__14_,r_253__13_,r_253__12_,r_253__11_,
  r_253__10_,r_253__9_,r_253__8_,r_253__7_,r_253__6_,r_253__5_,r_253__4_,r_253__3_,
  r_253__2_,r_253__1_,r_253__0_,r_254__63_,r_254__62_,r_254__61_,r_254__60_,
  r_254__59_,r_254__58_,r_254__57_,r_254__56_,r_254__55_,r_254__54_,r_254__53_,
  r_254__52_,r_254__51_,r_254__50_,r_254__49_,r_254__48_,r_254__47_,r_254__46_,r_254__45_,
  r_254__44_,r_254__43_,r_254__42_,r_254__41_,r_254__40_,r_254__39_,r_254__38_,
  r_254__37_,r_254__36_,r_254__35_,r_254__34_,r_254__33_,r_254__32_,r_254__31_,
  r_254__30_,r_254__29_,r_254__28_,r_254__27_,r_254__26_,r_254__25_,r_254__24_,
  r_254__23_,r_254__22_,r_254__21_,r_254__20_,r_254__19_,r_254__18_,r_254__17_,r_254__16_,
  r_254__15_,r_254__14_,r_254__13_,r_254__12_,r_254__11_,r_254__10_,r_254__9_,
  r_254__8_,r_254__7_,r_254__6_,r_254__5_,r_254__4_,r_254__3_,r_254__2_,r_254__1_,
  r_254__0_,r_255__63_,r_255__62_,r_255__61_,r_255__60_,r_255__59_,r_255__58_,
  r_255__57_,r_255__56_,r_255__55_,r_255__54_,r_255__53_,r_255__52_,r_255__51_,r_255__50_,
  r_255__49_,r_255__48_,r_255__47_,r_255__46_,r_255__45_,r_255__44_,r_255__43_,
  r_255__42_,r_255__41_,r_255__40_,r_255__39_,r_255__38_,r_255__37_,r_255__36_,
  r_255__35_,r_255__34_,r_255__33_,r_255__32_,r_255__31_,r_255__30_,r_255__29_,r_255__28_,
  r_255__27_,r_255__26_,r_255__25_,r_255__24_,r_255__23_,r_255__22_,r_255__21_,
  r_255__20_,r_255__19_,r_255__18_,r_255__17_,r_255__16_,r_255__15_,r_255__14_,
  r_255__13_,r_255__12_,r_255__11_,r_255__10_,r_255__9_,r_255__8_,r_255__7_,r_255__6_,
  r_255__5_,r_255__4_,r_255__3_,r_255__2_,r_255__1_,r_255__0_,r_256__63_,r_256__62_,
  r_256__61_,r_256__60_,r_256__59_,r_256__58_,r_256__57_,r_256__56_,r_256__55_,
  r_256__54_,r_256__53_,r_256__52_,r_256__51_,r_256__50_,r_256__49_,r_256__48_,
  r_256__47_,r_256__46_,r_256__45_,r_256__44_,r_256__43_,r_256__42_,r_256__41_,
  r_256__40_,r_256__39_,r_256__38_,r_256__37_,r_256__36_,r_256__35_,r_256__34_,r_256__33_,
  r_256__32_,r_256__31_,r_256__30_,r_256__29_,r_256__28_,r_256__27_,r_256__26_,
  r_256__25_,r_256__24_,r_256__23_,r_256__22_,r_256__21_,r_256__20_,r_256__19_,
  r_256__18_,r_256__17_,r_256__16_,r_256__15_,r_256__14_,r_256__13_,r_256__12_,
  r_256__11_,r_256__10_,r_256__9_,r_256__8_,r_256__7_,r_256__6_,r_256__5_,r_256__4_,
  r_256__3_,r_256__2_,r_256__1_,r_256__0_,r_257__63_,r_257__62_,r_257__61_,r_257__60_,
  r_257__59_,r_257__58_,r_257__57_,r_257__56_,r_257__55_,r_257__54_,r_257__53_,
  r_257__52_,r_257__51_,r_257__50_,r_257__49_,r_257__48_,r_257__47_,r_257__46_,
  r_257__45_,r_257__44_,r_257__43_,r_257__42_,r_257__41_,r_257__40_,r_257__39_,r_257__38_,
  r_257__37_,r_257__36_,r_257__35_,r_257__34_,r_257__33_,r_257__32_,r_257__31_,
  r_257__30_,r_257__29_,r_257__28_,r_257__27_,r_257__26_,r_257__25_,r_257__24_,
  r_257__23_,r_257__22_,r_257__21_,r_257__20_,r_257__19_,r_257__18_,r_257__17_,r_257__16_,
  r_257__15_,r_257__14_,r_257__13_,r_257__12_,r_257__11_,r_257__10_,r_257__9_,
  r_257__8_,r_257__7_,r_257__6_,r_257__5_,r_257__4_,r_257__3_,r_257__2_,r_257__1_,
  r_257__0_,r_258__63_,r_258__62_,r_258__61_,r_258__60_,r_258__59_,r_258__58_,
  r_258__57_,r_258__56_,r_258__55_,r_258__54_,r_258__53_,r_258__52_,r_258__51_,r_258__50_,
  r_258__49_,r_258__48_,r_258__47_,r_258__46_,r_258__45_,r_258__44_,r_258__43_,
  r_258__42_,r_258__41_,r_258__40_,r_258__39_,r_258__38_,r_258__37_,r_258__36_,
  r_258__35_,r_258__34_,r_258__33_,r_258__32_,r_258__31_,r_258__30_,r_258__29_,
  r_258__28_,r_258__27_,r_258__26_,r_258__25_,r_258__24_,r_258__23_,r_258__22_,r_258__21_,
  r_258__20_,r_258__19_,r_258__18_,r_258__17_,r_258__16_,r_258__15_,r_258__14_,
  r_258__13_,r_258__12_,r_258__11_,r_258__10_,r_258__9_,r_258__8_,r_258__7_,r_258__6_,
  r_258__5_,r_258__4_,r_258__3_,r_258__2_,r_258__1_,r_258__0_,r_259__63_,
  r_259__62_,r_259__61_,r_259__60_,r_259__59_,r_259__58_,r_259__57_,r_259__56_,r_259__55_,
  r_259__54_,r_259__53_,r_259__52_,r_259__51_,r_259__50_,r_259__49_,r_259__48_,
  r_259__47_,r_259__46_,r_259__45_,r_259__44_,r_259__43_,r_259__42_,r_259__41_,
  r_259__40_,r_259__39_,r_259__38_,r_259__37_,r_259__36_,r_259__35_,r_259__34_,
  r_259__33_,r_259__32_,r_259__31_,r_259__30_,r_259__29_,r_259__28_,r_259__27_,r_259__26_,
  r_259__25_,r_259__24_,r_259__23_,r_259__22_,r_259__21_,r_259__20_,r_259__19_,
  r_259__18_,r_259__17_,r_259__16_,r_259__15_,r_259__14_,r_259__13_,r_259__12_,
  r_259__11_,r_259__10_,r_259__9_,r_259__8_,r_259__7_,r_259__6_,r_259__5_,r_259__4_,
  r_259__3_,r_259__2_,r_259__1_,r_259__0_,r_260__63_,r_260__62_,r_260__61_,r_260__60_,
  r_260__59_,r_260__58_,r_260__57_,r_260__56_,r_260__55_,r_260__54_,r_260__53_,
  r_260__52_,r_260__51_,r_260__50_,r_260__49_,r_260__48_,r_260__47_,r_260__46_,
  r_260__45_,r_260__44_,r_260__43_,r_260__42_,r_260__41_,r_260__40_,r_260__39_,r_260__38_,
  r_260__37_,r_260__36_,r_260__35_,r_260__34_,r_260__33_,r_260__32_,r_260__31_,
  r_260__30_,r_260__29_,r_260__28_,r_260__27_,r_260__26_,r_260__25_,r_260__24_,
  r_260__23_,r_260__22_,r_260__21_,r_260__20_,r_260__19_,r_260__18_,r_260__17_,
  r_260__16_,r_260__15_,r_260__14_,r_260__13_,r_260__12_,r_260__11_,r_260__10_,r_260__9_,
  r_260__8_,r_260__7_,r_260__6_,r_260__5_,r_260__4_,r_260__3_,r_260__2_,r_260__1_,
  r_260__0_,r_261__63_,r_261__62_,r_261__61_,r_261__60_,r_261__59_,r_261__58_,
  r_261__57_,r_261__56_,r_261__55_,r_261__54_,r_261__53_,r_261__52_,r_261__51_,
  r_261__50_,r_261__49_,r_261__48_,r_261__47_,r_261__46_,r_261__45_,r_261__44_,r_261__43_,
  r_261__42_,r_261__41_,r_261__40_,r_261__39_,r_261__38_,r_261__37_,r_261__36_,
  r_261__35_,r_261__34_,r_261__33_,r_261__32_,r_261__31_,r_261__30_,r_261__29_,
  r_261__28_,r_261__27_,r_261__26_,r_261__25_,r_261__24_,r_261__23_,r_261__22_,
  r_261__21_,r_261__20_,r_261__19_,r_261__18_,r_261__17_,r_261__16_,r_261__15_,r_261__14_,
  r_261__13_,r_261__12_,r_261__11_,r_261__10_,r_261__9_,r_261__8_,r_261__7_,
  r_261__6_,r_261__5_,r_261__4_,r_261__3_,r_261__2_,r_261__1_,r_261__0_,r_262__63_,
  r_262__62_,r_262__61_,r_262__60_,r_262__59_,r_262__58_,r_262__57_,r_262__56_,
  r_262__55_,r_262__54_,r_262__53_,r_262__52_,r_262__51_,r_262__50_,r_262__49_,r_262__48_,
  r_262__47_,r_262__46_,r_262__45_,r_262__44_,r_262__43_,r_262__42_,r_262__41_,
  r_262__40_,r_262__39_,r_262__38_,r_262__37_,r_262__36_,r_262__35_,r_262__34_,
  r_262__33_,r_262__32_,r_262__31_,r_262__30_,r_262__29_,r_262__28_,r_262__27_,r_262__26_,
  r_262__25_,r_262__24_,r_262__23_,r_262__22_,r_262__21_,r_262__20_,r_262__19_,
  r_262__18_,r_262__17_,r_262__16_,r_262__15_,r_262__14_,r_262__13_,r_262__12_,
  r_262__11_,r_262__10_,r_262__9_,r_262__8_,r_262__7_,r_262__6_,r_262__5_,r_262__4_,
  r_262__3_,r_262__2_,r_262__1_,r_262__0_,r_263__63_,r_263__62_,r_263__61_,r_263__60_,
  r_263__59_,r_263__58_,r_263__57_,r_263__56_,r_263__55_,r_263__54_,r_263__53_,
  r_263__52_,r_263__51_,r_263__50_,r_263__49_,r_263__48_,r_263__47_,r_263__46_,
  r_263__45_,r_263__44_,r_263__43_,r_263__42_,r_263__41_,r_263__40_,r_263__39_,
  r_263__38_,r_263__37_,r_263__36_,r_263__35_,r_263__34_,r_263__33_,r_263__32_,r_263__31_,
  r_263__30_,r_263__29_,r_263__28_,r_263__27_,r_263__26_,r_263__25_,r_263__24_,
  r_263__23_,r_263__22_,r_263__21_,r_263__20_,r_263__19_,r_263__18_,r_263__17_,
  r_263__16_,r_263__15_,r_263__14_,r_263__13_,r_263__12_,r_263__11_,r_263__10_,r_263__9_,
  r_263__8_,r_263__7_,r_263__6_,r_263__5_,r_263__4_,r_263__3_,r_263__2_,r_263__1_,
  r_263__0_,r_264__63_,r_264__62_,r_264__61_,r_264__60_,r_264__59_,r_264__58_,
  r_264__57_,r_264__56_,r_264__55_,r_264__54_,r_264__53_,r_264__52_,r_264__51_,
  r_264__50_,r_264__49_,r_264__48_,r_264__47_,r_264__46_,r_264__45_,r_264__44_,
  r_264__43_,r_264__42_,r_264__41_,r_264__40_,r_264__39_,r_264__38_,r_264__37_,r_264__36_,
  r_264__35_,r_264__34_,r_264__33_,r_264__32_,r_264__31_,r_264__30_,r_264__29_,
  r_264__28_,r_264__27_,r_264__26_,r_264__25_,r_264__24_,r_264__23_,r_264__22_,
  r_264__21_,r_264__20_,r_264__19_,r_264__18_,r_264__17_,r_264__16_,r_264__15_,r_264__14_,
  r_264__13_,r_264__12_,r_264__11_,r_264__10_,r_264__9_,r_264__8_,r_264__7_,
  r_264__6_,r_264__5_,r_264__4_,r_264__3_,r_264__2_,r_264__1_,r_264__0_,r_265__63_,
  r_265__62_,r_265__61_,r_265__60_,r_265__59_,r_265__58_,r_265__57_,r_265__56_,
  r_265__55_,r_265__54_,r_265__53_,r_265__52_,r_265__51_,r_265__50_,r_265__49_,r_265__48_,
  r_265__47_,r_265__46_,r_265__45_,r_265__44_,r_265__43_,r_265__42_,r_265__41_,
  r_265__40_,r_265__39_,r_265__38_,r_265__37_,r_265__36_,r_265__35_,r_265__34_,
  r_265__33_,r_265__32_,r_265__31_,r_265__30_,r_265__29_,r_265__28_,r_265__27_,
  r_265__26_,r_265__25_,r_265__24_,r_265__23_,r_265__22_,r_265__21_,r_265__20_,r_265__19_,
  r_265__18_,r_265__17_,r_265__16_,r_265__15_,r_265__14_,r_265__13_,r_265__12_,
  r_265__11_,r_265__10_,r_265__9_,r_265__8_,r_265__7_,r_265__6_,r_265__5_,r_265__4_,
  r_265__3_,r_265__2_,r_265__1_,r_265__0_,r_266__63_,r_266__62_,r_266__61_,
  r_266__60_,r_266__59_,r_266__58_,r_266__57_,r_266__56_,r_266__55_,r_266__54_,r_266__53_,
  r_266__52_,r_266__51_,r_266__50_,r_266__49_,r_266__48_,r_266__47_,r_266__46_,
  r_266__45_,r_266__44_,r_266__43_,r_266__42_,r_266__41_,r_266__40_,r_266__39_,
  r_266__38_,r_266__37_,r_266__36_,r_266__35_,r_266__34_,r_266__33_,r_266__32_,
  r_266__31_,r_266__30_,r_266__29_,r_266__28_,r_266__27_,r_266__26_,r_266__25_,r_266__24_,
  r_266__23_,r_266__22_,r_266__21_,r_266__20_,r_266__19_,r_266__18_,r_266__17_,
  r_266__16_,r_266__15_,r_266__14_,r_266__13_,r_266__12_,r_266__11_,r_266__10_,
  r_266__9_,r_266__8_,r_266__7_,r_266__6_,r_266__5_,r_266__4_,r_266__3_,r_266__2_,
  r_266__1_,r_266__0_,r_267__63_,r_267__62_,r_267__61_,r_267__60_,r_267__59_,r_267__58_,
  r_267__57_,r_267__56_,r_267__55_,r_267__54_,r_267__53_,r_267__52_,r_267__51_,
  r_267__50_,r_267__49_,r_267__48_,r_267__47_,r_267__46_,r_267__45_,r_267__44_,
  r_267__43_,r_267__42_,r_267__41_,r_267__40_,r_267__39_,r_267__38_,r_267__37_,r_267__36_,
  r_267__35_,r_267__34_,r_267__33_,r_267__32_,r_267__31_,r_267__30_,r_267__29_,
  r_267__28_,r_267__27_,r_267__26_,r_267__25_,r_267__24_,r_267__23_,r_267__22_,
  r_267__21_,r_267__20_,r_267__19_,r_267__18_,r_267__17_,r_267__16_,r_267__15_,
  r_267__14_,r_267__13_,r_267__12_,r_267__11_,r_267__10_,r_267__9_,r_267__8_,r_267__7_,
  r_267__6_,r_267__5_,r_267__4_,r_267__3_,r_267__2_,r_267__1_,r_267__0_,r_268__63_,
  r_268__62_,r_268__61_,r_268__60_,r_268__59_,r_268__58_,r_268__57_,r_268__56_,
  r_268__55_,r_268__54_,r_268__53_,r_268__52_,r_268__51_,r_268__50_,r_268__49_,
  r_268__48_,r_268__47_,r_268__46_,r_268__45_,r_268__44_,r_268__43_,r_268__42_,r_268__41_,
  r_268__40_,r_268__39_,r_268__38_,r_268__37_,r_268__36_,r_268__35_,r_268__34_,
  r_268__33_,r_268__32_,r_268__31_,r_268__30_,r_268__29_,r_268__28_,r_268__27_,
  r_268__26_,r_268__25_,r_268__24_,r_268__23_,r_268__22_,r_268__21_,r_268__20_,
  r_268__19_,r_268__18_,r_268__17_,r_268__16_,r_268__15_,r_268__14_,r_268__13_,r_268__12_,
  r_268__11_,r_268__10_,r_268__9_,r_268__8_,r_268__7_,r_268__6_,r_268__5_,r_268__4_,
  r_268__3_,r_268__2_,r_268__1_,r_268__0_,r_269__63_,r_269__62_,r_269__61_,
  r_269__60_,r_269__59_,r_269__58_,r_269__57_,r_269__56_,r_269__55_,r_269__54_,
  r_269__53_,r_269__52_,r_269__51_,r_269__50_,r_269__49_,r_269__48_,r_269__47_,r_269__46_,
  r_269__45_,r_269__44_,r_269__43_,r_269__42_,r_269__41_,r_269__40_,r_269__39_,
  r_269__38_,r_269__37_,r_269__36_,r_269__35_,r_269__34_,r_269__33_,r_269__32_,
  r_269__31_,r_269__30_,r_269__29_,r_269__28_,r_269__27_,r_269__26_,r_269__25_,r_269__24_,
  r_269__23_,r_269__22_,r_269__21_,r_269__20_,r_269__19_,r_269__18_,r_269__17_,
  r_269__16_,r_269__15_,r_269__14_,r_269__13_,r_269__12_,r_269__11_,r_269__10_,
  r_269__9_,r_269__8_,r_269__7_,r_269__6_,r_269__5_,r_269__4_,r_269__3_,r_269__2_,
  r_269__1_,r_269__0_,r_270__63_,r_270__62_,r_270__61_,r_270__60_,r_270__59_,r_270__58_,
  r_270__57_,r_270__56_,r_270__55_,r_270__54_,r_270__53_,r_270__52_,r_270__51_,
  r_270__50_,r_270__49_,r_270__48_,r_270__47_,r_270__46_,r_270__45_,r_270__44_,
  r_270__43_,r_270__42_,r_270__41_,r_270__40_,r_270__39_,r_270__38_,r_270__37_,
  r_270__36_,r_270__35_,r_270__34_,r_270__33_,r_270__32_,r_270__31_,r_270__30_,r_270__29_,
  r_270__28_,r_270__27_,r_270__26_,r_270__25_,r_270__24_,r_270__23_,r_270__22_,
  r_270__21_,r_270__20_,r_270__19_,r_270__18_,r_270__17_,r_270__16_,r_270__15_,
  r_270__14_,r_270__13_,r_270__12_,r_270__11_,r_270__10_,r_270__9_,r_270__8_,r_270__7_,
  r_270__6_,r_270__5_,r_270__4_,r_270__3_,r_270__2_,r_270__1_,r_270__0_,r_271__63_,
  r_271__62_,r_271__61_,r_271__60_,r_271__59_,r_271__58_,r_271__57_,r_271__56_,
  r_271__55_,r_271__54_,r_271__53_,r_271__52_,r_271__51_,r_271__50_,r_271__49_,
  r_271__48_,r_271__47_,r_271__46_,r_271__45_,r_271__44_,r_271__43_,r_271__42_,
  r_271__41_,r_271__40_,r_271__39_,r_271__38_,r_271__37_,r_271__36_,r_271__35_,r_271__34_,
  r_271__33_,r_271__32_,r_271__31_,r_271__30_,r_271__29_,r_271__28_,r_271__27_,
  r_271__26_,r_271__25_,r_271__24_,r_271__23_,r_271__22_,r_271__21_,r_271__20_,
  r_271__19_,r_271__18_,r_271__17_,r_271__16_,r_271__15_,r_271__14_,r_271__13_,r_271__12_,
  r_271__11_,r_271__10_,r_271__9_,r_271__8_,r_271__7_,r_271__6_,r_271__5_,
  r_271__4_,r_271__3_,r_271__2_,r_271__1_,r_271__0_,r_272__63_,r_272__62_,r_272__61_,
  r_272__60_,r_272__59_,r_272__58_,r_272__57_,r_272__56_,r_272__55_,r_272__54_,
  r_272__53_,r_272__52_,r_272__51_,r_272__50_,r_272__49_,r_272__48_,r_272__47_,r_272__46_,
  r_272__45_,r_272__44_,r_272__43_,r_272__42_,r_272__41_,r_272__40_,r_272__39_,
  r_272__38_,r_272__37_,r_272__36_,r_272__35_,r_272__34_,r_272__33_,r_272__32_,
  r_272__31_,r_272__30_,r_272__29_,r_272__28_,r_272__27_,r_272__26_,r_272__25_,
  r_272__24_,r_272__23_,r_272__22_,r_272__21_,r_272__20_,r_272__19_,r_272__18_,r_272__17_,
  r_272__16_,r_272__15_,r_272__14_,r_272__13_,r_272__12_,r_272__11_,r_272__10_,
  r_272__9_,r_272__8_,r_272__7_,r_272__6_,r_272__5_,r_272__4_,r_272__3_,r_272__2_,
  r_272__1_,r_272__0_,r_273__63_,r_273__62_,r_273__61_,r_273__60_,r_273__59_,
  r_273__58_,r_273__57_,r_273__56_,r_273__55_,r_273__54_,r_273__53_,r_273__52_,r_273__51_,
  r_273__50_,r_273__49_,r_273__48_,r_273__47_,r_273__46_,r_273__45_,r_273__44_,
  r_273__43_,r_273__42_,r_273__41_,r_273__40_,r_273__39_,r_273__38_,r_273__37_,
  r_273__36_,r_273__35_,r_273__34_,r_273__33_,r_273__32_,r_273__31_,r_273__30_,
  r_273__29_,r_273__28_,r_273__27_,r_273__26_,r_273__25_,r_273__24_,r_273__23_,r_273__22_,
  r_273__21_,r_273__20_,r_273__19_,r_273__18_,r_273__17_,r_273__16_,r_273__15_,
  r_273__14_,r_273__13_,r_273__12_,r_273__11_,r_273__10_,r_273__9_,r_273__8_,r_273__7_,
  r_273__6_,r_273__5_,r_273__4_,r_273__3_,r_273__2_,r_273__1_,r_273__0_,
  r_274__63_,r_274__62_,r_274__61_,r_274__60_,r_274__59_,r_274__58_,r_274__57_,r_274__56_,
  r_274__55_,r_274__54_,r_274__53_,r_274__52_,r_274__51_,r_274__50_,r_274__49_,
  r_274__48_,r_274__47_,r_274__46_,r_274__45_,r_274__44_,r_274__43_,r_274__42_,
  r_274__41_,r_274__40_,r_274__39_,r_274__38_,r_274__37_,r_274__36_,r_274__35_,r_274__34_,
  r_274__33_,r_274__32_,r_274__31_,r_274__30_,r_274__29_,r_274__28_,r_274__27_,
  r_274__26_,r_274__25_,r_274__24_,r_274__23_,r_274__22_,r_274__21_,r_274__20_,
  r_274__19_,r_274__18_,r_274__17_,r_274__16_,r_274__15_,r_274__14_,r_274__13_,
  r_274__12_,r_274__11_,r_274__10_,r_274__9_,r_274__8_,r_274__7_,r_274__6_,r_274__5_,
  r_274__4_,r_274__3_,r_274__2_,r_274__1_,r_274__0_,r_275__63_,r_275__62_,r_275__61_,
  r_275__60_,r_275__59_,r_275__58_,r_275__57_,r_275__56_,r_275__55_,r_275__54_,
  r_275__53_,r_275__52_,r_275__51_,r_275__50_,r_275__49_,r_275__48_,r_275__47_,
  r_275__46_,r_275__45_,r_275__44_,r_275__43_,r_275__42_,r_275__41_,r_275__40_,r_275__39_,
  r_275__38_,r_275__37_,r_275__36_,r_275__35_,r_275__34_,r_275__33_,r_275__32_,
  r_275__31_,r_275__30_,r_275__29_,r_275__28_,r_275__27_,r_275__26_,r_275__25_,
  r_275__24_,r_275__23_,r_275__22_,r_275__21_,r_275__20_,r_275__19_,r_275__18_,
  r_275__17_,r_275__16_,r_275__15_,r_275__14_,r_275__13_,r_275__12_,r_275__11_,r_275__10_,
  r_275__9_,r_275__8_,r_275__7_,r_275__6_,r_275__5_,r_275__4_,r_275__3_,r_275__2_,
  r_275__1_,r_275__0_,r_276__63_,r_276__62_,r_276__61_,r_276__60_,r_276__59_,
  r_276__58_,r_276__57_,r_276__56_,r_276__55_,r_276__54_,r_276__53_,r_276__52_,
  r_276__51_,r_276__50_,r_276__49_,r_276__48_,r_276__47_,r_276__46_,r_276__45_,r_276__44_,
  r_276__43_,r_276__42_,r_276__41_,r_276__40_,r_276__39_,r_276__38_,r_276__37_,
  r_276__36_,r_276__35_,r_276__34_,r_276__33_,r_276__32_,r_276__31_,r_276__30_,
  r_276__29_,r_276__28_,r_276__27_,r_276__26_,r_276__25_,r_276__24_,r_276__23_,r_276__22_,
  r_276__21_,r_276__20_,r_276__19_,r_276__18_,r_276__17_,r_276__16_,r_276__15_,
  r_276__14_,r_276__13_,r_276__12_,r_276__11_,r_276__10_,r_276__9_,r_276__8_,
  r_276__7_,r_276__6_,r_276__5_,r_276__4_,r_276__3_,r_276__2_,r_276__1_,r_276__0_,
  r_277__63_,r_277__62_,r_277__61_,r_277__60_,r_277__59_,r_277__58_,r_277__57_,r_277__56_,
  r_277__55_,r_277__54_,r_277__53_,r_277__52_,r_277__51_,r_277__50_,r_277__49_,
  r_277__48_,r_277__47_,r_277__46_,r_277__45_,r_277__44_,r_277__43_,r_277__42_,
  r_277__41_,r_277__40_,r_277__39_,r_277__38_,r_277__37_,r_277__36_,r_277__35_,
  r_277__34_,r_277__33_,r_277__32_,r_277__31_,r_277__30_,r_277__29_,r_277__28_,r_277__27_,
  r_277__26_,r_277__25_,r_277__24_,r_277__23_,r_277__22_,r_277__21_,r_277__20_,
  r_277__19_,r_277__18_,r_277__17_,r_277__16_,r_277__15_,r_277__14_,r_277__13_,
  r_277__12_,r_277__11_,r_277__10_,r_277__9_,r_277__8_,r_277__7_,r_277__6_,r_277__5_,
  r_277__4_,r_277__3_,r_277__2_,r_277__1_,r_277__0_,r_278__63_,r_278__62_,r_278__61_,
  r_278__60_,r_278__59_,r_278__58_,r_278__57_,r_278__56_,r_278__55_,r_278__54_,
  r_278__53_,r_278__52_,r_278__51_,r_278__50_,r_278__49_,r_278__48_,r_278__47_,
  r_278__46_,r_278__45_,r_278__44_,r_278__43_,r_278__42_,r_278__41_,r_278__40_,
  r_278__39_,r_278__38_,r_278__37_,r_278__36_,r_278__35_,r_278__34_,r_278__33_,r_278__32_,
  r_278__31_,r_278__30_,r_278__29_,r_278__28_,r_278__27_,r_278__26_,r_278__25_,
  r_278__24_,r_278__23_,r_278__22_,r_278__21_,r_278__20_,r_278__19_,r_278__18_,
  r_278__17_,r_278__16_,r_278__15_,r_278__14_,r_278__13_,r_278__12_,r_278__11_,r_278__10_,
  r_278__9_,r_278__8_,r_278__7_,r_278__6_,r_278__5_,r_278__4_,r_278__3_,r_278__2_,
  r_278__1_,r_278__0_,r_279__63_,r_279__62_,r_279__61_,r_279__60_,r_279__59_,
  r_279__58_,r_279__57_,r_279__56_,r_279__55_,r_279__54_,r_279__53_,r_279__52_,
  r_279__51_,r_279__50_,r_279__49_,r_279__48_,r_279__47_,r_279__46_,r_279__45_,r_279__44_,
  r_279__43_,r_279__42_,r_279__41_,r_279__40_,r_279__39_,r_279__38_,r_279__37_,
  r_279__36_,r_279__35_,r_279__34_,r_279__33_,r_279__32_,r_279__31_,r_279__30_,
  r_279__29_,r_279__28_,r_279__27_,r_279__26_,r_279__25_,r_279__24_,r_279__23_,
  r_279__22_,r_279__21_,r_279__20_,r_279__19_,r_279__18_,r_279__17_,r_279__16_,r_279__15_,
  r_279__14_,r_279__13_,r_279__12_,r_279__11_,r_279__10_,r_279__9_,r_279__8_,
  r_279__7_,r_279__6_,r_279__5_,r_279__4_,r_279__3_,r_279__2_,r_279__1_,r_279__0_,
  r_280__63_,r_280__62_,r_280__61_,r_280__60_,r_280__59_,r_280__58_,r_280__57_,
  r_280__56_,r_280__55_,r_280__54_,r_280__53_,r_280__52_,r_280__51_,r_280__50_,r_280__49_,
  r_280__48_,r_280__47_,r_280__46_,r_280__45_,r_280__44_,r_280__43_,r_280__42_,
  r_280__41_,r_280__40_,r_280__39_,r_280__38_,r_280__37_,r_280__36_,r_280__35_,
  r_280__34_,r_280__33_,r_280__32_,r_280__31_,r_280__30_,r_280__29_,r_280__28_,
  r_280__27_,r_280__26_,r_280__25_,r_280__24_,r_280__23_,r_280__22_,r_280__21_,r_280__20_,
  r_280__19_,r_280__18_,r_280__17_,r_280__16_,r_280__15_,r_280__14_,r_280__13_,
  r_280__12_,r_280__11_,r_280__10_,r_280__9_,r_280__8_,r_280__7_,r_280__6_,r_280__5_,
  r_280__4_,r_280__3_,r_280__2_,r_280__1_,r_280__0_,r_281__63_,r_281__62_,
  r_281__61_,r_281__60_,r_281__59_,r_281__58_,r_281__57_,r_281__56_,r_281__55_,r_281__54_,
  r_281__53_,r_281__52_,r_281__51_,r_281__50_,r_281__49_,r_281__48_,r_281__47_,
  r_281__46_,r_281__45_,r_281__44_,r_281__43_,r_281__42_,r_281__41_,r_281__40_,
  r_281__39_,r_281__38_,r_281__37_,r_281__36_,r_281__35_,r_281__34_,r_281__33_,r_281__32_,
  r_281__31_,r_281__30_,r_281__29_,r_281__28_,r_281__27_,r_281__26_,r_281__25_,
  r_281__24_,r_281__23_,r_281__22_,r_281__21_,r_281__20_,r_281__19_,r_281__18_,
  r_281__17_,r_281__16_,r_281__15_,r_281__14_,r_281__13_,r_281__12_,r_281__11_,
  r_281__10_,r_281__9_,r_281__8_,r_281__7_,r_281__6_,r_281__5_,r_281__4_,r_281__3_,
  r_281__2_,r_281__1_,r_281__0_,r_282__63_,r_282__62_,r_282__61_,r_282__60_,r_282__59_,
  r_282__58_,r_282__57_,r_282__56_,r_282__55_,r_282__54_,r_282__53_,r_282__52_,
  r_282__51_,r_282__50_,r_282__49_,r_282__48_,r_282__47_,r_282__46_,r_282__45_,
  r_282__44_,r_282__43_,r_282__42_,r_282__41_,r_282__40_,r_282__39_,r_282__38_,r_282__37_,
  r_282__36_,r_282__35_,r_282__34_,r_282__33_,r_282__32_,r_282__31_,r_282__30_,
  r_282__29_,r_282__28_,r_282__27_,r_282__26_,r_282__25_,r_282__24_,r_282__23_,
  r_282__22_,r_282__21_,r_282__20_,r_282__19_,r_282__18_,r_282__17_,r_282__16_,
  r_282__15_,r_282__14_,r_282__13_,r_282__12_,r_282__11_,r_282__10_,r_282__9_,r_282__8_,
  r_282__7_,r_282__6_,r_282__5_,r_282__4_,r_282__3_,r_282__2_,r_282__1_,r_282__0_,
  r_283__63_,r_283__62_,r_283__61_,r_283__60_,r_283__59_,r_283__58_,r_283__57_,
  r_283__56_,r_283__55_,r_283__54_,r_283__53_,r_283__52_,r_283__51_,r_283__50_,
  r_283__49_,r_283__48_,r_283__47_,r_283__46_,r_283__45_,r_283__44_,r_283__43_,r_283__42_,
  r_283__41_,r_283__40_,r_283__39_,r_283__38_,r_283__37_,r_283__36_,r_283__35_,
  r_283__34_,r_283__33_,r_283__32_,r_283__31_,r_283__30_,r_283__29_,r_283__28_,
  r_283__27_,r_283__26_,r_283__25_,r_283__24_,r_283__23_,r_283__22_,r_283__21_,r_283__20_,
  r_283__19_,r_283__18_,r_283__17_,r_283__16_,r_283__15_,r_283__14_,r_283__13_,
  r_283__12_,r_283__11_,r_283__10_,r_283__9_,r_283__8_,r_283__7_,r_283__6_,r_283__5_,
  r_283__4_,r_283__3_,r_283__2_,r_283__1_,r_283__0_,r_284__63_,r_284__62_,
  r_284__61_,r_284__60_,r_284__59_,r_284__58_,r_284__57_,r_284__56_,r_284__55_,r_284__54_,
  r_284__53_,r_284__52_,r_284__51_,r_284__50_,r_284__49_,r_284__48_,r_284__47_,
  r_284__46_,r_284__45_,r_284__44_,r_284__43_,r_284__42_,r_284__41_,r_284__40_,
  r_284__39_,r_284__38_,r_284__37_,r_284__36_,r_284__35_,r_284__34_,r_284__33_,
  r_284__32_,r_284__31_,r_284__30_,r_284__29_,r_284__28_,r_284__27_,r_284__26_,r_284__25_,
  r_284__24_,r_284__23_,r_284__22_,r_284__21_,r_284__20_,r_284__19_,r_284__18_,
  r_284__17_,r_284__16_,r_284__15_,r_284__14_,r_284__13_,r_284__12_,r_284__11_,
  r_284__10_,r_284__9_,r_284__8_,r_284__7_,r_284__6_,r_284__5_,r_284__4_,r_284__3_,
  r_284__2_,r_284__1_,r_284__0_,r_285__63_,r_285__62_,r_285__61_,r_285__60_,r_285__59_,
  r_285__58_,r_285__57_,r_285__56_,r_285__55_,r_285__54_,r_285__53_,r_285__52_,
  r_285__51_,r_285__50_,r_285__49_,r_285__48_,r_285__47_,r_285__46_,r_285__45_,
  r_285__44_,r_285__43_,r_285__42_,r_285__41_,r_285__40_,r_285__39_,r_285__38_,
  r_285__37_,r_285__36_,r_285__35_,r_285__34_,r_285__33_,r_285__32_,r_285__31_,r_285__30_,
  r_285__29_,r_285__28_,r_285__27_,r_285__26_,r_285__25_,r_285__24_,r_285__23_,
  r_285__22_,r_285__21_,r_285__20_,r_285__19_,r_285__18_,r_285__17_,r_285__16_,
  r_285__15_,r_285__14_,r_285__13_,r_285__12_,r_285__11_,r_285__10_,r_285__9_,r_285__8_,
  r_285__7_,r_285__6_,r_285__5_,r_285__4_,r_285__3_,r_285__2_,r_285__1_,r_285__0_,
  r_286__63_,r_286__62_,r_286__61_,r_286__60_,r_286__59_,r_286__58_,r_286__57_,
  r_286__56_,r_286__55_,r_286__54_,r_286__53_,r_286__52_,r_286__51_,r_286__50_,
  r_286__49_,r_286__48_,r_286__47_,r_286__46_,r_286__45_,r_286__44_,r_286__43_,r_286__42_,
  r_286__41_,r_286__40_,r_286__39_,r_286__38_,r_286__37_,r_286__36_,r_286__35_,
  r_286__34_,r_286__33_,r_286__32_,r_286__31_,r_286__30_,r_286__29_,r_286__28_,
  r_286__27_,r_286__26_,r_286__25_,r_286__24_,r_286__23_,r_286__22_,r_286__21_,
  r_286__20_,r_286__19_,r_286__18_,r_286__17_,r_286__16_,r_286__15_,r_286__14_,r_286__13_,
  r_286__12_,r_286__11_,r_286__10_,r_286__9_,r_286__8_,r_286__7_,r_286__6_,
  r_286__5_,r_286__4_,r_286__3_,r_286__2_,r_286__1_,r_286__0_,r_287__63_,r_287__62_,
  r_287__61_,r_287__60_,r_287__59_,r_287__58_,r_287__57_,r_287__56_,r_287__55_,
  r_287__54_,r_287__53_,r_287__52_,r_287__51_,r_287__50_,r_287__49_,r_287__48_,r_287__47_,
  r_287__46_,r_287__45_,r_287__44_,r_287__43_,r_287__42_,r_287__41_,r_287__40_,
  r_287__39_,r_287__38_,r_287__37_,r_287__36_,r_287__35_,r_287__34_,r_287__33_,
  r_287__32_,r_287__31_,r_287__30_,r_287__29_,r_287__28_,r_287__27_,r_287__26_,
  r_287__25_,r_287__24_,r_287__23_,r_287__22_,r_287__21_,r_287__20_,r_287__19_,r_287__18_,
  r_287__17_,r_287__16_,r_287__15_,r_287__14_,r_287__13_,r_287__12_,r_287__11_,
  r_287__10_,r_287__9_,r_287__8_,r_287__7_,r_287__6_,r_287__5_,r_287__4_,r_287__3_,
  r_287__2_,r_287__1_,r_287__0_,r_288__63_,r_288__62_,r_288__61_,r_288__60_,
  r_288__59_,r_288__58_,r_288__57_,r_288__56_,r_288__55_,r_288__54_,r_288__53_,r_288__52_,
  r_288__51_,r_288__50_,r_288__49_,r_288__48_,r_288__47_,r_288__46_,r_288__45_,
  r_288__44_,r_288__43_,r_288__42_,r_288__41_,r_288__40_,r_288__39_,r_288__38_,
  r_288__37_,r_288__36_,r_288__35_,r_288__34_,r_288__33_,r_288__32_,r_288__31_,r_288__30_,
  r_288__29_,r_288__28_,r_288__27_,r_288__26_,r_288__25_,r_288__24_,r_288__23_,
  r_288__22_,r_288__21_,r_288__20_,r_288__19_,r_288__18_,r_288__17_,r_288__16_,
  r_288__15_,r_288__14_,r_288__13_,r_288__12_,r_288__11_,r_288__10_,r_288__9_,r_288__8_,
  r_288__7_,r_288__6_,r_288__5_,r_288__4_,r_288__3_,r_288__2_,r_288__1_,r_288__0_,
  r_289__63_,r_289__62_,r_289__61_,r_289__60_,r_289__59_,r_289__58_,r_289__57_,
  r_289__56_,r_289__55_,r_289__54_,r_289__53_,r_289__52_,r_289__51_,r_289__50_,
  r_289__49_,r_289__48_,r_289__47_,r_289__46_,r_289__45_,r_289__44_,r_289__43_,
  r_289__42_,r_289__41_,r_289__40_,r_289__39_,r_289__38_,r_289__37_,r_289__36_,r_289__35_,
  r_289__34_,r_289__33_,r_289__32_,r_289__31_,r_289__30_,r_289__29_,r_289__28_,
  r_289__27_,r_289__26_,r_289__25_,r_289__24_,r_289__23_,r_289__22_,r_289__21_,
  r_289__20_,r_289__19_,r_289__18_,r_289__17_,r_289__16_,r_289__15_,r_289__14_,
  r_289__13_,r_289__12_,r_289__11_,r_289__10_,r_289__9_,r_289__8_,r_289__7_,r_289__6_,
  r_289__5_,r_289__4_,r_289__3_,r_289__2_,r_289__1_,r_289__0_,r_290__63_,r_290__62_,
  r_290__61_,r_290__60_,r_290__59_,r_290__58_,r_290__57_,r_290__56_,r_290__55_,
  r_290__54_,r_290__53_,r_290__52_,r_290__51_,r_290__50_,r_290__49_,r_290__48_,
  r_290__47_,r_290__46_,r_290__45_,r_290__44_,r_290__43_,r_290__42_,r_290__41_,r_290__40_,
  r_290__39_,r_290__38_,r_290__37_,r_290__36_,r_290__35_,r_290__34_,r_290__33_,
  r_290__32_,r_290__31_,r_290__30_,r_290__29_,r_290__28_,r_290__27_,r_290__26_,
  r_290__25_,r_290__24_,r_290__23_,r_290__22_,r_290__21_,r_290__20_,r_290__19_,r_290__18_,
  r_290__17_,r_290__16_,r_290__15_,r_290__14_,r_290__13_,r_290__12_,r_290__11_,
  r_290__10_,r_290__9_,r_290__8_,r_290__7_,r_290__6_,r_290__5_,r_290__4_,r_290__3_,
  r_290__2_,r_290__1_,r_290__0_,r_291__63_,r_291__62_,r_291__61_,r_291__60_,
  r_291__59_,r_291__58_,r_291__57_,r_291__56_,r_291__55_,r_291__54_,r_291__53_,r_291__52_,
  r_291__51_,r_291__50_,r_291__49_,r_291__48_,r_291__47_,r_291__46_,r_291__45_,
  r_291__44_,r_291__43_,r_291__42_,r_291__41_,r_291__40_,r_291__39_,r_291__38_,
  r_291__37_,r_291__36_,r_291__35_,r_291__34_,r_291__33_,r_291__32_,r_291__31_,
  r_291__30_,r_291__29_,r_291__28_,r_291__27_,r_291__26_,r_291__25_,r_291__24_,r_291__23_,
  r_291__22_,r_291__21_,r_291__20_,r_291__19_,r_291__18_,r_291__17_,r_291__16_,
  r_291__15_,r_291__14_,r_291__13_,r_291__12_,r_291__11_,r_291__10_,r_291__9_,
  r_291__8_,r_291__7_,r_291__6_,r_291__5_,r_291__4_,r_291__3_,r_291__2_,r_291__1_,
  r_291__0_,r_292__63_,r_292__62_,r_292__61_,r_292__60_,r_292__59_,r_292__58_,r_292__57_,
  r_292__56_,r_292__55_,r_292__54_,r_292__53_,r_292__52_,r_292__51_,r_292__50_,
  r_292__49_,r_292__48_,r_292__47_,r_292__46_,r_292__45_,r_292__44_,r_292__43_,
  r_292__42_,r_292__41_,r_292__40_,r_292__39_,r_292__38_,r_292__37_,r_292__36_,
  r_292__35_,r_292__34_,r_292__33_,r_292__32_,r_292__31_,r_292__30_,r_292__29_,r_292__28_,
  r_292__27_,r_292__26_,r_292__25_,r_292__24_,r_292__23_,r_292__22_,r_292__21_,
  r_292__20_,r_292__19_,r_292__18_,r_292__17_,r_292__16_,r_292__15_,r_292__14_,
  r_292__13_,r_292__12_,r_292__11_,r_292__10_,r_292__9_,r_292__8_,r_292__7_,r_292__6_,
  r_292__5_,r_292__4_,r_292__3_,r_292__2_,r_292__1_,r_292__0_,r_293__63_,r_293__62_,
  r_293__61_,r_293__60_,r_293__59_,r_293__58_,r_293__57_,r_293__56_,r_293__55_,
  r_293__54_,r_293__53_,r_293__52_,r_293__51_,r_293__50_,r_293__49_,r_293__48_,
  r_293__47_,r_293__46_,r_293__45_,r_293__44_,r_293__43_,r_293__42_,r_293__41_,r_293__40_,
  r_293__39_,r_293__38_,r_293__37_,r_293__36_,r_293__35_,r_293__34_,r_293__33_,
  r_293__32_,r_293__31_,r_293__30_,r_293__29_,r_293__28_,r_293__27_,r_293__26_,
  r_293__25_,r_293__24_,r_293__23_,r_293__22_,r_293__21_,r_293__20_,r_293__19_,
  r_293__18_,r_293__17_,r_293__16_,r_293__15_,r_293__14_,r_293__13_,r_293__12_,r_293__11_,
  r_293__10_,r_293__9_,r_293__8_,r_293__7_,r_293__6_,r_293__5_,r_293__4_,r_293__3_,
  r_293__2_,r_293__1_,r_293__0_,r_294__63_,r_294__62_,r_294__61_,r_294__60_,
  r_294__59_,r_294__58_,r_294__57_,r_294__56_,r_294__55_,r_294__54_,r_294__53_,
  r_294__52_,r_294__51_,r_294__50_,r_294__49_,r_294__48_,r_294__47_,r_294__46_,r_294__45_,
  r_294__44_,r_294__43_,r_294__42_,r_294__41_,r_294__40_,r_294__39_,r_294__38_,
  r_294__37_,r_294__36_,r_294__35_,r_294__34_,r_294__33_,r_294__32_,r_294__31_,
  r_294__30_,r_294__29_,r_294__28_,r_294__27_,r_294__26_,r_294__25_,r_294__24_,
  r_294__23_,r_294__22_,r_294__21_,r_294__20_,r_294__19_,r_294__18_,r_294__17_,r_294__16_,
  r_294__15_,r_294__14_,r_294__13_,r_294__12_,r_294__11_,r_294__10_,r_294__9_,
  r_294__8_,r_294__7_,r_294__6_,r_294__5_,r_294__4_,r_294__3_,r_294__2_,r_294__1_,
  r_294__0_,r_295__63_,r_295__62_,r_295__61_,r_295__60_,r_295__59_,r_295__58_,
  r_295__57_,r_295__56_,r_295__55_,r_295__54_,r_295__53_,r_295__52_,r_295__51_,r_295__50_,
  r_295__49_,r_295__48_,r_295__47_,r_295__46_,r_295__45_,r_295__44_,r_295__43_,
  r_295__42_,r_295__41_,r_295__40_,r_295__39_,r_295__38_,r_295__37_,r_295__36_,
  r_295__35_,r_295__34_,r_295__33_,r_295__32_,r_295__31_,r_295__30_,r_295__29_,r_295__28_,
  r_295__27_,r_295__26_,r_295__25_,r_295__24_,r_295__23_,r_295__22_,r_295__21_,
  r_295__20_,r_295__19_,r_295__18_,r_295__17_,r_295__16_,r_295__15_,r_295__14_,
  r_295__13_,r_295__12_,r_295__11_,r_295__10_,r_295__9_,r_295__8_,r_295__7_,r_295__6_,
  r_295__5_,r_295__4_,r_295__3_,r_295__2_,r_295__1_,r_295__0_,r_296__63_,r_296__62_,
  r_296__61_,r_296__60_,r_296__59_,r_296__58_,r_296__57_,r_296__56_,r_296__55_,
  r_296__54_,r_296__53_,r_296__52_,r_296__51_,r_296__50_,r_296__49_,r_296__48_,
  r_296__47_,r_296__46_,r_296__45_,r_296__44_,r_296__43_,r_296__42_,r_296__41_,
  r_296__40_,r_296__39_,r_296__38_,r_296__37_,r_296__36_,r_296__35_,r_296__34_,r_296__33_,
  r_296__32_,r_296__31_,r_296__30_,r_296__29_,r_296__28_,r_296__27_,r_296__26_,
  r_296__25_,r_296__24_,r_296__23_,r_296__22_,r_296__21_,r_296__20_,r_296__19_,
  r_296__18_,r_296__17_,r_296__16_,r_296__15_,r_296__14_,r_296__13_,r_296__12_,
  r_296__11_,r_296__10_,r_296__9_,r_296__8_,r_296__7_,r_296__6_,r_296__5_,r_296__4_,
  r_296__3_,r_296__2_,r_296__1_,r_296__0_,r_297__63_,r_297__62_,r_297__61_,r_297__60_,
  r_297__59_,r_297__58_,r_297__57_,r_297__56_,r_297__55_,r_297__54_,r_297__53_,
  r_297__52_,r_297__51_,r_297__50_,r_297__49_,r_297__48_,r_297__47_,r_297__46_,
  r_297__45_,r_297__44_,r_297__43_,r_297__42_,r_297__41_,r_297__40_,r_297__39_,r_297__38_,
  r_297__37_,r_297__36_,r_297__35_,r_297__34_,r_297__33_,r_297__32_,r_297__31_,
  r_297__30_,r_297__29_,r_297__28_,r_297__27_,r_297__26_,r_297__25_,r_297__24_,
  r_297__23_,r_297__22_,r_297__21_,r_297__20_,r_297__19_,r_297__18_,r_297__17_,r_297__16_,
  r_297__15_,r_297__14_,r_297__13_,r_297__12_,r_297__11_,r_297__10_,r_297__9_,
  r_297__8_,r_297__7_,r_297__6_,r_297__5_,r_297__4_,r_297__3_,r_297__2_,r_297__1_,
  r_297__0_,r_298__63_,r_298__62_,r_298__61_,r_298__60_,r_298__59_,r_298__58_,
  r_298__57_,r_298__56_,r_298__55_,r_298__54_,r_298__53_,r_298__52_,r_298__51_,r_298__50_,
  r_298__49_,r_298__48_,r_298__47_,r_298__46_,r_298__45_,r_298__44_,r_298__43_,
  r_298__42_,r_298__41_,r_298__40_,r_298__39_,r_298__38_,r_298__37_,r_298__36_,
  r_298__35_,r_298__34_,r_298__33_,r_298__32_,r_298__31_,r_298__30_,r_298__29_,
  r_298__28_,r_298__27_,r_298__26_,r_298__25_,r_298__24_,r_298__23_,r_298__22_,r_298__21_,
  r_298__20_,r_298__19_,r_298__18_,r_298__17_,r_298__16_,r_298__15_,r_298__14_,
  r_298__13_,r_298__12_,r_298__11_,r_298__10_,r_298__9_,r_298__8_,r_298__7_,r_298__6_,
  r_298__5_,r_298__4_,r_298__3_,r_298__2_,r_298__1_,r_298__0_,r_299__63_,
  r_299__62_,r_299__61_,r_299__60_,r_299__59_,r_299__58_,r_299__57_,r_299__56_,r_299__55_,
  r_299__54_,r_299__53_,r_299__52_,r_299__51_,r_299__50_,r_299__49_,r_299__48_,
  r_299__47_,r_299__46_,r_299__45_,r_299__44_,r_299__43_,r_299__42_,r_299__41_,
  r_299__40_,r_299__39_,r_299__38_,r_299__37_,r_299__36_,r_299__35_,r_299__34_,
  r_299__33_,r_299__32_,r_299__31_,r_299__30_,r_299__29_,r_299__28_,r_299__27_,r_299__26_,
  r_299__25_,r_299__24_,r_299__23_,r_299__22_,r_299__21_,r_299__20_,r_299__19_,
  r_299__18_,r_299__17_,r_299__16_,r_299__15_,r_299__14_,r_299__13_,r_299__12_,
  r_299__11_,r_299__10_,r_299__9_,r_299__8_,r_299__7_,r_299__6_,r_299__5_,r_299__4_,
  r_299__3_,r_299__2_,r_299__1_,r_299__0_,r_300__63_,r_300__62_,r_300__61_,r_300__60_,
  r_300__59_,r_300__58_,r_300__57_,r_300__56_,r_300__55_,r_300__54_,r_300__53_,
  r_300__52_,r_300__51_,r_300__50_,r_300__49_,r_300__48_,r_300__47_,r_300__46_,
  r_300__45_,r_300__44_,r_300__43_,r_300__42_,r_300__41_,r_300__40_,r_300__39_,r_300__38_,
  r_300__37_,r_300__36_,r_300__35_,r_300__34_,r_300__33_,r_300__32_,r_300__31_,
  r_300__30_,r_300__29_,r_300__28_,r_300__27_,r_300__26_,r_300__25_,r_300__24_,
  r_300__23_,r_300__22_,r_300__21_,r_300__20_,r_300__19_,r_300__18_,r_300__17_,
  r_300__16_,r_300__15_,r_300__14_,r_300__13_,r_300__12_,r_300__11_,r_300__10_,r_300__9_,
  r_300__8_,r_300__7_,r_300__6_,r_300__5_,r_300__4_,r_300__3_,r_300__2_,r_300__1_,
  r_300__0_,r_301__63_,r_301__62_,r_301__61_,r_301__60_,r_301__59_,r_301__58_,
  r_301__57_,r_301__56_,r_301__55_,r_301__54_,r_301__53_,r_301__52_,r_301__51_,
  r_301__50_,r_301__49_,r_301__48_,r_301__47_,r_301__46_,r_301__45_,r_301__44_,r_301__43_,
  r_301__42_,r_301__41_,r_301__40_,r_301__39_,r_301__38_,r_301__37_,r_301__36_,
  r_301__35_,r_301__34_,r_301__33_,r_301__32_,r_301__31_,r_301__30_,r_301__29_,
  r_301__28_,r_301__27_,r_301__26_,r_301__25_,r_301__24_,r_301__23_,r_301__22_,
  r_301__21_,r_301__20_,r_301__19_,r_301__18_,r_301__17_,r_301__16_,r_301__15_,r_301__14_,
  r_301__13_,r_301__12_,r_301__11_,r_301__10_,r_301__9_,r_301__8_,r_301__7_,
  r_301__6_,r_301__5_,r_301__4_,r_301__3_,r_301__2_,r_301__1_,r_301__0_,r_302__63_,
  r_302__62_,r_302__61_,r_302__60_,r_302__59_,r_302__58_,r_302__57_,r_302__56_,
  r_302__55_,r_302__54_,r_302__53_,r_302__52_,r_302__51_,r_302__50_,r_302__49_,r_302__48_,
  r_302__47_,r_302__46_,r_302__45_,r_302__44_,r_302__43_,r_302__42_,r_302__41_,
  r_302__40_,r_302__39_,r_302__38_,r_302__37_,r_302__36_,r_302__35_,r_302__34_,
  r_302__33_,r_302__32_,r_302__31_,r_302__30_,r_302__29_,r_302__28_,r_302__27_,r_302__26_,
  r_302__25_,r_302__24_,r_302__23_,r_302__22_,r_302__21_,r_302__20_,r_302__19_,
  r_302__18_,r_302__17_,r_302__16_,r_302__15_,r_302__14_,r_302__13_,r_302__12_,
  r_302__11_,r_302__10_,r_302__9_,r_302__8_,r_302__7_,r_302__6_,r_302__5_,r_302__4_,
  r_302__3_,r_302__2_,r_302__1_,r_302__0_,r_303__63_,r_303__62_,r_303__61_,r_303__60_,
  r_303__59_,r_303__58_,r_303__57_,r_303__56_,r_303__55_,r_303__54_,r_303__53_,
  r_303__52_,r_303__51_,r_303__50_,r_303__49_,r_303__48_,r_303__47_,r_303__46_,
  r_303__45_,r_303__44_,r_303__43_,r_303__42_,r_303__41_,r_303__40_,r_303__39_,
  r_303__38_,r_303__37_,r_303__36_,r_303__35_,r_303__34_,r_303__33_,r_303__32_,r_303__31_,
  r_303__30_,r_303__29_,r_303__28_,r_303__27_,r_303__26_,r_303__25_,r_303__24_,
  r_303__23_,r_303__22_,r_303__21_,r_303__20_,r_303__19_,r_303__18_,r_303__17_,
  r_303__16_,r_303__15_,r_303__14_,r_303__13_,r_303__12_,r_303__11_,r_303__10_,r_303__9_,
  r_303__8_,r_303__7_,r_303__6_,r_303__5_,r_303__4_,r_303__3_,r_303__2_,r_303__1_,
  r_303__0_,r_304__63_,r_304__62_,r_304__61_,r_304__60_,r_304__59_,r_304__58_,
  r_304__57_,r_304__56_,r_304__55_,r_304__54_,r_304__53_,r_304__52_,r_304__51_,
  r_304__50_,r_304__49_,r_304__48_,r_304__47_,r_304__46_,r_304__45_,r_304__44_,
  r_304__43_,r_304__42_,r_304__41_,r_304__40_,r_304__39_,r_304__38_,r_304__37_,r_304__36_,
  r_304__35_,r_304__34_,r_304__33_,r_304__32_,r_304__31_,r_304__30_,r_304__29_,
  r_304__28_,r_304__27_,r_304__26_,r_304__25_,r_304__24_,r_304__23_,r_304__22_,
  r_304__21_,r_304__20_,r_304__19_,r_304__18_,r_304__17_,r_304__16_,r_304__15_,r_304__14_,
  r_304__13_,r_304__12_,r_304__11_,r_304__10_,r_304__9_,r_304__8_,r_304__7_,
  r_304__6_,r_304__5_,r_304__4_,r_304__3_,r_304__2_,r_304__1_,r_304__0_,r_305__63_,
  r_305__62_,r_305__61_,r_305__60_,r_305__59_,r_305__58_,r_305__57_,r_305__56_,
  r_305__55_,r_305__54_,r_305__53_,r_305__52_,r_305__51_,r_305__50_,r_305__49_,r_305__48_,
  r_305__47_,r_305__46_,r_305__45_,r_305__44_,r_305__43_,r_305__42_,r_305__41_,
  r_305__40_,r_305__39_,r_305__38_,r_305__37_,r_305__36_,r_305__35_,r_305__34_,
  r_305__33_,r_305__32_,r_305__31_,r_305__30_,r_305__29_,r_305__28_,r_305__27_,
  r_305__26_,r_305__25_,r_305__24_,r_305__23_,r_305__22_,r_305__21_,r_305__20_,r_305__19_,
  r_305__18_,r_305__17_,r_305__16_,r_305__15_,r_305__14_,r_305__13_,r_305__12_,
  r_305__11_,r_305__10_,r_305__9_,r_305__8_,r_305__7_,r_305__6_,r_305__5_,r_305__4_,
  r_305__3_,r_305__2_,r_305__1_,r_305__0_,r_306__63_,r_306__62_,r_306__61_,
  r_306__60_,r_306__59_,r_306__58_,r_306__57_,r_306__56_,r_306__55_,r_306__54_,r_306__53_,
  r_306__52_,r_306__51_,r_306__50_,r_306__49_,r_306__48_,r_306__47_,r_306__46_,
  r_306__45_,r_306__44_,r_306__43_,r_306__42_,r_306__41_,r_306__40_,r_306__39_,
  r_306__38_,r_306__37_,r_306__36_,r_306__35_,r_306__34_,r_306__33_,r_306__32_,
  r_306__31_,r_306__30_,r_306__29_,r_306__28_,r_306__27_,r_306__26_,r_306__25_,r_306__24_,
  r_306__23_,r_306__22_,r_306__21_,r_306__20_,r_306__19_,r_306__18_,r_306__17_,
  r_306__16_,r_306__15_,r_306__14_,r_306__13_,r_306__12_,r_306__11_,r_306__10_,
  r_306__9_,r_306__8_,r_306__7_,r_306__6_,r_306__5_,r_306__4_,r_306__3_,r_306__2_,
  r_306__1_,r_306__0_,r_307__63_,r_307__62_,r_307__61_,r_307__60_,r_307__59_,r_307__58_,
  r_307__57_,r_307__56_,r_307__55_,r_307__54_,r_307__53_,r_307__52_,r_307__51_,
  r_307__50_,r_307__49_,r_307__48_,r_307__47_,r_307__46_,r_307__45_,r_307__44_,
  r_307__43_,r_307__42_,r_307__41_,r_307__40_,r_307__39_,r_307__38_,r_307__37_,r_307__36_,
  r_307__35_,r_307__34_,r_307__33_,r_307__32_,r_307__31_,r_307__30_,r_307__29_,
  r_307__28_,r_307__27_,r_307__26_,r_307__25_,r_307__24_,r_307__23_,r_307__22_,
  r_307__21_,r_307__20_,r_307__19_,r_307__18_,r_307__17_,r_307__16_,r_307__15_,
  r_307__14_,r_307__13_,r_307__12_,r_307__11_,r_307__10_,r_307__9_,r_307__8_,r_307__7_,
  r_307__6_,r_307__5_,r_307__4_,r_307__3_,r_307__2_,r_307__1_,r_307__0_,r_308__63_,
  r_308__62_,r_308__61_,r_308__60_,r_308__59_,r_308__58_,r_308__57_,r_308__56_,
  r_308__55_,r_308__54_,r_308__53_,r_308__52_,r_308__51_,r_308__50_,r_308__49_,
  r_308__48_,r_308__47_,r_308__46_,r_308__45_,r_308__44_,r_308__43_,r_308__42_,r_308__41_,
  r_308__40_,r_308__39_,r_308__38_,r_308__37_,r_308__36_,r_308__35_,r_308__34_,
  r_308__33_,r_308__32_,r_308__31_,r_308__30_,r_308__29_,r_308__28_,r_308__27_,
  r_308__26_,r_308__25_,r_308__24_,r_308__23_,r_308__22_,r_308__21_,r_308__20_,
  r_308__19_,r_308__18_,r_308__17_,r_308__16_,r_308__15_,r_308__14_,r_308__13_,r_308__12_,
  r_308__11_,r_308__10_,r_308__9_,r_308__8_,r_308__7_,r_308__6_,r_308__5_,r_308__4_,
  r_308__3_,r_308__2_,r_308__1_,r_308__0_,r_309__63_,r_309__62_,r_309__61_,
  r_309__60_,r_309__59_,r_309__58_,r_309__57_,r_309__56_,r_309__55_,r_309__54_,
  r_309__53_,r_309__52_,r_309__51_,r_309__50_,r_309__49_,r_309__48_,r_309__47_,r_309__46_,
  r_309__45_,r_309__44_,r_309__43_,r_309__42_,r_309__41_,r_309__40_,r_309__39_,
  r_309__38_,r_309__37_,r_309__36_,r_309__35_,r_309__34_,r_309__33_,r_309__32_,
  r_309__31_,r_309__30_,r_309__29_,r_309__28_,r_309__27_,r_309__26_,r_309__25_,r_309__24_,
  r_309__23_,r_309__22_,r_309__21_,r_309__20_,r_309__19_,r_309__18_,r_309__17_,
  r_309__16_,r_309__15_,r_309__14_,r_309__13_,r_309__12_,r_309__11_,r_309__10_,
  r_309__9_,r_309__8_,r_309__7_,r_309__6_,r_309__5_,r_309__4_,r_309__3_,r_309__2_,
  r_309__1_,r_309__0_,r_310__63_,r_310__62_,r_310__61_,r_310__60_,r_310__59_,r_310__58_,
  r_310__57_,r_310__56_,r_310__55_,r_310__54_,r_310__53_,r_310__52_,r_310__51_,
  r_310__50_,r_310__49_,r_310__48_,r_310__47_,r_310__46_,r_310__45_,r_310__44_,
  r_310__43_,r_310__42_,r_310__41_,r_310__40_,r_310__39_,r_310__38_,r_310__37_,
  r_310__36_,r_310__35_,r_310__34_,r_310__33_,r_310__32_,r_310__31_,r_310__30_,r_310__29_,
  r_310__28_,r_310__27_,r_310__26_,r_310__25_,r_310__24_,r_310__23_,r_310__22_,
  r_310__21_,r_310__20_,r_310__19_,r_310__18_,r_310__17_,r_310__16_,r_310__15_,
  r_310__14_,r_310__13_,r_310__12_,r_310__11_,r_310__10_,r_310__9_,r_310__8_,r_310__7_,
  r_310__6_,r_310__5_,r_310__4_,r_310__3_,r_310__2_,r_310__1_,r_310__0_,r_311__63_,
  r_311__62_,r_311__61_,r_311__60_,r_311__59_,r_311__58_,r_311__57_,r_311__56_,
  r_311__55_,r_311__54_,r_311__53_,r_311__52_,r_311__51_,r_311__50_,r_311__49_,
  r_311__48_,r_311__47_,r_311__46_,r_311__45_,r_311__44_,r_311__43_,r_311__42_,
  r_311__41_,r_311__40_,r_311__39_,r_311__38_,r_311__37_,r_311__36_,r_311__35_,r_311__34_,
  r_311__33_,r_311__32_,r_311__31_,r_311__30_,r_311__29_,r_311__28_,r_311__27_,
  r_311__26_,r_311__25_,r_311__24_,r_311__23_,r_311__22_,r_311__21_,r_311__20_,
  r_311__19_,r_311__18_,r_311__17_,r_311__16_,r_311__15_,r_311__14_,r_311__13_,r_311__12_,
  r_311__11_,r_311__10_,r_311__9_,r_311__8_,r_311__7_,r_311__6_,r_311__5_,
  r_311__4_,r_311__3_,r_311__2_,r_311__1_,r_311__0_,r_312__63_,r_312__62_,r_312__61_,
  r_312__60_,r_312__59_,r_312__58_,r_312__57_,r_312__56_,r_312__55_,r_312__54_,
  r_312__53_,r_312__52_,r_312__51_,r_312__50_,r_312__49_,r_312__48_,r_312__47_,r_312__46_,
  r_312__45_,r_312__44_,r_312__43_,r_312__42_,r_312__41_,r_312__40_,r_312__39_,
  r_312__38_,r_312__37_,r_312__36_,r_312__35_,r_312__34_,r_312__33_,r_312__32_,
  r_312__31_,r_312__30_,r_312__29_,r_312__28_,r_312__27_,r_312__26_,r_312__25_,
  r_312__24_,r_312__23_,r_312__22_,r_312__21_,r_312__20_,r_312__19_,r_312__18_,r_312__17_,
  r_312__16_,r_312__15_,r_312__14_,r_312__13_,r_312__12_,r_312__11_,r_312__10_,
  r_312__9_,r_312__8_,r_312__7_,r_312__6_,r_312__5_,r_312__4_,r_312__3_,r_312__2_,
  r_312__1_,r_312__0_,r_313__63_,r_313__62_,r_313__61_,r_313__60_,r_313__59_,
  r_313__58_,r_313__57_,r_313__56_,r_313__55_,r_313__54_,r_313__53_,r_313__52_,r_313__51_,
  r_313__50_,r_313__49_,r_313__48_,r_313__47_,r_313__46_,r_313__45_,r_313__44_,
  r_313__43_,r_313__42_,r_313__41_,r_313__40_,r_313__39_,r_313__38_,r_313__37_,
  r_313__36_,r_313__35_,r_313__34_,r_313__33_,r_313__32_,r_313__31_,r_313__30_,
  r_313__29_,r_313__28_,r_313__27_,r_313__26_,r_313__25_,r_313__24_,r_313__23_,r_313__22_,
  r_313__21_,r_313__20_,r_313__19_,r_313__18_,r_313__17_,r_313__16_,r_313__15_,
  r_313__14_,r_313__13_,r_313__12_,r_313__11_,r_313__10_,r_313__9_,r_313__8_,r_313__7_,
  r_313__6_,r_313__5_,r_313__4_,r_313__3_,r_313__2_,r_313__1_,r_313__0_,
  r_314__63_,r_314__62_,r_314__61_,r_314__60_,r_314__59_,r_314__58_,r_314__57_,r_314__56_,
  r_314__55_,r_314__54_,r_314__53_,r_314__52_,r_314__51_,r_314__50_,r_314__49_,
  r_314__48_,r_314__47_,r_314__46_,r_314__45_,r_314__44_,r_314__43_,r_314__42_,
  r_314__41_,r_314__40_,r_314__39_,r_314__38_,r_314__37_,r_314__36_,r_314__35_,r_314__34_,
  r_314__33_,r_314__32_,r_314__31_,r_314__30_,r_314__29_,r_314__28_,r_314__27_,
  r_314__26_,r_314__25_,r_314__24_,r_314__23_,r_314__22_,r_314__21_,r_314__20_,
  r_314__19_,r_314__18_,r_314__17_,r_314__16_,r_314__15_,r_314__14_,r_314__13_,
  r_314__12_,r_314__11_,r_314__10_,r_314__9_,r_314__8_,r_314__7_,r_314__6_,r_314__5_,
  r_314__4_,r_314__3_,r_314__2_,r_314__1_,r_314__0_,r_315__63_,r_315__62_,r_315__61_,
  r_315__60_,r_315__59_,r_315__58_,r_315__57_,r_315__56_,r_315__55_,r_315__54_,
  r_315__53_,r_315__52_,r_315__51_,r_315__50_,r_315__49_,r_315__48_,r_315__47_,
  r_315__46_,r_315__45_,r_315__44_,r_315__43_,r_315__42_,r_315__41_,r_315__40_,r_315__39_,
  r_315__38_,r_315__37_,r_315__36_,r_315__35_,r_315__34_,r_315__33_,r_315__32_,
  r_315__31_,r_315__30_,r_315__29_,r_315__28_,r_315__27_,r_315__26_,r_315__25_,
  r_315__24_,r_315__23_,r_315__22_,r_315__21_,r_315__20_,r_315__19_,r_315__18_,
  r_315__17_,r_315__16_,r_315__15_,r_315__14_,r_315__13_,r_315__12_,r_315__11_,r_315__10_,
  r_315__9_,r_315__8_,r_315__7_,r_315__6_,r_315__5_,r_315__4_,r_315__3_,r_315__2_,
  r_315__1_,r_315__0_,r_316__63_,r_316__62_,r_316__61_,r_316__60_,r_316__59_,
  r_316__58_,r_316__57_,r_316__56_,r_316__55_,r_316__54_,r_316__53_,r_316__52_,
  r_316__51_,r_316__50_,r_316__49_,r_316__48_,r_316__47_,r_316__46_,r_316__45_,r_316__44_,
  r_316__43_,r_316__42_,r_316__41_,r_316__40_,r_316__39_,r_316__38_,r_316__37_,
  r_316__36_,r_316__35_,r_316__34_,r_316__33_,r_316__32_,r_316__31_,r_316__30_,
  r_316__29_,r_316__28_,r_316__27_,r_316__26_,r_316__25_,r_316__24_,r_316__23_,r_316__22_,
  r_316__21_,r_316__20_,r_316__19_,r_316__18_,r_316__17_,r_316__16_,r_316__15_,
  r_316__14_,r_316__13_,r_316__12_,r_316__11_,r_316__10_,r_316__9_,r_316__8_,
  r_316__7_,r_316__6_,r_316__5_,r_316__4_,r_316__3_,r_316__2_,r_316__1_,r_316__0_,
  r_317__63_,r_317__62_,r_317__61_,r_317__60_,r_317__59_,r_317__58_,r_317__57_,r_317__56_,
  r_317__55_,r_317__54_,r_317__53_,r_317__52_,r_317__51_,r_317__50_,r_317__49_,
  r_317__48_,r_317__47_,r_317__46_,r_317__45_,r_317__44_,r_317__43_,r_317__42_,
  r_317__41_,r_317__40_,r_317__39_,r_317__38_,r_317__37_,r_317__36_,r_317__35_,
  r_317__34_,r_317__33_,r_317__32_,r_317__31_,r_317__30_,r_317__29_,r_317__28_,r_317__27_,
  r_317__26_,r_317__25_,r_317__24_,r_317__23_,r_317__22_,r_317__21_,r_317__20_,
  r_317__19_,r_317__18_,r_317__17_,r_317__16_,r_317__15_,r_317__14_,r_317__13_,
  r_317__12_,r_317__11_,r_317__10_,r_317__9_,r_317__8_,r_317__7_,r_317__6_,r_317__5_,
  r_317__4_,r_317__3_,r_317__2_,r_317__1_,r_317__0_,r_318__63_,r_318__62_,r_318__61_,
  r_318__60_,r_318__59_,r_318__58_,r_318__57_,r_318__56_,r_318__55_,r_318__54_,
  r_318__53_,r_318__52_,r_318__51_,r_318__50_,r_318__49_,r_318__48_,r_318__47_,
  r_318__46_,r_318__45_,r_318__44_,r_318__43_,r_318__42_,r_318__41_,r_318__40_,
  r_318__39_,r_318__38_,r_318__37_,r_318__36_,r_318__35_,r_318__34_,r_318__33_,r_318__32_,
  r_318__31_,r_318__30_,r_318__29_,r_318__28_,r_318__27_,r_318__26_,r_318__25_,
  r_318__24_,r_318__23_,r_318__22_,r_318__21_,r_318__20_,r_318__19_,r_318__18_,
  r_318__17_,r_318__16_,r_318__15_,r_318__14_,r_318__13_,r_318__12_,r_318__11_,r_318__10_,
  r_318__9_,r_318__8_,r_318__7_,r_318__6_,r_318__5_,r_318__4_,r_318__3_,r_318__2_,
  r_318__1_,r_318__0_,r_319__63_,r_319__62_,r_319__61_,r_319__60_,r_319__59_,
  r_319__58_,r_319__57_,r_319__56_,r_319__55_,r_319__54_,r_319__53_,r_319__52_,
  r_319__51_,r_319__50_,r_319__49_,r_319__48_,r_319__47_,r_319__46_,r_319__45_,r_319__44_,
  r_319__43_,r_319__42_,r_319__41_,r_319__40_,r_319__39_,r_319__38_,r_319__37_,
  r_319__36_,r_319__35_,r_319__34_,r_319__33_,r_319__32_,r_319__31_,r_319__30_,
  r_319__29_,r_319__28_,r_319__27_,r_319__26_,r_319__25_,r_319__24_,r_319__23_,
  r_319__22_,r_319__21_,r_319__20_,r_319__19_,r_319__18_,r_319__17_,r_319__16_,r_319__15_,
  r_319__14_,r_319__13_,r_319__12_,r_319__11_,r_319__10_,r_319__9_,r_319__8_,
  r_319__7_,r_319__6_,r_319__5_,r_319__4_,r_319__3_,r_319__2_,r_319__1_,r_319__0_,
  r_320__63_,r_320__62_,r_320__61_,r_320__60_,r_320__59_,r_320__58_,r_320__57_,
  r_320__56_,r_320__55_,r_320__54_,r_320__53_,r_320__52_,r_320__51_,r_320__50_,r_320__49_,
  r_320__48_,r_320__47_,r_320__46_,r_320__45_,r_320__44_,r_320__43_,r_320__42_,
  r_320__41_,r_320__40_,r_320__39_,r_320__38_,r_320__37_,r_320__36_,r_320__35_,
  r_320__34_,r_320__33_,r_320__32_,r_320__31_,r_320__30_,r_320__29_,r_320__28_,
  r_320__27_,r_320__26_,r_320__25_,r_320__24_,r_320__23_,r_320__22_,r_320__21_,r_320__20_,
  r_320__19_,r_320__18_,r_320__17_,r_320__16_,r_320__15_,r_320__14_,r_320__13_,
  r_320__12_,r_320__11_,r_320__10_,r_320__9_,r_320__8_,r_320__7_,r_320__6_,r_320__5_,
  r_320__4_,r_320__3_,r_320__2_,r_320__1_,r_320__0_,r_321__63_,r_321__62_,
  r_321__61_,r_321__60_,r_321__59_,r_321__58_,r_321__57_,r_321__56_,r_321__55_,r_321__54_,
  r_321__53_,r_321__52_,r_321__51_,r_321__50_,r_321__49_,r_321__48_,r_321__47_,
  r_321__46_,r_321__45_,r_321__44_,r_321__43_,r_321__42_,r_321__41_,r_321__40_,
  r_321__39_,r_321__38_,r_321__37_,r_321__36_,r_321__35_,r_321__34_,r_321__33_,r_321__32_,
  r_321__31_,r_321__30_,r_321__29_,r_321__28_,r_321__27_,r_321__26_,r_321__25_,
  r_321__24_,r_321__23_,r_321__22_,r_321__21_,r_321__20_,r_321__19_,r_321__18_,
  r_321__17_,r_321__16_,r_321__15_,r_321__14_,r_321__13_,r_321__12_,r_321__11_,
  r_321__10_,r_321__9_,r_321__8_,r_321__7_,r_321__6_,r_321__5_,r_321__4_,r_321__3_,
  r_321__2_,r_321__1_,r_321__0_,r_322__63_,r_322__62_,r_322__61_,r_322__60_,r_322__59_,
  r_322__58_,r_322__57_,r_322__56_,r_322__55_,r_322__54_,r_322__53_,r_322__52_,
  r_322__51_,r_322__50_,r_322__49_,r_322__48_,r_322__47_,r_322__46_,r_322__45_,
  r_322__44_,r_322__43_,r_322__42_,r_322__41_,r_322__40_,r_322__39_,r_322__38_,r_322__37_,
  r_322__36_,r_322__35_,r_322__34_,r_322__33_,r_322__32_,r_322__31_,r_322__30_,
  r_322__29_,r_322__28_,r_322__27_,r_322__26_,r_322__25_,r_322__24_,r_322__23_,
  r_322__22_,r_322__21_,r_322__20_,r_322__19_,r_322__18_,r_322__17_,r_322__16_,
  r_322__15_,r_322__14_,r_322__13_,r_322__12_,r_322__11_,r_322__10_,r_322__9_,r_322__8_,
  r_322__7_,r_322__6_,r_322__5_,r_322__4_,r_322__3_,r_322__2_,r_322__1_,r_322__0_,
  r_323__63_,r_323__62_,r_323__61_,r_323__60_,r_323__59_,r_323__58_,r_323__57_,
  r_323__56_,r_323__55_,r_323__54_,r_323__53_,r_323__52_,r_323__51_,r_323__50_,
  r_323__49_,r_323__48_,r_323__47_,r_323__46_,r_323__45_,r_323__44_,r_323__43_,r_323__42_,
  r_323__41_,r_323__40_,r_323__39_,r_323__38_,r_323__37_,r_323__36_,r_323__35_,
  r_323__34_,r_323__33_,r_323__32_,r_323__31_,r_323__30_,r_323__29_,r_323__28_,
  r_323__27_,r_323__26_,r_323__25_,r_323__24_,r_323__23_,r_323__22_,r_323__21_,r_323__20_,
  r_323__19_,r_323__18_,r_323__17_,r_323__16_,r_323__15_,r_323__14_,r_323__13_,
  r_323__12_,r_323__11_,r_323__10_,r_323__9_,r_323__8_,r_323__7_,r_323__6_,r_323__5_,
  r_323__4_,r_323__3_,r_323__2_,r_323__1_,r_323__0_,r_324__63_,r_324__62_,
  r_324__61_,r_324__60_,r_324__59_,r_324__58_,r_324__57_,r_324__56_,r_324__55_,r_324__54_,
  r_324__53_,r_324__52_,r_324__51_,r_324__50_,r_324__49_,r_324__48_,r_324__47_,
  r_324__46_,r_324__45_,r_324__44_,r_324__43_,r_324__42_,r_324__41_,r_324__40_,
  r_324__39_,r_324__38_,r_324__37_,r_324__36_,r_324__35_,r_324__34_,r_324__33_,
  r_324__32_,r_324__31_,r_324__30_,r_324__29_,r_324__28_,r_324__27_,r_324__26_,r_324__25_,
  r_324__24_,r_324__23_,r_324__22_,r_324__21_,r_324__20_,r_324__19_,r_324__18_,
  r_324__17_,r_324__16_,r_324__15_,r_324__14_,r_324__13_,r_324__12_,r_324__11_,
  r_324__10_,r_324__9_,r_324__8_,r_324__7_,r_324__6_,r_324__5_,r_324__4_,r_324__3_,
  r_324__2_,r_324__1_,r_324__0_,r_325__63_,r_325__62_,r_325__61_,r_325__60_,r_325__59_,
  r_325__58_,r_325__57_,r_325__56_,r_325__55_,r_325__54_,r_325__53_,r_325__52_,
  r_325__51_,r_325__50_,r_325__49_,r_325__48_,r_325__47_,r_325__46_,r_325__45_,
  r_325__44_,r_325__43_,r_325__42_,r_325__41_,r_325__40_,r_325__39_,r_325__38_,
  r_325__37_,r_325__36_,r_325__35_,r_325__34_,r_325__33_,r_325__32_,r_325__31_,r_325__30_,
  r_325__29_,r_325__28_,r_325__27_,r_325__26_,r_325__25_,r_325__24_,r_325__23_,
  r_325__22_,r_325__21_,r_325__20_,r_325__19_,r_325__18_,r_325__17_,r_325__16_,
  r_325__15_,r_325__14_,r_325__13_,r_325__12_,r_325__11_,r_325__10_,r_325__9_,r_325__8_,
  r_325__7_,r_325__6_,r_325__5_,r_325__4_,r_325__3_,r_325__2_,r_325__1_,r_325__0_,
  r_326__63_,r_326__62_,r_326__61_,r_326__60_,r_326__59_,r_326__58_,r_326__57_,
  r_326__56_,r_326__55_,r_326__54_,r_326__53_,r_326__52_,r_326__51_,r_326__50_,
  r_326__49_,r_326__48_,r_326__47_,r_326__46_,r_326__45_,r_326__44_,r_326__43_,r_326__42_,
  r_326__41_,r_326__40_,r_326__39_,r_326__38_,r_326__37_,r_326__36_,r_326__35_,
  r_326__34_,r_326__33_,r_326__32_,r_326__31_,r_326__30_,r_326__29_,r_326__28_,
  r_326__27_,r_326__26_,r_326__25_,r_326__24_,r_326__23_,r_326__22_,r_326__21_,
  r_326__20_,r_326__19_,r_326__18_,r_326__17_,r_326__16_,r_326__15_,r_326__14_,r_326__13_,
  r_326__12_,r_326__11_,r_326__10_,r_326__9_,r_326__8_,r_326__7_,r_326__6_,
  r_326__5_,r_326__4_,r_326__3_,r_326__2_,r_326__1_,r_326__0_,r_327__63_,r_327__62_,
  r_327__61_,r_327__60_,r_327__59_,r_327__58_,r_327__57_,r_327__56_,r_327__55_,
  r_327__54_,r_327__53_,r_327__52_,r_327__51_,r_327__50_,r_327__49_,r_327__48_,r_327__47_,
  r_327__46_,r_327__45_,r_327__44_,r_327__43_,r_327__42_,r_327__41_,r_327__40_,
  r_327__39_,r_327__38_,r_327__37_,r_327__36_,r_327__35_,r_327__34_,r_327__33_,
  r_327__32_,r_327__31_,r_327__30_,r_327__29_,r_327__28_,r_327__27_,r_327__26_,
  r_327__25_,r_327__24_,r_327__23_,r_327__22_,r_327__21_,r_327__20_,r_327__19_,r_327__18_,
  r_327__17_,r_327__16_,r_327__15_,r_327__14_,r_327__13_,r_327__12_,r_327__11_,
  r_327__10_,r_327__9_,r_327__8_,r_327__7_,r_327__6_,r_327__5_,r_327__4_,r_327__3_,
  r_327__2_,r_327__1_,r_327__0_,r_328__63_,r_328__62_,r_328__61_,r_328__60_,
  r_328__59_,r_328__58_,r_328__57_,r_328__56_,r_328__55_,r_328__54_,r_328__53_,r_328__52_,
  r_328__51_,r_328__50_,r_328__49_,r_328__48_,r_328__47_,r_328__46_,r_328__45_,
  r_328__44_,r_328__43_,r_328__42_,r_328__41_,r_328__40_,r_328__39_,r_328__38_,
  r_328__37_,r_328__36_,r_328__35_,r_328__34_,r_328__33_,r_328__32_,r_328__31_,r_328__30_,
  r_328__29_,r_328__28_,r_328__27_,r_328__26_,r_328__25_,r_328__24_,r_328__23_,
  r_328__22_,r_328__21_,r_328__20_,r_328__19_,r_328__18_,r_328__17_,r_328__16_,
  r_328__15_,r_328__14_,r_328__13_,r_328__12_,r_328__11_,r_328__10_,r_328__9_,r_328__8_,
  r_328__7_,r_328__6_,r_328__5_,r_328__4_,r_328__3_,r_328__2_,r_328__1_,r_328__0_,
  r_329__63_,r_329__62_,r_329__61_,r_329__60_,r_329__59_,r_329__58_,r_329__57_,
  r_329__56_,r_329__55_,r_329__54_,r_329__53_,r_329__52_,r_329__51_,r_329__50_,
  r_329__49_,r_329__48_,r_329__47_,r_329__46_,r_329__45_,r_329__44_,r_329__43_,
  r_329__42_,r_329__41_,r_329__40_,r_329__39_,r_329__38_,r_329__37_,r_329__36_,r_329__35_,
  r_329__34_,r_329__33_,r_329__32_,r_329__31_,r_329__30_,r_329__29_,r_329__28_,
  r_329__27_,r_329__26_,r_329__25_,r_329__24_,r_329__23_,r_329__22_,r_329__21_,
  r_329__20_,r_329__19_,r_329__18_,r_329__17_,r_329__16_,r_329__15_,r_329__14_,
  r_329__13_,r_329__12_,r_329__11_,r_329__10_,r_329__9_,r_329__8_,r_329__7_,r_329__6_,
  r_329__5_,r_329__4_,r_329__3_,r_329__2_,r_329__1_,r_329__0_,r_330__63_,r_330__62_,
  r_330__61_,r_330__60_,r_330__59_,r_330__58_,r_330__57_,r_330__56_,r_330__55_,
  r_330__54_,r_330__53_,r_330__52_,r_330__51_,r_330__50_,r_330__49_,r_330__48_,
  r_330__47_,r_330__46_,r_330__45_,r_330__44_,r_330__43_,r_330__42_,r_330__41_,r_330__40_,
  r_330__39_,r_330__38_,r_330__37_,r_330__36_,r_330__35_,r_330__34_,r_330__33_,
  r_330__32_,r_330__31_,r_330__30_,r_330__29_,r_330__28_,r_330__27_,r_330__26_,
  r_330__25_,r_330__24_,r_330__23_,r_330__22_,r_330__21_,r_330__20_,r_330__19_,r_330__18_,
  r_330__17_,r_330__16_,r_330__15_,r_330__14_,r_330__13_,r_330__12_,r_330__11_,
  r_330__10_,r_330__9_,r_330__8_,r_330__7_,r_330__6_,r_330__5_,r_330__4_,r_330__3_,
  r_330__2_,r_330__1_,r_330__0_,r_331__63_,r_331__62_,r_331__61_,r_331__60_,
  r_331__59_,r_331__58_,r_331__57_,r_331__56_,r_331__55_,r_331__54_,r_331__53_,r_331__52_,
  r_331__51_,r_331__50_,r_331__49_,r_331__48_,r_331__47_,r_331__46_,r_331__45_,
  r_331__44_,r_331__43_,r_331__42_,r_331__41_,r_331__40_,r_331__39_,r_331__38_,
  r_331__37_,r_331__36_,r_331__35_,r_331__34_,r_331__33_,r_331__32_,r_331__31_,
  r_331__30_,r_331__29_,r_331__28_,r_331__27_,r_331__26_,r_331__25_,r_331__24_,r_331__23_,
  r_331__22_,r_331__21_,r_331__20_,r_331__19_,r_331__18_,r_331__17_,r_331__16_,
  r_331__15_,r_331__14_,r_331__13_,r_331__12_,r_331__11_,r_331__10_,r_331__9_,
  r_331__8_,r_331__7_,r_331__6_,r_331__5_,r_331__4_,r_331__3_,r_331__2_,r_331__1_,
  r_331__0_,r_332__63_,r_332__62_,r_332__61_,r_332__60_,r_332__59_,r_332__58_,r_332__57_,
  r_332__56_,r_332__55_,r_332__54_,r_332__53_,r_332__52_,r_332__51_,r_332__50_,
  r_332__49_,r_332__48_,r_332__47_,r_332__46_,r_332__45_,r_332__44_,r_332__43_,
  r_332__42_,r_332__41_,r_332__40_,r_332__39_,r_332__38_,r_332__37_,r_332__36_,
  r_332__35_,r_332__34_,r_332__33_,r_332__32_,r_332__31_,r_332__30_,r_332__29_,r_332__28_,
  r_332__27_,r_332__26_,r_332__25_,r_332__24_,r_332__23_,r_332__22_,r_332__21_,
  r_332__20_,r_332__19_,r_332__18_,r_332__17_,r_332__16_,r_332__15_,r_332__14_,
  r_332__13_,r_332__12_,r_332__11_,r_332__10_,r_332__9_,r_332__8_,r_332__7_,r_332__6_,
  r_332__5_,r_332__4_,r_332__3_,r_332__2_,r_332__1_,r_332__0_,r_333__63_,r_333__62_,
  r_333__61_,r_333__60_,r_333__59_,r_333__58_,r_333__57_,r_333__56_,r_333__55_,
  r_333__54_,r_333__53_,r_333__52_,r_333__51_,r_333__50_,r_333__49_,r_333__48_,
  r_333__47_,r_333__46_,r_333__45_,r_333__44_,r_333__43_,r_333__42_,r_333__41_,r_333__40_,
  r_333__39_,r_333__38_,r_333__37_,r_333__36_,r_333__35_,r_333__34_,r_333__33_,
  r_333__32_,r_333__31_,r_333__30_,r_333__29_,r_333__28_,r_333__27_,r_333__26_,
  r_333__25_,r_333__24_,r_333__23_,r_333__22_,r_333__21_,r_333__20_,r_333__19_,
  r_333__18_,r_333__17_,r_333__16_,r_333__15_,r_333__14_,r_333__13_,r_333__12_,r_333__11_,
  r_333__10_,r_333__9_,r_333__8_,r_333__7_,r_333__6_,r_333__5_,r_333__4_,r_333__3_,
  r_333__2_,r_333__1_,r_333__0_,r_334__63_,r_334__62_,r_334__61_,r_334__60_,
  r_334__59_,r_334__58_,r_334__57_,r_334__56_,r_334__55_,r_334__54_,r_334__53_,
  r_334__52_,r_334__51_,r_334__50_,r_334__49_,r_334__48_,r_334__47_,r_334__46_,r_334__45_,
  r_334__44_,r_334__43_,r_334__42_,r_334__41_,r_334__40_,r_334__39_,r_334__38_,
  r_334__37_,r_334__36_,r_334__35_,r_334__34_,r_334__33_,r_334__32_,r_334__31_,
  r_334__30_,r_334__29_,r_334__28_,r_334__27_,r_334__26_,r_334__25_,r_334__24_,
  r_334__23_,r_334__22_,r_334__21_,r_334__20_,r_334__19_,r_334__18_,r_334__17_,r_334__16_,
  r_334__15_,r_334__14_,r_334__13_,r_334__12_,r_334__11_,r_334__10_,r_334__9_,
  r_334__8_,r_334__7_,r_334__6_,r_334__5_,r_334__4_,r_334__3_,r_334__2_,r_334__1_,
  r_334__0_,r_335__63_,r_335__62_,r_335__61_,r_335__60_,r_335__59_,r_335__58_,
  r_335__57_,r_335__56_,r_335__55_,r_335__54_,r_335__53_,r_335__52_,r_335__51_,r_335__50_,
  r_335__49_,r_335__48_,r_335__47_,r_335__46_,r_335__45_,r_335__44_,r_335__43_,
  r_335__42_,r_335__41_,r_335__40_,r_335__39_,r_335__38_,r_335__37_,r_335__36_,
  r_335__35_,r_335__34_,r_335__33_,r_335__32_,r_335__31_,r_335__30_,r_335__29_,r_335__28_,
  r_335__27_,r_335__26_,r_335__25_,r_335__24_,r_335__23_,r_335__22_,r_335__21_,
  r_335__20_,r_335__19_,r_335__18_,r_335__17_,r_335__16_,r_335__15_,r_335__14_,
  r_335__13_,r_335__12_,r_335__11_,r_335__10_,r_335__9_,r_335__8_,r_335__7_,r_335__6_,
  r_335__5_,r_335__4_,r_335__3_,r_335__2_,r_335__1_,r_335__0_,r_336__63_,r_336__62_,
  r_336__61_,r_336__60_,r_336__59_,r_336__58_,r_336__57_,r_336__56_,r_336__55_,
  r_336__54_,r_336__53_,r_336__52_,r_336__51_,r_336__50_,r_336__49_,r_336__48_,
  r_336__47_,r_336__46_,r_336__45_,r_336__44_,r_336__43_,r_336__42_,r_336__41_,
  r_336__40_,r_336__39_,r_336__38_,r_336__37_,r_336__36_,r_336__35_,r_336__34_,r_336__33_,
  r_336__32_,r_336__31_,r_336__30_,r_336__29_,r_336__28_,r_336__27_,r_336__26_,
  r_336__25_,r_336__24_,r_336__23_,r_336__22_,r_336__21_,r_336__20_,r_336__19_,
  r_336__18_,r_336__17_,r_336__16_,r_336__15_,r_336__14_,r_336__13_,r_336__12_,
  r_336__11_,r_336__10_,r_336__9_,r_336__8_,r_336__7_,r_336__6_,r_336__5_,r_336__4_,
  r_336__3_,r_336__2_,r_336__1_,r_336__0_,r_337__63_,r_337__62_,r_337__61_,r_337__60_,
  r_337__59_,r_337__58_,r_337__57_,r_337__56_,r_337__55_,r_337__54_,r_337__53_,
  r_337__52_,r_337__51_,r_337__50_,r_337__49_,r_337__48_,r_337__47_,r_337__46_,
  r_337__45_,r_337__44_,r_337__43_,r_337__42_,r_337__41_,r_337__40_,r_337__39_,r_337__38_,
  r_337__37_,r_337__36_,r_337__35_,r_337__34_,r_337__33_,r_337__32_,r_337__31_,
  r_337__30_,r_337__29_,r_337__28_,r_337__27_,r_337__26_,r_337__25_,r_337__24_,
  r_337__23_,r_337__22_,r_337__21_,r_337__20_,r_337__19_,r_337__18_,r_337__17_,r_337__16_,
  r_337__15_,r_337__14_,r_337__13_,r_337__12_,r_337__11_,r_337__10_,r_337__9_,
  r_337__8_,r_337__7_,r_337__6_,r_337__5_,r_337__4_,r_337__3_,r_337__2_,r_337__1_,
  r_337__0_,r_338__63_,r_338__62_,r_338__61_,r_338__60_,r_338__59_,r_338__58_,
  r_338__57_,r_338__56_,r_338__55_,r_338__54_,r_338__53_,r_338__52_,r_338__51_,r_338__50_,
  r_338__49_,r_338__48_,r_338__47_,r_338__46_,r_338__45_,r_338__44_,r_338__43_,
  r_338__42_,r_338__41_,r_338__40_,r_338__39_,r_338__38_,r_338__37_,r_338__36_,
  r_338__35_,r_338__34_,r_338__33_,r_338__32_,r_338__31_,r_338__30_,r_338__29_,
  r_338__28_,r_338__27_,r_338__26_,r_338__25_,r_338__24_,r_338__23_,r_338__22_,r_338__21_,
  r_338__20_,r_338__19_,r_338__18_,r_338__17_,r_338__16_,r_338__15_,r_338__14_,
  r_338__13_,r_338__12_,r_338__11_,r_338__10_,r_338__9_,r_338__8_,r_338__7_,r_338__6_,
  r_338__5_,r_338__4_,r_338__3_,r_338__2_,r_338__1_,r_338__0_,r_339__63_,
  r_339__62_,r_339__61_,r_339__60_,r_339__59_,r_339__58_,r_339__57_,r_339__56_,r_339__55_,
  r_339__54_,r_339__53_,r_339__52_,r_339__51_,r_339__50_,r_339__49_,r_339__48_,
  r_339__47_,r_339__46_,r_339__45_,r_339__44_,r_339__43_,r_339__42_,r_339__41_,
  r_339__40_,r_339__39_,r_339__38_,r_339__37_,r_339__36_,r_339__35_,r_339__34_,
  r_339__33_,r_339__32_,r_339__31_,r_339__30_,r_339__29_,r_339__28_,r_339__27_,r_339__26_,
  r_339__25_,r_339__24_,r_339__23_,r_339__22_,r_339__21_,r_339__20_,r_339__19_,
  r_339__18_,r_339__17_,r_339__16_,r_339__15_,r_339__14_,r_339__13_,r_339__12_,
  r_339__11_,r_339__10_,r_339__9_,r_339__8_,r_339__7_,r_339__6_,r_339__5_,r_339__4_,
  r_339__3_,r_339__2_,r_339__1_,r_339__0_,r_340__63_,r_340__62_,r_340__61_,r_340__60_,
  r_340__59_,r_340__58_,r_340__57_,r_340__56_,r_340__55_,r_340__54_,r_340__53_,
  r_340__52_,r_340__51_,r_340__50_,r_340__49_,r_340__48_,r_340__47_,r_340__46_,
  r_340__45_,r_340__44_,r_340__43_,r_340__42_,r_340__41_,r_340__40_,r_340__39_,r_340__38_,
  r_340__37_,r_340__36_,r_340__35_,r_340__34_,r_340__33_,r_340__32_,r_340__31_,
  r_340__30_,r_340__29_,r_340__28_,r_340__27_,r_340__26_,r_340__25_,r_340__24_,
  r_340__23_,r_340__22_,r_340__21_,r_340__20_,r_340__19_,r_340__18_,r_340__17_,
  r_340__16_,r_340__15_,r_340__14_,r_340__13_,r_340__12_,r_340__11_,r_340__10_,r_340__9_,
  r_340__8_,r_340__7_,r_340__6_,r_340__5_,r_340__4_,r_340__3_,r_340__2_,r_340__1_,
  r_340__0_,r_341__63_,r_341__62_,r_341__61_,r_341__60_,r_341__59_,r_341__58_,
  r_341__57_,r_341__56_,r_341__55_,r_341__54_,r_341__53_,r_341__52_,r_341__51_,
  r_341__50_,r_341__49_,r_341__48_,r_341__47_,r_341__46_,r_341__45_,r_341__44_,r_341__43_,
  r_341__42_,r_341__41_,r_341__40_,r_341__39_,r_341__38_,r_341__37_,r_341__36_,
  r_341__35_,r_341__34_,r_341__33_,r_341__32_,r_341__31_,r_341__30_,r_341__29_,
  r_341__28_,r_341__27_,r_341__26_,r_341__25_,r_341__24_,r_341__23_,r_341__22_,
  r_341__21_,r_341__20_,r_341__19_,r_341__18_,r_341__17_,r_341__16_,r_341__15_,r_341__14_,
  r_341__13_,r_341__12_,r_341__11_,r_341__10_,r_341__9_,r_341__8_,r_341__7_,
  r_341__6_,r_341__5_,r_341__4_,r_341__3_,r_341__2_,r_341__1_,r_341__0_,r_342__63_,
  r_342__62_,r_342__61_,r_342__60_,r_342__59_,r_342__58_,r_342__57_,r_342__56_,
  r_342__55_,r_342__54_,r_342__53_,r_342__52_,r_342__51_,r_342__50_,r_342__49_,r_342__48_,
  r_342__47_,r_342__46_,r_342__45_,r_342__44_,r_342__43_,r_342__42_,r_342__41_,
  r_342__40_,r_342__39_,r_342__38_,r_342__37_,r_342__36_,r_342__35_,r_342__34_,
  r_342__33_,r_342__32_,r_342__31_,r_342__30_,r_342__29_,r_342__28_,r_342__27_,r_342__26_,
  r_342__25_,r_342__24_,r_342__23_,r_342__22_,r_342__21_,r_342__20_,r_342__19_,
  r_342__18_,r_342__17_,r_342__16_,r_342__15_,r_342__14_,r_342__13_,r_342__12_,
  r_342__11_,r_342__10_,r_342__9_,r_342__8_,r_342__7_,r_342__6_,r_342__5_,r_342__4_,
  r_342__3_,r_342__2_,r_342__1_,r_342__0_,r_343__63_,r_343__62_,r_343__61_,r_343__60_,
  r_343__59_,r_343__58_,r_343__57_,r_343__56_,r_343__55_,r_343__54_,r_343__53_,
  r_343__52_,r_343__51_,r_343__50_,r_343__49_,r_343__48_,r_343__47_,r_343__46_,
  r_343__45_,r_343__44_,r_343__43_,r_343__42_,r_343__41_,r_343__40_,r_343__39_,
  r_343__38_,r_343__37_,r_343__36_,r_343__35_,r_343__34_,r_343__33_,r_343__32_,r_343__31_,
  r_343__30_,r_343__29_,r_343__28_,r_343__27_,r_343__26_,r_343__25_,r_343__24_,
  r_343__23_,r_343__22_,r_343__21_,r_343__20_,r_343__19_,r_343__18_,r_343__17_,
  r_343__16_,r_343__15_,r_343__14_,r_343__13_,r_343__12_,r_343__11_,r_343__10_,r_343__9_,
  r_343__8_,r_343__7_,r_343__6_,r_343__5_,r_343__4_,r_343__3_,r_343__2_,r_343__1_,
  r_343__0_,r_344__63_,r_344__62_,r_344__61_,r_344__60_,r_344__59_,r_344__58_,
  r_344__57_,r_344__56_,r_344__55_,r_344__54_,r_344__53_,r_344__52_,r_344__51_,
  r_344__50_,r_344__49_,r_344__48_,r_344__47_,r_344__46_,r_344__45_,r_344__44_,
  r_344__43_,r_344__42_,r_344__41_,r_344__40_,r_344__39_,r_344__38_,r_344__37_,r_344__36_,
  r_344__35_,r_344__34_,r_344__33_,r_344__32_,r_344__31_,r_344__30_,r_344__29_,
  r_344__28_,r_344__27_,r_344__26_,r_344__25_,r_344__24_,r_344__23_,r_344__22_,
  r_344__21_,r_344__20_,r_344__19_,r_344__18_,r_344__17_,r_344__16_,r_344__15_,r_344__14_,
  r_344__13_,r_344__12_,r_344__11_,r_344__10_,r_344__9_,r_344__8_,r_344__7_,
  r_344__6_,r_344__5_,r_344__4_,r_344__3_,r_344__2_,r_344__1_,r_344__0_,r_345__63_,
  r_345__62_,r_345__61_,r_345__60_,r_345__59_,r_345__58_,r_345__57_,r_345__56_,
  r_345__55_,r_345__54_,r_345__53_,r_345__52_,r_345__51_,r_345__50_,r_345__49_,r_345__48_,
  r_345__47_,r_345__46_,r_345__45_,r_345__44_,r_345__43_,r_345__42_,r_345__41_,
  r_345__40_,r_345__39_,r_345__38_,r_345__37_,r_345__36_,r_345__35_,r_345__34_,
  r_345__33_,r_345__32_,r_345__31_,r_345__30_,r_345__29_,r_345__28_,r_345__27_,
  r_345__26_,r_345__25_,r_345__24_,r_345__23_,r_345__22_,r_345__21_,r_345__20_,r_345__19_,
  r_345__18_,r_345__17_,r_345__16_,r_345__15_,r_345__14_,r_345__13_,r_345__12_,
  r_345__11_,r_345__10_,r_345__9_,r_345__8_,r_345__7_,r_345__6_,r_345__5_,r_345__4_,
  r_345__3_,r_345__2_,r_345__1_,r_345__0_,r_346__63_,r_346__62_,r_346__61_,
  r_346__60_,r_346__59_,r_346__58_,r_346__57_,r_346__56_,r_346__55_,r_346__54_,r_346__53_,
  r_346__52_,r_346__51_,r_346__50_,r_346__49_,r_346__48_,r_346__47_,r_346__46_,
  r_346__45_,r_346__44_,r_346__43_,r_346__42_,r_346__41_,r_346__40_,r_346__39_,
  r_346__38_,r_346__37_,r_346__36_,r_346__35_,r_346__34_,r_346__33_,r_346__32_,
  r_346__31_,r_346__30_,r_346__29_,r_346__28_,r_346__27_,r_346__26_,r_346__25_,r_346__24_,
  r_346__23_,r_346__22_,r_346__21_,r_346__20_,r_346__19_,r_346__18_,r_346__17_,
  r_346__16_,r_346__15_,r_346__14_,r_346__13_,r_346__12_,r_346__11_,r_346__10_,
  r_346__9_,r_346__8_,r_346__7_,r_346__6_,r_346__5_,r_346__4_,r_346__3_,r_346__2_,
  r_346__1_,r_346__0_,r_347__63_,r_347__62_,r_347__61_,r_347__60_,r_347__59_,r_347__58_,
  r_347__57_,r_347__56_,r_347__55_,r_347__54_,r_347__53_,r_347__52_,r_347__51_,
  r_347__50_,r_347__49_,r_347__48_,r_347__47_,r_347__46_,r_347__45_,r_347__44_,
  r_347__43_,r_347__42_,r_347__41_,r_347__40_,r_347__39_,r_347__38_,r_347__37_,r_347__36_,
  r_347__35_,r_347__34_,r_347__33_,r_347__32_,r_347__31_,r_347__30_,r_347__29_,
  r_347__28_,r_347__27_,r_347__26_,r_347__25_,r_347__24_,r_347__23_,r_347__22_,
  r_347__21_,r_347__20_,r_347__19_,r_347__18_,r_347__17_,r_347__16_,r_347__15_,
  r_347__14_,r_347__13_,r_347__12_,r_347__11_,r_347__10_,r_347__9_,r_347__8_,r_347__7_,
  r_347__6_,r_347__5_,r_347__4_,r_347__3_,r_347__2_,r_347__1_,r_347__0_,r_348__63_,
  r_348__62_,r_348__61_,r_348__60_,r_348__59_,r_348__58_,r_348__57_,r_348__56_,
  r_348__55_,r_348__54_,r_348__53_,r_348__52_,r_348__51_,r_348__50_,r_348__49_,
  r_348__48_,r_348__47_,r_348__46_,r_348__45_,r_348__44_,r_348__43_,r_348__42_,r_348__41_,
  r_348__40_,r_348__39_,r_348__38_,r_348__37_,r_348__36_,r_348__35_,r_348__34_,
  r_348__33_,r_348__32_,r_348__31_,r_348__30_,r_348__29_,r_348__28_,r_348__27_,
  r_348__26_,r_348__25_,r_348__24_,r_348__23_,r_348__22_,r_348__21_,r_348__20_,
  r_348__19_,r_348__18_,r_348__17_,r_348__16_,r_348__15_,r_348__14_,r_348__13_,r_348__12_,
  r_348__11_,r_348__10_,r_348__9_,r_348__8_,r_348__7_,r_348__6_,r_348__5_,r_348__4_,
  r_348__3_,r_348__2_,r_348__1_,r_348__0_,r_349__63_,r_349__62_,r_349__61_,
  r_349__60_,r_349__59_,r_349__58_,r_349__57_,r_349__56_,r_349__55_,r_349__54_,
  r_349__53_,r_349__52_,r_349__51_,r_349__50_,r_349__49_,r_349__48_,r_349__47_,r_349__46_,
  r_349__45_,r_349__44_,r_349__43_,r_349__42_,r_349__41_,r_349__40_,r_349__39_,
  r_349__38_,r_349__37_,r_349__36_,r_349__35_,r_349__34_,r_349__33_,r_349__32_,
  r_349__31_,r_349__30_,r_349__29_,r_349__28_,r_349__27_,r_349__26_,r_349__25_,r_349__24_,
  r_349__23_,r_349__22_,r_349__21_,r_349__20_,r_349__19_,r_349__18_,r_349__17_,
  r_349__16_,r_349__15_,r_349__14_,r_349__13_,r_349__12_,r_349__11_,r_349__10_,
  r_349__9_,r_349__8_,r_349__7_,r_349__6_,r_349__5_,r_349__4_,r_349__3_,r_349__2_,
  r_349__1_,r_349__0_,r_350__63_,r_350__62_,r_350__61_,r_350__60_,r_350__59_,r_350__58_,
  r_350__57_,r_350__56_,r_350__55_,r_350__54_,r_350__53_,r_350__52_,r_350__51_,
  r_350__50_,r_350__49_,r_350__48_,r_350__47_,r_350__46_,r_350__45_,r_350__44_,
  r_350__43_,r_350__42_,r_350__41_,r_350__40_,r_350__39_,r_350__38_,r_350__37_,
  r_350__36_,r_350__35_,r_350__34_,r_350__33_,r_350__32_,r_350__31_,r_350__30_,r_350__29_,
  r_350__28_,r_350__27_,r_350__26_,r_350__25_,r_350__24_,r_350__23_,r_350__22_,
  r_350__21_,r_350__20_,r_350__19_,r_350__18_,r_350__17_,r_350__16_,r_350__15_,
  r_350__14_,r_350__13_,r_350__12_,r_350__11_,r_350__10_,r_350__9_,r_350__8_,r_350__7_,
  r_350__6_,r_350__5_,r_350__4_,r_350__3_,r_350__2_,r_350__1_,r_350__0_,r_351__63_,
  r_351__62_,r_351__61_,r_351__60_,r_351__59_,r_351__58_,r_351__57_,r_351__56_,
  r_351__55_,r_351__54_,r_351__53_,r_351__52_,r_351__51_,r_351__50_,r_351__49_,
  r_351__48_,r_351__47_,r_351__46_,r_351__45_,r_351__44_,r_351__43_,r_351__42_,
  r_351__41_,r_351__40_,r_351__39_,r_351__38_,r_351__37_,r_351__36_,r_351__35_,r_351__34_,
  r_351__33_,r_351__32_,r_351__31_,r_351__30_,r_351__29_,r_351__28_,r_351__27_,
  r_351__26_,r_351__25_,r_351__24_,r_351__23_,r_351__22_,r_351__21_,r_351__20_,
  r_351__19_,r_351__18_,r_351__17_,r_351__16_,r_351__15_,r_351__14_,r_351__13_,r_351__12_,
  r_351__11_,r_351__10_,r_351__9_,r_351__8_,r_351__7_,r_351__6_,r_351__5_,
  r_351__4_,r_351__3_,r_351__2_,r_351__1_,r_351__0_,r_352__63_,r_352__62_,r_352__61_,
  r_352__60_,r_352__59_,r_352__58_,r_352__57_,r_352__56_,r_352__55_,r_352__54_,
  r_352__53_,r_352__52_,r_352__51_,r_352__50_,r_352__49_,r_352__48_,r_352__47_,r_352__46_,
  r_352__45_,r_352__44_,r_352__43_,r_352__42_,r_352__41_,r_352__40_,r_352__39_,
  r_352__38_,r_352__37_,r_352__36_,r_352__35_,r_352__34_,r_352__33_,r_352__32_,
  r_352__31_,r_352__30_,r_352__29_,r_352__28_,r_352__27_,r_352__26_,r_352__25_,
  r_352__24_,r_352__23_,r_352__22_,r_352__21_,r_352__20_,r_352__19_,r_352__18_,r_352__17_,
  r_352__16_,r_352__15_,r_352__14_,r_352__13_,r_352__12_,r_352__11_,r_352__10_,
  r_352__9_,r_352__8_,r_352__7_,r_352__6_,r_352__5_,r_352__4_,r_352__3_,r_352__2_,
  r_352__1_,r_352__0_,r_353__63_,r_353__62_,r_353__61_,r_353__60_,r_353__59_,
  r_353__58_,r_353__57_,r_353__56_,r_353__55_,r_353__54_,r_353__53_,r_353__52_,r_353__51_,
  r_353__50_,r_353__49_,r_353__48_,r_353__47_,r_353__46_,r_353__45_,r_353__44_,
  r_353__43_,r_353__42_,r_353__41_,r_353__40_,r_353__39_,r_353__38_,r_353__37_,
  r_353__36_,r_353__35_,r_353__34_,r_353__33_,r_353__32_,r_353__31_,r_353__30_,
  r_353__29_,r_353__28_,r_353__27_,r_353__26_,r_353__25_,r_353__24_,r_353__23_,r_353__22_,
  r_353__21_,r_353__20_,r_353__19_,r_353__18_,r_353__17_,r_353__16_,r_353__15_,
  r_353__14_,r_353__13_,r_353__12_,r_353__11_,r_353__10_,r_353__9_,r_353__8_,r_353__7_,
  r_353__6_,r_353__5_,r_353__4_,r_353__3_,r_353__2_,r_353__1_,r_353__0_,
  r_354__63_,r_354__62_,r_354__61_,r_354__60_,r_354__59_,r_354__58_,r_354__57_,r_354__56_,
  r_354__55_,r_354__54_,r_354__53_,r_354__52_,r_354__51_,r_354__50_,r_354__49_,
  r_354__48_,r_354__47_,r_354__46_,r_354__45_,r_354__44_,r_354__43_,r_354__42_,
  r_354__41_,r_354__40_,r_354__39_,r_354__38_,r_354__37_,r_354__36_,r_354__35_,r_354__34_,
  r_354__33_,r_354__32_,r_354__31_,r_354__30_,r_354__29_,r_354__28_,r_354__27_,
  r_354__26_,r_354__25_,r_354__24_,r_354__23_,r_354__22_,r_354__21_,r_354__20_,
  r_354__19_,r_354__18_,r_354__17_,r_354__16_,r_354__15_,r_354__14_,r_354__13_,
  r_354__12_,r_354__11_,r_354__10_,r_354__9_,r_354__8_,r_354__7_,r_354__6_,r_354__5_,
  r_354__4_,r_354__3_,r_354__2_,r_354__1_,r_354__0_,r_355__63_,r_355__62_,r_355__61_,
  r_355__60_,r_355__59_,r_355__58_,r_355__57_,r_355__56_,r_355__55_,r_355__54_,
  r_355__53_,r_355__52_,r_355__51_,r_355__50_,r_355__49_,r_355__48_,r_355__47_,
  r_355__46_,r_355__45_,r_355__44_,r_355__43_,r_355__42_,r_355__41_,r_355__40_,r_355__39_,
  r_355__38_,r_355__37_,r_355__36_,r_355__35_,r_355__34_,r_355__33_,r_355__32_,
  r_355__31_,r_355__30_,r_355__29_,r_355__28_,r_355__27_,r_355__26_,r_355__25_,
  r_355__24_,r_355__23_,r_355__22_,r_355__21_,r_355__20_,r_355__19_,r_355__18_,
  r_355__17_,r_355__16_,r_355__15_,r_355__14_,r_355__13_,r_355__12_,r_355__11_,r_355__10_,
  r_355__9_,r_355__8_,r_355__7_,r_355__6_,r_355__5_,r_355__4_,r_355__3_,r_355__2_,
  r_355__1_,r_355__0_,r_356__63_,r_356__62_,r_356__61_,r_356__60_,r_356__59_,
  r_356__58_,r_356__57_,r_356__56_,r_356__55_,r_356__54_,r_356__53_,r_356__52_,
  r_356__51_,r_356__50_,r_356__49_,r_356__48_,r_356__47_,r_356__46_,r_356__45_,r_356__44_,
  r_356__43_,r_356__42_,r_356__41_,r_356__40_,r_356__39_,r_356__38_,r_356__37_,
  r_356__36_,r_356__35_,r_356__34_,r_356__33_,r_356__32_,r_356__31_,r_356__30_,
  r_356__29_,r_356__28_,r_356__27_,r_356__26_,r_356__25_,r_356__24_,r_356__23_,r_356__22_,
  r_356__21_,r_356__20_,r_356__19_,r_356__18_,r_356__17_,r_356__16_,r_356__15_,
  r_356__14_,r_356__13_,r_356__12_,r_356__11_,r_356__10_,r_356__9_,r_356__8_,
  r_356__7_,r_356__6_,r_356__5_,r_356__4_,r_356__3_,r_356__2_,r_356__1_,r_356__0_,
  r_357__63_,r_357__62_,r_357__61_,r_357__60_,r_357__59_,r_357__58_,r_357__57_,r_357__56_,
  r_357__55_,r_357__54_,r_357__53_,r_357__52_,r_357__51_,r_357__50_,r_357__49_,
  r_357__48_,r_357__47_,r_357__46_,r_357__45_,r_357__44_,r_357__43_,r_357__42_,
  r_357__41_,r_357__40_,r_357__39_,r_357__38_,r_357__37_,r_357__36_,r_357__35_,
  r_357__34_,r_357__33_,r_357__32_,r_357__31_,r_357__30_,r_357__29_,r_357__28_,r_357__27_,
  r_357__26_,r_357__25_,r_357__24_,r_357__23_,r_357__22_,r_357__21_,r_357__20_,
  r_357__19_,r_357__18_,r_357__17_,r_357__16_,r_357__15_,r_357__14_,r_357__13_,
  r_357__12_,r_357__11_,r_357__10_,r_357__9_,r_357__8_,r_357__7_,r_357__6_,r_357__5_,
  r_357__4_,r_357__3_,r_357__2_,r_357__1_,r_357__0_,r_358__63_,r_358__62_,r_358__61_,
  r_358__60_,r_358__59_,r_358__58_,r_358__57_,r_358__56_,r_358__55_,r_358__54_,
  r_358__53_,r_358__52_,r_358__51_,r_358__50_,r_358__49_,r_358__48_,r_358__47_,
  r_358__46_,r_358__45_,r_358__44_,r_358__43_,r_358__42_,r_358__41_,r_358__40_,
  r_358__39_,r_358__38_,r_358__37_,r_358__36_,r_358__35_,r_358__34_,r_358__33_,r_358__32_,
  r_358__31_,r_358__30_,r_358__29_,r_358__28_,r_358__27_,r_358__26_,r_358__25_,
  r_358__24_,r_358__23_,r_358__22_,r_358__21_,r_358__20_,r_358__19_,r_358__18_,
  r_358__17_,r_358__16_,r_358__15_,r_358__14_,r_358__13_,r_358__12_,r_358__11_,r_358__10_,
  r_358__9_,r_358__8_,r_358__7_,r_358__6_,r_358__5_,r_358__4_,r_358__3_,r_358__2_,
  r_358__1_,r_358__0_,r_359__63_,r_359__62_,r_359__61_,r_359__60_,r_359__59_,
  r_359__58_,r_359__57_,r_359__56_,r_359__55_,r_359__54_,r_359__53_,r_359__52_,
  r_359__51_,r_359__50_,r_359__49_,r_359__48_,r_359__47_,r_359__46_,r_359__45_,r_359__44_,
  r_359__43_,r_359__42_,r_359__41_,r_359__40_,r_359__39_,r_359__38_,r_359__37_,
  r_359__36_,r_359__35_,r_359__34_,r_359__33_,r_359__32_,r_359__31_,r_359__30_,
  r_359__29_,r_359__28_,r_359__27_,r_359__26_,r_359__25_,r_359__24_,r_359__23_,
  r_359__22_,r_359__21_,r_359__20_,r_359__19_,r_359__18_,r_359__17_,r_359__16_,r_359__15_,
  r_359__14_,r_359__13_,r_359__12_,r_359__11_,r_359__10_,r_359__9_,r_359__8_,
  r_359__7_,r_359__6_,r_359__5_,r_359__4_,r_359__3_,r_359__2_,r_359__1_,r_359__0_,
  r_360__63_,r_360__62_,r_360__61_,r_360__60_,r_360__59_,r_360__58_,r_360__57_,
  r_360__56_,r_360__55_,r_360__54_,r_360__53_,r_360__52_,r_360__51_,r_360__50_,r_360__49_,
  r_360__48_,r_360__47_,r_360__46_,r_360__45_,r_360__44_,r_360__43_,r_360__42_,
  r_360__41_,r_360__40_,r_360__39_,r_360__38_,r_360__37_,r_360__36_,r_360__35_,
  r_360__34_,r_360__33_,r_360__32_,r_360__31_,r_360__30_,r_360__29_,r_360__28_,
  r_360__27_,r_360__26_,r_360__25_,r_360__24_,r_360__23_,r_360__22_,r_360__21_,r_360__20_,
  r_360__19_,r_360__18_,r_360__17_,r_360__16_,r_360__15_,r_360__14_,r_360__13_,
  r_360__12_,r_360__11_,r_360__10_,r_360__9_,r_360__8_,r_360__7_,r_360__6_,r_360__5_,
  r_360__4_,r_360__3_,r_360__2_,r_360__1_,r_360__0_,r_361__63_,r_361__62_,
  r_361__61_,r_361__60_,r_361__59_,r_361__58_,r_361__57_,r_361__56_,r_361__55_,r_361__54_,
  r_361__53_,r_361__52_,r_361__51_,r_361__50_,r_361__49_,r_361__48_,r_361__47_,
  r_361__46_,r_361__45_,r_361__44_,r_361__43_,r_361__42_,r_361__41_,r_361__40_,
  r_361__39_,r_361__38_,r_361__37_,r_361__36_,r_361__35_,r_361__34_,r_361__33_,r_361__32_,
  r_361__31_,r_361__30_,r_361__29_,r_361__28_,r_361__27_,r_361__26_,r_361__25_,
  r_361__24_,r_361__23_,r_361__22_,r_361__21_,r_361__20_,r_361__19_,r_361__18_,
  r_361__17_,r_361__16_,r_361__15_,r_361__14_,r_361__13_,r_361__12_,r_361__11_,
  r_361__10_,r_361__9_,r_361__8_,r_361__7_,r_361__6_,r_361__5_,r_361__4_,r_361__3_,
  r_361__2_,r_361__1_,r_361__0_,r_362__63_,r_362__62_,r_362__61_,r_362__60_,r_362__59_,
  r_362__58_,r_362__57_,r_362__56_,r_362__55_,r_362__54_,r_362__53_,r_362__52_,
  r_362__51_,r_362__50_,r_362__49_,r_362__48_,r_362__47_,r_362__46_,r_362__45_,
  r_362__44_,r_362__43_,r_362__42_,r_362__41_,r_362__40_,r_362__39_,r_362__38_,r_362__37_,
  r_362__36_,r_362__35_,r_362__34_,r_362__33_,r_362__32_,r_362__31_,r_362__30_,
  r_362__29_,r_362__28_,r_362__27_,r_362__26_,r_362__25_,r_362__24_,r_362__23_,
  r_362__22_,r_362__21_,r_362__20_,r_362__19_,r_362__18_,r_362__17_,r_362__16_,
  r_362__15_,r_362__14_,r_362__13_,r_362__12_,r_362__11_,r_362__10_,r_362__9_,r_362__8_,
  r_362__7_,r_362__6_,r_362__5_,r_362__4_,r_362__3_,r_362__2_,r_362__1_,r_362__0_,
  r_363__63_,r_363__62_,r_363__61_,r_363__60_,r_363__59_,r_363__58_,r_363__57_,
  r_363__56_,r_363__55_,r_363__54_,r_363__53_,r_363__52_,r_363__51_,r_363__50_,
  r_363__49_,r_363__48_,r_363__47_,r_363__46_,r_363__45_,r_363__44_,r_363__43_,r_363__42_,
  r_363__41_,r_363__40_,r_363__39_,r_363__38_,r_363__37_,r_363__36_,r_363__35_,
  r_363__34_,r_363__33_,r_363__32_,r_363__31_,r_363__30_,r_363__29_,r_363__28_,
  r_363__27_,r_363__26_,r_363__25_,r_363__24_,r_363__23_,r_363__22_,r_363__21_,r_363__20_,
  r_363__19_,r_363__18_,r_363__17_,r_363__16_,r_363__15_,r_363__14_,r_363__13_,
  r_363__12_,r_363__11_,r_363__10_,r_363__9_,r_363__8_,r_363__7_,r_363__6_,r_363__5_,
  r_363__4_,r_363__3_,r_363__2_,r_363__1_,r_363__0_,r_364__63_,r_364__62_,
  r_364__61_,r_364__60_,r_364__59_,r_364__58_,r_364__57_,r_364__56_,r_364__55_,r_364__54_,
  r_364__53_,r_364__52_,r_364__51_,r_364__50_,r_364__49_,r_364__48_,r_364__47_,
  r_364__46_,r_364__45_,r_364__44_,r_364__43_,r_364__42_,r_364__41_,r_364__40_,
  r_364__39_,r_364__38_,r_364__37_,r_364__36_,r_364__35_,r_364__34_,r_364__33_,
  r_364__32_,r_364__31_,r_364__30_,r_364__29_,r_364__28_,r_364__27_,r_364__26_,r_364__25_,
  r_364__24_,r_364__23_,r_364__22_,r_364__21_,r_364__20_,r_364__19_,r_364__18_,
  r_364__17_,r_364__16_,r_364__15_,r_364__14_,r_364__13_,r_364__12_,r_364__11_,
  r_364__10_,r_364__9_,r_364__8_,r_364__7_,r_364__6_,r_364__5_,r_364__4_,r_364__3_,
  r_364__2_,r_364__1_,r_364__0_,r_365__63_,r_365__62_,r_365__61_,r_365__60_,r_365__59_,
  r_365__58_,r_365__57_,r_365__56_,r_365__55_,r_365__54_,r_365__53_,r_365__52_,
  r_365__51_,r_365__50_,r_365__49_,r_365__48_,r_365__47_,r_365__46_,r_365__45_,
  r_365__44_,r_365__43_,r_365__42_,r_365__41_,r_365__40_,r_365__39_,r_365__38_,
  r_365__37_,r_365__36_,r_365__35_,r_365__34_,r_365__33_,r_365__32_,r_365__31_,r_365__30_,
  r_365__29_,r_365__28_,r_365__27_,r_365__26_,r_365__25_,r_365__24_,r_365__23_,
  r_365__22_,r_365__21_,r_365__20_,r_365__19_,r_365__18_,r_365__17_,r_365__16_,
  r_365__15_,r_365__14_,r_365__13_,r_365__12_,r_365__11_,r_365__10_,r_365__9_,r_365__8_,
  r_365__7_,r_365__6_,r_365__5_,r_365__4_,r_365__3_,r_365__2_,r_365__1_,r_365__0_,
  r_366__63_,r_366__62_,r_366__61_,r_366__60_,r_366__59_,r_366__58_,r_366__57_,
  r_366__56_,r_366__55_,r_366__54_,r_366__53_,r_366__52_,r_366__51_,r_366__50_,
  r_366__49_,r_366__48_,r_366__47_,r_366__46_,r_366__45_,r_366__44_,r_366__43_,r_366__42_,
  r_366__41_,r_366__40_,r_366__39_,r_366__38_,r_366__37_,r_366__36_,r_366__35_,
  r_366__34_,r_366__33_,r_366__32_,r_366__31_,r_366__30_,r_366__29_,r_366__28_,
  r_366__27_,r_366__26_,r_366__25_,r_366__24_,r_366__23_,r_366__22_,r_366__21_,
  r_366__20_,r_366__19_,r_366__18_,r_366__17_,r_366__16_,r_366__15_,r_366__14_,r_366__13_,
  r_366__12_,r_366__11_,r_366__10_,r_366__9_,r_366__8_,r_366__7_,r_366__6_,
  r_366__5_,r_366__4_,r_366__3_,r_366__2_,r_366__1_,r_366__0_,r_367__63_,r_367__62_,
  r_367__61_,r_367__60_,r_367__59_,r_367__58_,r_367__57_,r_367__56_,r_367__55_,
  r_367__54_,r_367__53_,r_367__52_,r_367__51_,r_367__50_,r_367__49_,r_367__48_,r_367__47_,
  r_367__46_,r_367__45_,r_367__44_,r_367__43_,r_367__42_,r_367__41_,r_367__40_,
  r_367__39_,r_367__38_,r_367__37_,r_367__36_,r_367__35_,r_367__34_,r_367__33_,
  r_367__32_,r_367__31_,r_367__30_,r_367__29_,r_367__28_,r_367__27_,r_367__26_,
  r_367__25_,r_367__24_,r_367__23_,r_367__22_,r_367__21_,r_367__20_,r_367__19_,r_367__18_,
  r_367__17_,r_367__16_,r_367__15_,r_367__14_,r_367__13_,r_367__12_,r_367__11_,
  r_367__10_,r_367__9_,r_367__8_,r_367__7_,r_367__6_,r_367__5_,r_367__4_,r_367__3_,
  r_367__2_,r_367__1_,r_367__0_,r_368__63_,r_368__62_,r_368__61_,r_368__60_,
  r_368__59_,r_368__58_,r_368__57_,r_368__56_,r_368__55_,r_368__54_,r_368__53_,r_368__52_,
  r_368__51_,r_368__50_,r_368__49_,r_368__48_,r_368__47_,r_368__46_,r_368__45_,
  r_368__44_,r_368__43_,r_368__42_,r_368__41_,r_368__40_,r_368__39_,r_368__38_,
  r_368__37_,r_368__36_,r_368__35_,r_368__34_,r_368__33_,r_368__32_,r_368__31_,r_368__30_,
  r_368__29_,r_368__28_,r_368__27_,r_368__26_,r_368__25_,r_368__24_,r_368__23_,
  r_368__22_,r_368__21_,r_368__20_,r_368__19_,r_368__18_,r_368__17_,r_368__16_,
  r_368__15_,r_368__14_,r_368__13_,r_368__12_,r_368__11_,r_368__10_,r_368__9_,r_368__8_,
  r_368__7_,r_368__6_,r_368__5_,r_368__4_,r_368__3_,r_368__2_,r_368__1_,r_368__0_,
  r_369__63_,r_369__62_,r_369__61_,r_369__60_,r_369__59_,r_369__58_,r_369__57_,
  r_369__56_,r_369__55_,r_369__54_,r_369__53_,r_369__52_,r_369__51_,r_369__50_,
  r_369__49_,r_369__48_,r_369__47_,r_369__46_,r_369__45_,r_369__44_,r_369__43_,
  r_369__42_,r_369__41_,r_369__40_,r_369__39_,r_369__38_,r_369__37_,r_369__36_,r_369__35_,
  r_369__34_,r_369__33_,r_369__32_,r_369__31_,r_369__30_,r_369__29_,r_369__28_,
  r_369__27_,r_369__26_,r_369__25_,r_369__24_,r_369__23_,r_369__22_,r_369__21_,
  r_369__20_,r_369__19_,r_369__18_,r_369__17_,r_369__16_,r_369__15_,r_369__14_,
  r_369__13_,r_369__12_,r_369__11_,r_369__10_,r_369__9_,r_369__8_,r_369__7_,r_369__6_,
  r_369__5_,r_369__4_,r_369__3_,r_369__2_,r_369__1_,r_369__0_,r_370__63_,r_370__62_,
  r_370__61_,r_370__60_,r_370__59_,r_370__58_,r_370__57_,r_370__56_,r_370__55_,
  r_370__54_,r_370__53_,r_370__52_,r_370__51_,r_370__50_,r_370__49_,r_370__48_,
  r_370__47_,r_370__46_,r_370__45_,r_370__44_,r_370__43_,r_370__42_,r_370__41_,r_370__40_,
  r_370__39_,r_370__38_,r_370__37_,r_370__36_,r_370__35_,r_370__34_,r_370__33_,
  r_370__32_,r_370__31_,r_370__30_,r_370__29_,r_370__28_,r_370__27_,r_370__26_,
  r_370__25_,r_370__24_,r_370__23_,r_370__22_,r_370__21_,r_370__20_,r_370__19_,r_370__18_,
  r_370__17_,r_370__16_,r_370__15_,r_370__14_,r_370__13_,r_370__12_,r_370__11_,
  r_370__10_,r_370__9_,r_370__8_,r_370__7_,r_370__6_,r_370__5_,r_370__4_,r_370__3_,
  r_370__2_,r_370__1_,r_370__0_,r_371__63_,r_371__62_,r_371__61_,r_371__60_,
  r_371__59_,r_371__58_,r_371__57_,r_371__56_,r_371__55_,r_371__54_,r_371__53_,r_371__52_,
  r_371__51_,r_371__50_,r_371__49_,r_371__48_,r_371__47_,r_371__46_,r_371__45_,
  r_371__44_,r_371__43_,r_371__42_,r_371__41_,r_371__40_,r_371__39_,r_371__38_,
  r_371__37_,r_371__36_,r_371__35_,r_371__34_,r_371__33_,r_371__32_,r_371__31_,
  r_371__30_,r_371__29_,r_371__28_,r_371__27_,r_371__26_,r_371__25_,r_371__24_,r_371__23_,
  r_371__22_,r_371__21_,r_371__20_,r_371__19_,r_371__18_,r_371__17_,r_371__16_,
  r_371__15_,r_371__14_,r_371__13_,r_371__12_,r_371__11_,r_371__10_,r_371__9_,
  r_371__8_,r_371__7_,r_371__6_,r_371__5_,r_371__4_,r_371__3_,r_371__2_,r_371__1_,
  r_371__0_,r_372__63_,r_372__62_,r_372__61_,r_372__60_,r_372__59_,r_372__58_,r_372__57_,
  r_372__56_,r_372__55_,r_372__54_,r_372__53_,r_372__52_,r_372__51_,r_372__50_,
  r_372__49_,r_372__48_,r_372__47_,r_372__46_,r_372__45_,r_372__44_,r_372__43_,
  r_372__42_,r_372__41_,r_372__40_,r_372__39_,r_372__38_,r_372__37_,r_372__36_,
  r_372__35_,r_372__34_,r_372__33_,r_372__32_,r_372__31_,r_372__30_,r_372__29_,r_372__28_,
  r_372__27_,r_372__26_,r_372__25_,r_372__24_,r_372__23_,r_372__22_,r_372__21_,
  r_372__20_,r_372__19_,r_372__18_,r_372__17_,r_372__16_,r_372__15_,r_372__14_,
  r_372__13_,r_372__12_,r_372__11_,r_372__10_,r_372__9_,r_372__8_,r_372__7_,r_372__6_,
  r_372__5_,r_372__4_,r_372__3_,r_372__2_,r_372__1_,r_372__0_,r_373__63_,r_373__62_,
  r_373__61_,r_373__60_,r_373__59_,r_373__58_,r_373__57_,r_373__56_,r_373__55_,
  r_373__54_,r_373__53_,r_373__52_,r_373__51_,r_373__50_,r_373__49_,r_373__48_,
  r_373__47_,r_373__46_,r_373__45_,r_373__44_,r_373__43_,r_373__42_,r_373__41_,r_373__40_,
  r_373__39_,r_373__38_,r_373__37_,r_373__36_,r_373__35_,r_373__34_,r_373__33_,
  r_373__32_,r_373__31_,r_373__30_,r_373__29_,r_373__28_,r_373__27_,r_373__26_,
  r_373__25_,r_373__24_,r_373__23_,r_373__22_,r_373__21_,r_373__20_,r_373__19_,
  r_373__18_,r_373__17_,r_373__16_,r_373__15_,r_373__14_,r_373__13_,r_373__12_,r_373__11_,
  r_373__10_,r_373__9_,r_373__8_,r_373__7_,r_373__6_,r_373__5_,r_373__4_,r_373__3_,
  r_373__2_,r_373__1_,r_373__0_,r_374__63_,r_374__62_,r_374__61_,r_374__60_,
  r_374__59_,r_374__58_,r_374__57_,r_374__56_,r_374__55_,r_374__54_,r_374__53_,
  r_374__52_,r_374__51_,r_374__50_,r_374__49_,r_374__48_,r_374__47_,r_374__46_,r_374__45_,
  r_374__44_,r_374__43_,r_374__42_,r_374__41_,r_374__40_,r_374__39_,r_374__38_,
  r_374__37_,r_374__36_,r_374__35_,r_374__34_,r_374__33_,r_374__32_,r_374__31_,
  r_374__30_,r_374__29_,r_374__28_,r_374__27_,r_374__26_,r_374__25_,r_374__24_,
  r_374__23_,r_374__22_,r_374__21_,r_374__20_,r_374__19_,r_374__18_,r_374__17_,r_374__16_,
  r_374__15_,r_374__14_,r_374__13_,r_374__12_,r_374__11_,r_374__10_,r_374__9_,
  r_374__8_,r_374__7_,r_374__6_,r_374__5_,r_374__4_,r_374__3_,r_374__2_,r_374__1_,
  r_374__0_,r_375__63_,r_375__62_,r_375__61_,r_375__60_,r_375__59_,r_375__58_,
  r_375__57_,r_375__56_,r_375__55_,r_375__54_,r_375__53_,r_375__52_,r_375__51_,r_375__50_,
  r_375__49_,r_375__48_,r_375__47_,r_375__46_,r_375__45_,r_375__44_,r_375__43_,
  r_375__42_,r_375__41_,r_375__40_,r_375__39_,r_375__38_,r_375__37_,r_375__36_,
  r_375__35_,r_375__34_,r_375__33_,r_375__32_,r_375__31_,r_375__30_,r_375__29_,r_375__28_,
  r_375__27_,r_375__26_,r_375__25_,r_375__24_,r_375__23_,r_375__22_,r_375__21_,
  r_375__20_,r_375__19_,r_375__18_,r_375__17_,r_375__16_,r_375__15_,r_375__14_,
  r_375__13_,r_375__12_,r_375__11_,r_375__10_,r_375__9_,r_375__8_,r_375__7_,r_375__6_,
  r_375__5_,r_375__4_,r_375__3_,r_375__2_,r_375__1_,r_375__0_,r_376__63_,r_376__62_,
  r_376__61_,r_376__60_,r_376__59_,r_376__58_,r_376__57_,r_376__56_,r_376__55_,
  r_376__54_,r_376__53_,r_376__52_,r_376__51_,r_376__50_,r_376__49_,r_376__48_,
  r_376__47_,r_376__46_,r_376__45_,r_376__44_,r_376__43_,r_376__42_,r_376__41_,
  r_376__40_,r_376__39_,r_376__38_,r_376__37_,r_376__36_,r_376__35_,r_376__34_,r_376__33_,
  r_376__32_,r_376__31_,r_376__30_,r_376__29_,r_376__28_,r_376__27_,r_376__26_,
  r_376__25_,r_376__24_,r_376__23_,r_376__22_,r_376__21_,r_376__20_,r_376__19_,
  r_376__18_,r_376__17_,r_376__16_,r_376__15_,r_376__14_,r_376__13_,r_376__12_,
  r_376__11_,r_376__10_,r_376__9_,r_376__8_,r_376__7_,r_376__6_,r_376__5_,r_376__4_,
  r_376__3_,r_376__2_,r_376__1_,r_376__0_,r_377__63_,r_377__62_,r_377__61_,r_377__60_,
  r_377__59_,r_377__58_,r_377__57_,r_377__56_,r_377__55_,r_377__54_,r_377__53_,
  r_377__52_,r_377__51_,r_377__50_,r_377__49_,r_377__48_,r_377__47_,r_377__46_,
  r_377__45_,r_377__44_,r_377__43_,r_377__42_,r_377__41_,r_377__40_,r_377__39_,r_377__38_,
  r_377__37_,r_377__36_,r_377__35_,r_377__34_,r_377__33_,r_377__32_,r_377__31_,
  r_377__30_,r_377__29_,r_377__28_,r_377__27_,r_377__26_,r_377__25_,r_377__24_,
  r_377__23_,r_377__22_,r_377__21_,r_377__20_,r_377__19_,r_377__18_,r_377__17_,r_377__16_,
  r_377__15_,r_377__14_,r_377__13_,r_377__12_,r_377__11_,r_377__10_,r_377__9_,
  r_377__8_,r_377__7_,r_377__6_,r_377__5_,r_377__4_,r_377__3_,r_377__2_,r_377__1_,
  r_377__0_,r_378__63_,r_378__62_,r_378__61_,r_378__60_,r_378__59_,r_378__58_,
  r_378__57_,r_378__56_,r_378__55_,r_378__54_,r_378__53_,r_378__52_,r_378__51_,r_378__50_,
  r_378__49_,r_378__48_,r_378__47_,r_378__46_,r_378__45_,r_378__44_,r_378__43_,
  r_378__42_,r_378__41_,r_378__40_,r_378__39_,r_378__38_,r_378__37_,r_378__36_,
  r_378__35_,r_378__34_,r_378__33_,r_378__32_,r_378__31_,r_378__30_,r_378__29_,
  r_378__28_,r_378__27_,r_378__26_,r_378__25_,r_378__24_,r_378__23_,r_378__22_,r_378__21_,
  r_378__20_,r_378__19_,r_378__18_,r_378__17_,r_378__16_,r_378__15_,r_378__14_,
  r_378__13_,r_378__12_,r_378__11_,r_378__10_,r_378__9_,r_378__8_,r_378__7_,r_378__6_,
  r_378__5_,r_378__4_,r_378__3_,r_378__2_,r_378__1_,r_378__0_,r_379__63_,
  r_379__62_,r_379__61_,r_379__60_,r_379__59_,r_379__58_,r_379__57_,r_379__56_,r_379__55_,
  r_379__54_,r_379__53_,r_379__52_,r_379__51_,r_379__50_,r_379__49_,r_379__48_,
  r_379__47_,r_379__46_,r_379__45_,r_379__44_,r_379__43_,r_379__42_,r_379__41_,
  r_379__40_,r_379__39_,r_379__38_,r_379__37_,r_379__36_,r_379__35_,r_379__34_,
  r_379__33_,r_379__32_,r_379__31_,r_379__30_,r_379__29_,r_379__28_,r_379__27_,r_379__26_,
  r_379__25_,r_379__24_,r_379__23_,r_379__22_,r_379__21_,r_379__20_,r_379__19_,
  r_379__18_,r_379__17_,r_379__16_,r_379__15_,r_379__14_,r_379__13_,r_379__12_,
  r_379__11_,r_379__10_,r_379__9_,r_379__8_,r_379__7_,r_379__6_,r_379__5_,r_379__4_,
  r_379__3_,r_379__2_,r_379__1_,r_379__0_,r_380__63_,r_380__62_,r_380__61_,r_380__60_,
  r_380__59_,r_380__58_,r_380__57_,r_380__56_,r_380__55_,r_380__54_,r_380__53_,
  r_380__52_,r_380__51_,r_380__50_,r_380__49_,r_380__48_,r_380__47_,r_380__46_,
  r_380__45_,r_380__44_,r_380__43_,r_380__42_,r_380__41_,r_380__40_,r_380__39_,r_380__38_,
  r_380__37_,r_380__36_,r_380__35_,r_380__34_,r_380__33_,r_380__32_,r_380__31_,
  r_380__30_,r_380__29_,r_380__28_,r_380__27_,r_380__26_,r_380__25_,r_380__24_,
  r_380__23_,r_380__22_,r_380__21_,r_380__20_,r_380__19_,r_380__18_,r_380__17_,
  r_380__16_,r_380__15_,r_380__14_,r_380__13_,r_380__12_,r_380__11_,r_380__10_,r_380__9_,
  r_380__8_,r_380__7_,r_380__6_,r_380__5_,r_380__4_,r_380__3_,r_380__2_,r_380__1_,
  r_380__0_,r_381__63_,r_381__62_,r_381__61_,r_381__60_,r_381__59_,r_381__58_,
  r_381__57_,r_381__56_,r_381__55_,r_381__54_,r_381__53_,r_381__52_,r_381__51_,
  r_381__50_,r_381__49_,r_381__48_,r_381__47_,r_381__46_,r_381__45_,r_381__44_,r_381__43_,
  r_381__42_,r_381__41_,r_381__40_,r_381__39_,r_381__38_,r_381__37_,r_381__36_,
  r_381__35_,r_381__34_,r_381__33_,r_381__32_,r_381__31_,r_381__30_,r_381__29_,
  r_381__28_,r_381__27_,r_381__26_,r_381__25_,r_381__24_,r_381__23_,r_381__22_,
  r_381__21_,r_381__20_,r_381__19_,r_381__18_,r_381__17_,r_381__16_,r_381__15_,r_381__14_,
  r_381__13_,r_381__12_,r_381__11_,r_381__10_,r_381__9_,r_381__8_,r_381__7_,
  r_381__6_,r_381__5_,r_381__4_,r_381__3_,r_381__2_,r_381__1_,r_381__0_,r_382__63_,
  r_382__62_,r_382__61_,r_382__60_,r_382__59_,r_382__58_,r_382__57_,r_382__56_,
  r_382__55_,r_382__54_,r_382__53_,r_382__52_,r_382__51_,r_382__50_,r_382__49_,r_382__48_,
  r_382__47_,r_382__46_,r_382__45_,r_382__44_,r_382__43_,r_382__42_,r_382__41_,
  r_382__40_,r_382__39_,r_382__38_,r_382__37_,r_382__36_,r_382__35_,r_382__34_,
  r_382__33_,r_382__32_,r_382__31_,r_382__30_,r_382__29_,r_382__28_,r_382__27_,r_382__26_,
  r_382__25_,r_382__24_,r_382__23_,r_382__22_,r_382__21_,r_382__20_,r_382__19_,
  r_382__18_,r_382__17_,r_382__16_,r_382__15_,r_382__14_,r_382__13_,r_382__12_,
  r_382__11_,r_382__10_,r_382__9_,r_382__8_,r_382__7_,r_382__6_,r_382__5_,r_382__4_,
  r_382__3_,r_382__2_,r_382__1_,r_382__0_,r_383__63_,r_383__62_,r_383__61_,r_383__60_,
  r_383__59_,r_383__58_,r_383__57_,r_383__56_,r_383__55_,r_383__54_,r_383__53_,
  r_383__52_,r_383__51_,r_383__50_,r_383__49_,r_383__48_,r_383__47_,r_383__46_,
  r_383__45_,r_383__44_,r_383__43_,r_383__42_,r_383__41_,r_383__40_,r_383__39_,
  r_383__38_,r_383__37_,r_383__36_,r_383__35_,r_383__34_,r_383__33_,r_383__32_,r_383__31_,
  r_383__30_,r_383__29_,r_383__28_,r_383__27_,r_383__26_,r_383__25_,r_383__24_,
  r_383__23_,r_383__22_,r_383__21_,r_383__20_,r_383__19_,r_383__18_,r_383__17_,
  r_383__16_,r_383__15_,r_383__14_,r_383__13_,r_383__12_,r_383__11_,r_383__10_,r_383__9_,
  r_383__8_,r_383__7_,r_383__6_,r_383__5_,r_383__4_,r_383__3_,r_383__2_,r_383__1_,
  r_383__0_,r_384__63_,r_384__62_,r_384__61_,r_384__60_,r_384__59_,r_384__58_,
  r_384__57_,r_384__56_,r_384__55_,r_384__54_,r_384__53_,r_384__52_,r_384__51_,
  r_384__50_,r_384__49_,r_384__48_,r_384__47_,r_384__46_,r_384__45_,r_384__44_,
  r_384__43_,r_384__42_,r_384__41_,r_384__40_,r_384__39_,r_384__38_,r_384__37_,r_384__36_,
  r_384__35_,r_384__34_,r_384__33_,r_384__32_,r_384__31_,r_384__30_,r_384__29_,
  r_384__28_,r_384__27_,r_384__26_,r_384__25_,r_384__24_,r_384__23_,r_384__22_,
  r_384__21_,r_384__20_,r_384__19_,r_384__18_,r_384__17_,r_384__16_,r_384__15_,r_384__14_,
  r_384__13_,r_384__12_,r_384__11_,r_384__10_,r_384__9_,r_384__8_,r_384__7_,
  r_384__6_,r_384__5_,r_384__4_,r_384__3_,r_384__2_,r_384__1_,r_384__0_,r_385__63_,
  r_385__62_,r_385__61_,r_385__60_,r_385__59_,r_385__58_,r_385__57_,r_385__56_,
  r_385__55_,r_385__54_,r_385__53_,r_385__52_,r_385__51_,r_385__50_,r_385__49_,r_385__48_,
  r_385__47_,r_385__46_,r_385__45_,r_385__44_,r_385__43_,r_385__42_,r_385__41_,
  r_385__40_,r_385__39_,r_385__38_,r_385__37_,r_385__36_,r_385__35_,r_385__34_,
  r_385__33_,r_385__32_,r_385__31_,r_385__30_,r_385__29_,r_385__28_,r_385__27_,
  r_385__26_,r_385__25_,r_385__24_,r_385__23_,r_385__22_,r_385__21_,r_385__20_,r_385__19_,
  r_385__18_,r_385__17_,r_385__16_,r_385__15_,r_385__14_,r_385__13_,r_385__12_,
  r_385__11_,r_385__10_,r_385__9_,r_385__8_,r_385__7_,r_385__6_,r_385__5_,r_385__4_,
  r_385__3_,r_385__2_,r_385__1_,r_385__0_,r_386__63_,r_386__62_,r_386__61_,
  r_386__60_,r_386__59_,r_386__58_,r_386__57_,r_386__56_,r_386__55_,r_386__54_,r_386__53_,
  r_386__52_,r_386__51_,r_386__50_,r_386__49_,r_386__48_,r_386__47_,r_386__46_,
  r_386__45_,r_386__44_,r_386__43_,r_386__42_,r_386__41_,r_386__40_,r_386__39_,
  r_386__38_,r_386__37_,r_386__36_,r_386__35_,r_386__34_,r_386__33_,r_386__32_,
  r_386__31_,r_386__30_,r_386__29_,r_386__28_,r_386__27_,r_386__26_,r_386__25_,r_386__24_,
  r_386__23_,r_386__22_,r_386__21_,r_386__20_,r_386__19_,r_386__18_,r_386__17_,
  r_386__16_,r_386__15_,r_386__14_,r_386__13_,r_386__12_,r_386__11_,r_386__10_,
  r_386__9_,r_386__8_,r_386__7_,r_386__6_,r_386__5_,r_386__4_,r_386__3_,r_386__2_,
  r_386__1_,r_386__0_,r_387__63_,r_387__62_,r_387__61_,r_387__60_,r_387__59_,r_387__58_,
  r_387__57_,r_387__56_,r_387__55_,r_387__54_,r_387__53_,r_387__52_,r_387__51_,
  r_387__50_,r_387__49_,r_387__48_,r_387__47_,r_387__46_,r_387__45_,r_387__44_,
  r_387__43_,r_387__42_,r_387__41_,r_387__40_,r_387__39_,r_387__38_,r_387__37_,r_387__36_,
  r_387__35_,r_387__34_,r_387__33_,r_387__32_,r_387__31_,r_387__30_,r_387__29_,
  r_387__28_,r_387__27_,r_387__26_,r_387__25_,r_387__24_,r_387__23_,r_387__22_,
  r_387__21_,r_387__20_,r_387__19_,r_387__18_,r_387__17_,r_387__16_,r_387__15_,
  r_387__14_,r_387__13_,r_387__12_,r_387__11_,r_387__10_,r_387__9_,r_387__8_,r_387__7_,
  r_387__6_,r_387__5_,r_387__4_,r_387__3_,r_387__2_,r_387__1_,r_387__0_,r_388__63_,
  r_388__62_,r_388__61_,r_388__60_,r_388__59_,r_388__58_,r_388__57_,r_388__56_,
  r_388__55_,r_388__54_,r_388__53_,r_388__52_,r_388__51_,r_388__50_,r_388__49_,
  r_388__48_,r_388__47_,r_388__46_,r_388__45_,r_388__44_,r_388__43_,r_388__42_,r_388__41_,
  r_388__40_,r_388__39_,r_388__38_,r_388__37_,r_388__36_,r_388__35_,r_388__34_,
  r_388__33_,r_388__32_,r_388__31_,r_388__30_,r_388__29_,r_388__28_,r_388__27_,
  r_388__26_,r_388__25_,r_388__24_,r_388__23_,r_388__22_,r_388__21_,r_388__20_,
  r_388__19_,r_388__18_,r_388__17_,r_388__16_,r_388__15_,r_388__14_,r_388__13_,r_388__12_,
  r_388__11_,r_388__10_,r_388__9_,r_388__8_,r_388__7_,r_388__6_,r_388__5_,r_388__4_,
  r_388__3_,r_388__2_,r_388__1_,r_388__0_,r_389__63_,r_389__62_,r_389__61_,
  r_389__60_,r_389__59_,r_389__58_,r_389__57_,r_389__56_,r_389__55_,r_389__54_,
  r_389__53_,r_389__52_,r_389__51_,r_389__50_,r_389__49_,r_389__48_,r_389__47_,r_389__46_,
  r_389__45_,r_389__44_,r_389__43_,r_389__42_,r_389__41_,r_389__40_,r_389__39_,
  r_389__38_,r_389__37_,r_389__36_,r_389__35_,r_389__34_,r_389__33_,r_389__32_,
  r_389__31_,r_389__30_,r_389__29_,r_389__28_,r_389__27_,r_389__26_,r_389__25_,r_389__24_,
  r_389__23_,r_389__22_,r_389__21_,r_389__20_,r_389__19_,r_389__18_,r_389__17_,
  r_389__16_,r_389__15_,r_389__14_,r_389__13_,r_389__12_,r_389__11_,r_389__10_,
  r_389__9_,r_389__8_,r_389__7_,r_389__6_,r_389__5_,r_389__4_,r_389__3_,r_389__2_,
  r_389__1_,r_389__0_,r_390__63_,r_390__62_,r_390__61_,r_390__60_,r_390__59_,r_390__58_,
  r_390__57_,r_390__56_,r_390__55_,r_390__54_,r_390__53_,r_390__52_,r_390__51_,
  r_390__50_,r_390__49_,r_390__48_,r_390__47_,r_390__46_,r_390__45_,r_390__44_,
  r_390__43_,r_390__42_,r_390__41_,r_390__40_,r_390__39_,r_390__38_,r_390__37_,
  r_390__36_,r_390__35_,r_390__34_,r_390__33_,r_390__32_,r_390__31_,r_390__30_,r_390__29_,
  r_390__28_,r_390__27_,r_390__26_,r_390__25_,r_390__24_,r_390__23_,r_390__22_,
  r_390__21_,r_390__20_,r_390__19_,r_390__18_,r_390__17_,r_390__16_,r_390__15_,
  r_390__14_,r_390__13_,r_390__12_,r_390__11_,r_390__10_,r_390__9_,r_390__8_,r_390__7_,
  r_390__6_,r_390__5_,r_390__4_,r_390__3_,r_390__2_,r_390__1_,r_390__0_,r_391__63_,
  r_391__62_,r_391__61_,r_391__60_,r_391__59_,r_391__58_,r_391__57_,r_391__56_,
  r_391__55_,r_391__54_,r_391__53_,r_391__52_,r_391__51_,r_391__50_,r_391__49_,
  r_391__48_,r_391__47_,r_391__46_,r_391__45_,r_391__44_,r_391__43_,r_391__42_,
  r_391__41_,r_391__40_,r_391__39_,r_391__38_,r_391__37_,r_391__36_,r_391__35_,r_391__34_,
  r_391__33_,r_391__32_,r_391__31_,r_391__30_,r_391__29_,r_391__28_,r_391__27_,
  r_391__26_,r_391__25_,r_391__24_,r_391__23_,r_391__22_,r_391__21_,r_391__20_,
  r_391__19_,r_391__18_,r_391__17_,r_391__16_,r_391__15_,r_391__14_,r_391__13_,r_391__12_,
  r_391__11_,r_391__10_,r_391__9_,r_391__8_,r_391__7_,r_391__6_,r_391__5_,
  r_391__4_,r_391__3_,r_391__2_,r_391__1_,r_391__0_,r_392__63_,r_392__62_,r_392__61_,
  r_392__60_,r_392__59_,r_392__58_,r_392__57_,r_392__56_,r_392__55_,r_392__54_,
  r_392__53_,r_392__52_,r_392__51_,r_392__50_,r_392__49_,r_392__48_,r_392__47_,r_392__46_,
  r_392__45_,r_392__44_,r_392__43_,r_392__42_,r_392__41_,r_392__40_,r_392__39_,
  r_392__38_,r_392__37_,r_392__36_,r_392__35_,r_392__34_,r_392__33_,r_392__32_,
  r_392__31_,r_392__30_,r_392__29_,r_392__28_,r_392__27_,r_392__26_,r_392__25_,
  r_392__24_,r_392__23_,r_392__22_,r_392__21_,r_392__20_,r_392__19_,r_392__18_,r_392__17_,
  r_392__16_,r_392__15_,r_392__14_,r_392__13_,r_392__12_,r_392__11_,r_392__10_,
  r_392__9_,r_392__8_,r_392__7_,r_392__6_,r_392__5_,r_392__4_,r_392__3_,r_392__2_,
  r_392__1_,r_392__0_,r_393__63_,r_393__62_,r_393__61_,r_393__60_,r_393__59_,
  r_393__58_,r_393__57_,r_393__56_,r_393__55_,r_393__54_,r_393__53_,r_393__52_,r_393__51_,
  r_393__50_,r_393__49_,r_393__48_,r_393__47_,r_393__46_,r_393__45_,r_393__44_,
  r_393__43_,r_393__42_,r_393__41_,r_393__40_,r_393__39_,r_393__38_,r_393__37_,
  r_393__36_,r_393__35_,r_393__34_,r_393__33_,r_393__32_,r_393__31_,r_393__30_,
  r_393__29_,r_393__28_,r_393__27_,r_393__26_,r_393__25_,r_393__24_,r_393__23_,r_393__22_,
  r_393__21_,r_393__20_,r_393__19_,r_393__18_,r_393__17_,r_393__16_,r_393__15_,
  r_393__14_,r_393__13_,r_393__12_,r_393__11_,r_393__10_,r_393__9_,r_393__8_,r_393__7_,
  r_393__6_,r_393__5_,r_393__4_,r_393__3_,r_393__2_,r_393__1_,r_393__0_,
  r_394__63_,r_394__62_,r_394__61_,r_394__60_,r_394__59_,r_394__58_,r_394__57_,r_394__56_,
  r_394__55_,r_394__54_,r_394__53_,r_394__52_,r_394__51_,r_394__50_,r_394__49_,
  r_394__48_,r_394__47_,r_394__46_,r_394__45_,r_394__44_,r_394__43_,r_394__42_,
  r_394__41_,r_394__40_,r_394__39_,r_394__38_,r_394__37_,r_394__36_,r_394__35_,r_394__34_,
  r_394__33_,r_394__32_,r_394__31_,r_394__30_,r_394__29_,r_394__28_,r_394__27_,
  r_394__26_,r_394__25_,r_394__24_,r_394__23_,r_394__22_,r_394__21_,r_394__20_,
  r_394__19_,r_394__18_,r_394__17_,r_394__16_,r_394__15_,r_394__14_,r_394__13_,
  r_394__12_,r_394__11_,r_394__10_,r_394__9_,r_394__8_,r_394__7_,r_394__6_,r_394__5_,
  r_394__4_,r_394__3_,r_394__2_,r_394__1_,r_394__0_,r_395__63_,r_395__62_,r_395__61_,
  r_395__60_,r_395__59_,r_395__58_,r_395__57_,r_395__56_,r_395__55_,r_395__54_,
  r_395__53_,r_395__52_,r_395__51_,r_395__50_,r_395__49_,r_395__48_,r_395__47_,
  r_395__46_,r_395__45_,r_395__44_,r_395__43_,r_395__42_,r_395__41_,r_395__40_,r_395__39_,
  r_395__38_,r_395__37_,r_395__36_,r_395__35_,r_395__34_,r_395__33_,r_395__32_,
  r_395__31_,r_395__30_,r_395__29_,r_395__28_,r_395__27_,r_395__26_,r_395__25_,
  r_395__24_,r_395__23_,r_395__22_,r_395__21_,r_395__20_,r_395__19_,r_395__18_,
  r_395__17_,r_395__16_,r_395__15_,r_395__14_,r_395__13_,r_395__12_,r_395__11_,r_395__10_,
  r_395__9_,r_395__8_,r_395__7_,r_395__6_,r_395__5_,r_395__4_,r_395__3_,r_395__2_,
  r_395__1_,r_395__0_,r_396__63_,r_396__62_,r_396__61_,r_396__60_,r_396__59_,
  r_396__58_,r_396__57_,r_396__56_,r_396__55_,r_396__54_,r_396__53_,r_396__52_,
  r_396__51_,r_396__50_,r_396__49_,r_396__48_,r_396__47_,r_396__46_,r_396__45_,r_396__44_,
  r_396__43_,r_396__42_,r_396__41_,r_396__40_,r_396__39_,r_396__38_,r_396__37_,
  r_396__36_,r_396__35_,r_396__34_,r_396__33_,r_396__32_,r_396__31_,r_396__30_,
  r_396__29_,r_396__28_,r_396__27_,r_396__26_,r_396__25_,r_396__24_,r_396__23_,r_396__22_,
  r_396__21_,r_396__20_,r_396__19_,r_396__18_,r_396__17_,r_396__16_,r_396__15_,
  r_396__14_,r_396__13_,r_396__12_,r_396__11_,r_396__10_,r_396__9_,r_396__8_,
  r_396__7_,r_396__6_,r_396__5_,r_396__4_,r_396__3_,r_396__2_,r_396__1_,r_396__0_,
  r_397__63_,r_397__62_,r_397__61_,r_397__60_,r_397__59_,r_397__58_,r_397__57_,r_397__56_,
  r_397__55_,r_397__54_,r_397__53_,r_397__52_,r_397__51_,r_397__50_,r_397__49_,
  r_397__48_,r_397__47_,r_397__46_,r_397__45_,r_397__44_,r_397__43_,r_397__42_,
  r_397__41_,r_397__40_,r_397__39_,r_397__38_,r_397__37_,r_397__36_,r_397__35_,
  r_397__34_,r_397__33_,r_397__32_,r_397__31_,r_397__30_,r_397__29_,r_397__28_,r_397__27_,
  r_397__26_,r_397__25_,r_397__24_,r_397__23_,r_397__22_,r_397__21_,r_397__20_,
  r_397__19_,r_397__18_,r_397__17_,r_397__16_,r_397__15_,r_397__14_,r_397__13_,
  r_397__12_,r_397__11_,r_397__10_,r_397__9_,r_397__8_,r_397__7_,r_397__6_,r_397__5_,
  r_397__4_,r_397__3_,r_397__2_,r_397__1_,r_397__0_,r_398__63_,r_398__62_,r_398__61_,
  r_398__60_,r_398__59_,r_398__58_,r_398__57_,r_398__56_,r_398__55_,r_398__54_,
  r_398__53_,r_398__52_,r_398__51_,r_398__50_,r_398__49_,r_398__48_,r_398__47_,
  r_398__46_,r_398__45_,r_398__44_,r_398__43_,r_398__42_,r_398__41_,r_398__40_,
  r_398__39_,r_398__38_,r_398__37_,r_398__36_,r_398__35_,r_398__34_,r_398__33_,r_398__32_,
  r_398__31_,r_398__30_,r_398__29_,r_398__28_,r_398__27_,r_398__26_,r_398__25_,
  r_398__24_,r_398__23_,r_398__22_,r_398__21_,r_398__20_,r_398__19_,r_398__18_,
  r_398__17_,r_398__16_,r_398__15_,r_398__14_,r_398__13_,r_398__12_,r_398__11_,r_398__10_,
  r_398__9_,r_398__8_,r_398__7_,r_398__6_,r_398__5_,r_398__4_,r_398__3_,r_398__2_,
  r_398__1_,r_398__0_,r_399__63_,r_399__62_,r_399__61_,r_399__60_,r_399__59_,
  r_399__58_,r_399__57_,r_399__56_,r_399__55_,r_399__54_,r_399__53_,r_399__52_,
  r_399__51_,r_399__50_,r_399__49_,r_399__48_,r_399__47_,r_399__46_,r_399__45_,r_399__44_,
  r_399__43_,r_399__42_,r_399__41_,r_399__40_,r_399__39_,r_399__38_,r_399__37_,
  r_399__36_,r_399__35_,r_399__34_,r_399__33_,r_399__32_,r_399__31_,r_399__30_,
  r_399__29_,r_399__28_,r_399__27_,r_399__26_,r_399__25_,r_399__24_,r_399__23_,
  r_399__22_,r_399__21_,r_399__20_,r_399__19_,r_399__18_,r_399__17_,r_399__16_,r_399__15_,
  r_399__14_,r_399__13_,r_399__12_,r_399__11_,r_399__10_,r_399__9_,r_399__8_,
  r_399__7_,r_399__6_,r_399__5_,r_399__4_,r_399__3_,r_399__2_,r_399__1_,r_399__0_,
  r_400__63_,r_400__62_,r_400__61_,r_400__60_,r_400__59_,r_400__58_,r_400__57_,
  r_400__56_,r_400__55_,r_400__54_,r_400__53_,r_400__52_,r_400__51_,r_400__50_,r_400__49_,
  r_400__48_,r_400__47_,r_400__46_,r_400__45_,r_400__44_,r_400__43_,r_400__42_,
  r_400__41_,r_400__40_,r_400__39_,r_400__38_,r_400__37_,r_400__36_,r_400__35_,
  r_400__34_,r_400__33_,r_400__32_,r_400__31_,r_400__30_,r_400__29_,r_400__28_,
  r_400__27_,r_400__26_,r_400__25_,r_400__24_,r_400__23_,r_400__22_,r_400__21_,r_400__20_,
  r_400__19_,r_400__18_,r_400__17_,r_400__16_,r_400__15_,r_400__14_,r_400__13_,
  r_400__12_,r_400__11_,r_400__10_,r_400__9_,r_400__8_,r_400__7_,r_400__6_,r_400__5_,
  r_400__4_,r_400__3_,r_400__2_,r_400__1_,r_400__0_,r_401__63_,r_401__62_,
  r_401__61_,r_401__60_,r_401__59_,r_401__58_,r_401__57_,r_401__56_,r_401__55_,r_401__54_,
  r_401__53_,r_401__52_,r_401__51_,r_401__50_,r_401__49_,r_401__48_,r_401__47_,
  r_401__46_,r_401__45_,r_401__44_,r_401__43_,r_401__42_,r_401__41_,r_401__40_,
  r_401__39_,r_401__38_,r_401__37_,r_401__36_,r_401__35_,r_401__34_,r_401__33_,r_401__32_,
  r_401__31_,r_401__30_,r_401__29_,r_401__28_,r_401__27_,r_401__26_,r_401__25_,
  r_401__24_,r_401__23_,r_401__22_,r_401__21_,r_401__20_,r_401__19_,r_401__18_,
  r_401__17_,r_401__16_,r_401__15_,r_401__14_,r_401__13_,r_401__12_,r_401__11_,
  r_401__10_,r_401__9_,r_401__8_,r_401__7_,r_401__6_,r_401__5_,r_401__4_,r_401__3_,
  r_401__2_,r_401__1_,r_401__0_,r_402__63_,r_402__62_,r_402__61_,r_402__60_,r_402__59_,
  r_402__58_,r_402__57_,r_402__56_,r_402__55_,r_402__54_,r_402__53_,r_402__52_,
  r_402__51_,r_402__50_,r_402__49_,r_402__48_,r_402__47_,r_402__46_,r_402__45_,
  r_402__44_,r_402__43_,r_402__42_,r_402__41_,r_402__40_,r_402__39_,r_402__38_,r_402__37_,
  r_402__36_,r_402__35_,r_402__34_,r_402__33_,r_402__32_,r_402__31_,r_402__30_,
  r_402__29_,r_402__28_,r_402__27_,r_402__26_,r_402__25_,r_402__24_,r_402__23_,
  r_402__22_,r_402__21_,r_402__20_,r_402__19_,r_402__18_,r_402__17_,r_402__16_,
  r_402__15_,r_402__14_,r_402__13_,r_402__12_,r_402__11_,r_402__10_,r_402__9_,r_402__8_,
  r_402__7_,r_402__6_,r_402__5_,r_402__4_,r_402__3_,r_402__2_,r_402__1_,r_402__0_,
  r_403__63_,r_403__62_,r_403__61_,r_403__60_,r_403__59_,r_403__58_,r_403__57_,
  r_403__56_,r_403__55_,r_403__54_,r_403__53_,r_403__52_,r_403__51_,r_403__50_,
  r_403__49_,r_403__48_,r_403__47_,r_403__46_,r_403__45_,r_403__44_,r_403__43_,r_403__42_,
  r_403__41_,r_403__40_,r_403__39_,r_403__38_,r_403__37_,r_403__36_,r_403__35_,
  r_403__34_,r_403__33_,r_403__32_,r_403__31_,r_403__30_,r_403__29_,r_403__28_,
  r_403__27_,r_403__26_,r_403__25_,r_403__24_,r_403__23_,r_403__22_,r_403__21_,r_403__20_,
  r_403__19_,r_403__18_,r_403__17_,r_403__16_,r_403__15_,r_403__14_,r_403__13_,
  r_403__12_,r_403__11_,r_403__10_,r_403__9_,r_403__8_,r_403__7_,r_403__6_,r_403__5_,
  r_403__4_,r_403__3_,r_403__2_,r_403__1_,r_403__0_,r_404__63_,r_404__62_,
  r_404__61_,r_404__60_,r_404__59_,r_404__58_,r_404__57_,r_404__56_,r_404__55_,r_404__54_,
  r_404__53_,r_404__52_,r_404__51_,r_404__50_,r_404__49_,r_404__48_,r_404__47_,
  r_404__46_,r_404__45_,r_404__44_,r_404__43_,r_404__42_,r_404__41_,r_404__40_,
  r_404__39_,r_404__38_,r_404__37_,r_404__36_,r_404__35_,r_404__34_,r_404__33_,
  r_404__32_,r_404__31_,r_404__30_,r_404__29_,r_404__28_,r_404__27_,r_404__26_,r_404__25_,
  r_404__24_,r_404__23_,r_404__22_,r_404__21_,r_404__20_,r_404__19_,r_404__18_,
  r_404__17_,r_404__16_,r_404__15_,r_404__14_,r_404__13_,r_404__12_,r_404__11_,
  r_404__10_,r_404__9_,r_404__8_,r_404__7_,r_404__6_,r_404__5_,r_404__4_,r_404__3_,
  r_404__2_,r_404__1_,r_404__0_,r_405__63_,r_405__62_,r_405__61_,r_405__60_,r_405__59_,
  r_405__58_,r_405__57_,r_405__56_,r_405__55_,r_405__54_,r_405__53_,r_405__52_,
  r_405__51_,r_405__50_,r_405__49_,r_405__48_,r_405__47_,r_405__46_,r_405__45_,
  r_405__44_,r_405__43_,r_405__42_,r_405__41_,r_405__40_,r_405__39_,r_405__38_,
  r_405__37_,r_405__36_,r_405__35_,r_405__34_,r_405__33_,r_405__32_,r_405__31_,r_405__30_,
  r_405__29_,r_405__28_,r_405__27_,r_405__26_,r_405__25_,r_405__24_,r_405__23_,
  r_405__22_,r_405__21_,r_405__20_,r_405__19_,r_405__18_,r_405__17_,r_405__16_,
  r_405__15_,r_405__14_,r_405__13_,r_405__12_,r_405__11_,r_405__10_,r_405__9_,r_405__8_,
  r_405__7_,r_405__6_,r_405__5_,r_405__4_,r_405__3_,r_405__2_,r_405__1_,r_405__0_,
  r_406__63_,r_406__62_,r_406__61_,r_406__60_,r_406__59_,r_406__58_,r_406__57_,
  r_406__56_,r_406__55_,r_406__54_,r_406__53_,r_406__52_,r_406__51_,r_406__50_,
  r_406__49_,r_406__48_,r_406__47_,r_406__46_,r_406__45_,r_406__44_,r_406__43_,r_406__42_,
  r_406__41_,r_406__40_,r_406__39_,r_406__38_,r_406__37_,r_406__36_,r_406__35_,
  r_406__34_,r_406__33_,r_406__32_,r_406__31_,r_406__30_,r_406__29_,r_406__28_,
  r_406__27_,r_406__26_,r_406__25_,r_406__24_,r_406__23_,r_406__22_,r_406__21_,
  r_406__20_,r_406__19_,r_406__18_,r_406__17_,r_406__16_,r_406__15_,r_406__14_,r_406__13_,
  r_406__12_,r_406__11_,r_406__10_,r_406__9_,r_406__8_,r_406__7_,r_406__6_,
  r_406__5_,r_406__4_,r_406__3_,r_406__2_,r_406__1_,r_406__0_,r_407__63_,r_407__62_,
  r_407__61_,r_407__60_,r_407__59_,r_407__58_,r_407__57_,r_407__56_,r_407__55_,
  r_407__54_,r_407__53_,r_407__52_,r_407__51_,r_407__50_,r_407__49_,r_407__48_,r_407__47_,
  r_407__46_,r_407__45_,r_407__44_,r_407__43_,r_407__42_,r_407__41_,r_407__40_,
  r_407__39_,r_407__38_,r_407__37_,r_407__36_,r_407__35_,r_407__34_,r_407__33_,
  r_407__32_,r_407__31_,r_407__30_,r_407__29_,r_407__28_,r_407__27_,r_407__26_,
  r_407__25_,r_407__24_,r_407__23_,r_407__22_,r_407__21_,r_407__20_,r_407__19_,r_407__18_,
  r_407__17_,r_407__16_,r_407__15_,r_407__14_,r_407__13_,r_407__12_,r_407__11_,
  r_407__10_,r_407__9_,r_407__8_,r_407__7_,r_407__6_,r_407__5_,r_407__4_,r_407__3_,
  r_407__2_,r_407__1_,r_407__0_,r_408__63_,r_408__62_,r_408__61_,r_408__60_,
  r_408__59_,r_408__58_,r_408__57_,r_408__56_,r_408__55_,r_408__54_,r_408__53_,r_408__52_,
  r_408__51_,r_408__50_,r_408__49_,r_408__48_,r_408__47_,r_408__46_,r_408__45_,
  r_408__44_,r_408__43_,r_408__42_,r_408__41_,r_408__40_,r_408__39_,r_408__38_,
  r_408__37_,r_408__36_,r_408__35_,r_408__34_,r_408__33_,r_408__32_,r_408__31_,r_408__30_,
  r_408__29_,r_408__28_,r_408__27_,r_408__26_,r_408__25_,r_408__24_,r_408__23_,
  r_408__22_,r_408__21_,r_408__20_,r_408__19_,r_408__18_,r_408__17_,r_408__16_,
  r_408__15_,r_408__14_,r_408__13_,r_408__12_,r_408__11_,r_408__10_,r_408__9_,r_408__8_,
  r_408__7_,r_408__6_,r_408__5_,r_408__4_,r_408__3_,r_408__2_,r_408__1_,r_408__0_,
  r_409__63_,r_409__62_,r_409__61_,r_409__60_,r_409__59_,r_409__58_,r_409__57_,
  r_409__56_,r_409__55_,r_409__54_,r_409__53_,r_409__52_,r_409__51_,r_409__50_,
  r_409__49_,r_409__48_,r_409__47_,r_409__46_,r_409__45_,r_409__44_,r_409__43_,
  r_409__42_,r_409__41_,r_409__40_,r_409__39_,r_409__38_,r_409__37_,r_409__36_,r_409__35_,
  r_409__34_,r_409__33_,r_409__32_,r_409__31_,r_409__30_,r_409__29_,r_409__28_,
  r_409__27_,r_409__26_,r_409__25_,r_409__24_,r_409__23_,r_409__22_,r_409__21_,
  r_409__20_,r_409__19_,r_409__18_,r_409__17_,r_409__16_,r_409__15_,r_409__14_,
  r_409__13_,r_409__12_,r_409__11_,r_409__10_,r_409__9_,r_409__8_,r_409__7_,r_409__6_,
  r_409__5_,r_409__4_,r_409__3_,r_409__2_,r_409__1_,r_409__0_,r_410__63_,r_410__62_,
  r_410__61_,r_410__60_,r_410__59_,r_410__58_,r_410__57_,r_410__56_,r_410__55_,
  r_410__54_,r_410__53_,r_410__52_,r_410__51_,r_410__50_,r_410__49_,r_410__48_,
  r_410__47_,r_410__46_,r_410__45_,r_410__44_,r_410__43_,r_410__42_,r_410__41_,r_410__40_,
  r_410__39_,r_410__38_,r_410__37_,r_410__36_,r_410__35_,r_410__34_,r_410__33_,
  r_410__32_,r_410__31_,r_410__30_,r_410__29_,r_410__28_,r_410__27_,r_410__26_,
  r_410__25_,r_410__24_,r_410__23_,r_410__22_,r_410__21_,r_410__20_,r_410__19_,r_410__18_,
  r_410__17_,r_410__16_,r_410__15_,r_410__14_,r_410__13_,r_410__12_,r_410__11_,
  r_410__10_,r_410__9_,r_410__8_,r_410__7_,r_410__6_,r_410__5_,r_410__4_,r_410__3_,
  r_410__2_,r_410__1_,r_410__0_,r_411__63_,r_411__62_,r_411__61_,r_411__60_,
  r_411__59_,r_411__58_,r_411__57_,r_411__56_,r_411__55_,r_411__54_,r_411__53_,r_411__52_,
  r_411__51_,r_411__50_,r_411__49_,r_411__48_,r_411__47_,r_411__46_,r_411__45_,
  r_411__44_,r_411__43_,r_411__42_,r_411__41_,r_411__40_,r_411__39_,r_411__38_,
  r_411__37_,r_411__36_,r_411__35_,r_411__34_,r_411__33_,r_411__32_,r_411__31_,
  r_411__30_,r_411__29_,r_411__28_,r_411__27_,r_411__26_,r_411__25_,r_411__24_,r_411__23_,
  r_411__22_,r_411__21_,r_411__20_,r_411__19_,r_411__18_,r_411__17_,r_411__16_,
  r_411__15_,r_411__14_,r_411__13_,r_411__12_,r_411__11_,r_411__10_,r_411__9_,
  r_411__8_,r_411__7_,r_411__6_,r_411__5_,r_411__4_,r_411__3_,r_411__2_,r_411__1_,
  r_411__0_,r_412__63_,r_412__62_,r_412__61_,r_412__60_,r_412__59_,r_412__58_,r_412__57_,
  r_412__56_,r_412__55_,r_412__54_,r_412__53_,r_412__52_,r_412__51_,r_412__50_,
  r_412__49_,r_412__48_,r_412__47_,r_412__46_,r_412__45_,r_412__44_,r_412__43_,
  r_412__42_,r_412__41_,r_412__40_,r_412__39_,r_412__38_,r_412__37_,r_412__36_,
  r_412__35_,r_412__34_,r_412__33_,r_412__32_,r_412__31_,r_412__30_,r_412__29_,r_412__28_,
  r_412__27_,r_412__26_,r_412__25_,r_412__24_,r_412__23_,r_412__22_,r_412__21_,
  r_412__20_,r_412__19_,r_412__18_,r_412__17_,r_412__16_,r_412__15_,r_412__14_,
  r_412__13_,r_412__12_,r_412__11_,r_412__10_,r_412__9_,r_412__8_,r_412__7_,r_412__6_,
  r_412__5_,r_412__4_,r_412__3_,r_412__2_,r_412__1_,r_412__0_,r_413__63_,r_413__62_,
  r_413__61_,r_413__60_,r_413__59_,r_413__58_,r_413__57_,r_413__56_,r_413__55_,
  r_413__54_,r_413__53_,r_413__52_,r_413__51_,r_413__50_,r_413__49_,r_413__48_,
  r_413__47_,r_413__46_,r_413__45_,r_413__44_,r_413__43_,r_413__42_,r_413__41_,r_413__40_,
  r_413__39_,r_413__38_,r_413__37_,r_413__36_,r_413__35_,r_413__34_,r_413__33_,
  r_413__32_,r_413__31_,r_413__30_,r_413__29_,r_413__28_,r_413__27_,r_413__26_,
  r_413__25_,r_413__24_,r_413__23_,r_413__22_,r_413__21_,r_413__20_,r_413__19_,
  r_413__18_,r_413__17_,r_413__16_,r_413__15_,r_413__14_,r_413__13_,r_413__12_,r_413__11_,
  r_413__10_,r_413__9_,r_413__8_,r_413__7_,r_413__6_,r_413__5_,r_413__4_,r_413__3_,
  r_413__2_,r_413__1_,r_413__0_,r_414__63_,r_414__62_,r_414__61_,r_414__60_,
  r_414__59_,r_414__58_,r_414__57_,r_414__56_,r_414__55_,r_414__54_,r_414__53_,
  r_414__52_,r_414__51_,r_414__50_,r_414__49_,r_414__48_,r_414__47_,r_414__46_,r_414__45_,
  r_414__44_,r_414__43_,r_414__42_,r_414__41_,r_414__40_,r_414__39_,r_414__38_,
  r_414__37_,r_414__36_,r_414__35_,r_414__34_,r_414__33_,r_414__32_,r_414__31_,
  r_414__30_,r_414__29_,r_414__28_,r_414__27_,r_414__26_,r_414__25_,r_414__24_,
  r_414__23_,r_414__22_,r_414__21_,r_414__20_,r_414__19_,r_414__18_,r_414__17_,r_414__16_,
  r_414__15_,r_414__14_,r_414__13_,r_414__12_,r_414__11_,r_414__10_,r_414__9_,
  r_414__8_,r_414__7_,r_414__6_,r_414__5_,r_414__4_,r_414__3_,r_414__2_,r_414__1_,
  r_414__0_,r_415__63_,r_415__62_,r_415__61_,r_415__60_,r_415__59_,r_415__58_,
  r_415__57_,r_415__56_,r_415__55_,r_415__54_,r_415__53_,r_415__52_,r_415__51_,r_415__50_,
  r_415__49_,r_415__48_,r_415__47_,r_415__46_,r_415__45_,r_415__44_,r_415__43_,
  r_415__42_,r_415__41_,r_415__40_,r_415__39_,r_415__38_,r_415__37_,r_415__36_,
  r_415__35_,r_415__34_,r_415__33_,r_415__32_,r_415__31_,r_415__30_,r_415__29_,r_415__28_,
  r_415__27_,r_415__26_,r_415__25_,r_415__24_,r_415__23_,r_415__22_,r_415__21_,
  r_415__20_,r_415__19_,r_415__18_,r_415__17_,r_415__16_,r_415__15_,r_415__14_,
  r_415__13_,r_415__12_,r_415__11_,r_415__10_,r_415__9_,r_415__8_,r_415__7_,r_415__6_,
  r_415__5_,r_415__4_,r_415__3_,r_415__2_,r_415__1_,r_415__0_,r_416__63_,r_416__62_,
  r_416__61_,r_416__60_,r_416__59_,r_416__58_,r_416__57_,r_416__56_,r_416__55_,
  r_416__54_,r_416__53_,r_416__52_,r_416__51_,r_416__50_,r_416__49_,r_416__48_,
  r_416__47_,r_416__46_,r_416__45_,r_416__44_,r_416__43_,r_416__42_,r_416__41_,
  r_416__40_,r_416__39_,r_416__38_,r_416__37_,r_416__36_,r_416__35_,r_416__34_,r_416__33_,
  r_416__32_,r_416__31_,r_416__30_,r_416__29_,r_416__28_,r_416__27_,r_416__26_,
  r_416__25_,r_416__24_,r_416__23_,r_416__22_,r_416__21_,r_416__20_,r_416__19_,
  r_416__18_,r_416__17_,r_416__16_,r_416__15_,r_416__14_,r_416__13_,r_416__12_,
  r_416__11_,r_416__10_,r_416__9_,r_416__8_,r_416__7_,r_416__6_,r_416__5_,r_416__4_,
  r_416__3_,r_416__2_,r_416__1_,r_416__0_,r_417__63_,r_417__62_,r_417__61_,r_417__60_,
  r_417__59_,r_417__58_,r_417__57_,r_417__56_,r_417__55_,r_417__54_,r_417__53_,
  r_417__52_,r_417__51_,r_417__50_,r_417__49_,r_417__48_,r_417__47_,r_417__46_,
  r_417__45_,r_417__44_,r_417__43_,r_417__42_,r_417__41_,r_417__40_,r_417__39_,r_417__38_,
  r_417__37_,r_417__36_,r_417__35_,r_417__34_,r_417__33_,r_417__32_,r_417__31_,
  r_417__30_,r_417__29_,r_417__28_,r_417__27_,r_417__26_,r_417__25_,r_417__24_,
  r_417__23_,r_417__22_,r_417__21_,r_417__20_,r_417__19_,r_417__18_,r_417__17_,r_417__16_,
  r_417__15_,r_417__14_,r_417__13_,r_417__12_,r_417__11_,r_417__10_,r_417__9_,
  r_417__8_,r_417__7_,r_417__6_,r_417__5_,r_417__4_,r_417__3_,r_417__2_,r_417__1_,
  r_417__0_,r_418__63_,r_418__62_,r_418__61_,r_418__60_,r_418__59_,r_418__58_,
  r_418__57_,r_418__56_,r_418__55_,r_418__54_,r_418__53_,r_418__52_,r_418__51_,r_418__50_,
  r_418__49_,r_418__48_,r_418__47_,r_418__46_,r_418__45_,r_418__44_,r_418__43_,
  r_418__42_,r_418__41_,r_418__40_,r_418__39_,r_418__38_,r_418__37_,r_418__36_,
  r_418__35_,r_418__34_,r_418__33_,r_418__32_,r_418__31_,r_418__30_,r_418__29_,
  r_418__28_,r_418__27_,r_418__26_,r_418__25_,r_418__24_,r_418__23_,r_418__22_,r_418__21_,
  r_418__20_,r_418__19_,r_418__18_,r_418__17_,r_418__16_,r_418__15_,r_418__14_,
  r_418__13_,r_418__12_,r_418__11_,r_418__10_,r_418__9_,r_418__8_,r_418__7_,r_418__6_,
  r_418__5_,r_418__4_,r_418__3_,r_418__2_,r_418__1_,r_418__0_,r_419__63_,
  r_419__62_,r_419__61_,r_419__60_,r_419__59_,r_419__58_,r_419__57_,r_419__56_,r_419__55_,
  r_419__54_,r_419__53_,r_419__52_,r_419__51_,r_419__50_,r_419__49_,r_419__48_,
  r_419__47_,r_419__46_,r_419__45_,r_419__44_,r_419__43_,r_419__42_,r_419__41_,
  r_419__40_,r_419__39_,r_419__38_,r_419__37_,r_419__36_,r_419__35_,r_419__34_,
  r_419__33_,r_419__32_,r_419__31_,r_419__30_,r_419__29_,r_419__28_,r_419__27_,r_419__26_,
  r_419__25_,r_419__24_,r_419__23_,r_419__22_,r_419__21_,r_419__20_,r_419__19_,
  r_419__18_,r_419__17_,r_419__16_,r_419__15_,r_419__14_,r_419__13_,r_419__12_,
  r_419__11_,r_419__10_,r_419__9_,r_419__8_,r_419__7_,r_419__6_,r_419__5_,r_419__4_,
  r_419__3_,r_419__2_,r_419__1_,r_419__0_,r_420__63_,r_420__62_,r_420__61_,r_420__60_,
  r_420__59_,r_420__58_,r_420__57_,r_420__56_,r_420__55_,r_420__54_,r_420__53_,
  r_420__52_,r_420__51_,r_420__50_,r_420__49_,r_420__48_,r_420__47_,r_420__46_,
  r_420__45_,r_420__44_,r_420__43_,r_420__42_,r_420__41_,r_420__40_,r_420__39_,r_420__38_,
  r_420__37_,r_420__36_,r_420__35_,r_420__34_,r_420__33_,r_420__32_,r_420__31_,
  r_420__30_,r_420__29_,r_420__28_,r_420__27_,r_420__26_,r_420__25_,r_420__24_,
  r_420__23_,r_420__22_,r_420__21_,r_420__20_,r_420__19_,r_420__18_,r_420__17_,
  r_420__16_,r_420__15_,r_420__14_,r_420__13_,r_420__12_,r_420__11_,r_420__10_,r_420__9_,
  r_420__8_,r_420__7_,r_420__6_,r_420__5_,r_420__4_,r_420__3_,r_420__2_,r_420__1_,
  r_420__0_,r_421__63_,r_421__62_,r_421__61_,r_421__60_,r_421__59_,r_421__58_,
  r_421__57_,r_421__56_,r_421__55_,r_421__54_,r_421__53_,r_421__52_,r_421__51_,
  r_421__50_,r_421__49_,r_421__48_,r_421__47_,r_421__46_,r_421__45_,r_421__44_,r_421__43_,
  r_421__42_,r_421__41_,r_421__40_,r_421__39_,r_421__38_,r_421__37_,r_421__36_,
  r_421__35_,r_421__34_,r_421__33_,r_421__32_,r_421__31_,r_421__30_,r_421__29_,
  r_421__28_,r_421__27_,r_421__26_,r_421__25_,r_421__24_,r_421__23_,r_421__22_,
  r_421__21_,r_421__20_,r_421__19_,r_421__18_,r_421__17_,r_421__16_,r_421__15_,r_421__14_,
  r_421__13_,r_421__12_,r_421__11_,r_421__10_,r_421__9_,r_421__8_,r_421__7_,
  r_421__6_,r_421__5_,r_421__4_,r_421__3_,r_421__2_,r_421__1_,r_421__0_,r_422__63_,
  r_422__62_,r_422__61_,r_422__60_,r_422__59_,r_422__58_,r_422__57_,r_422__56_,
  r_422__55_,r_422__54_,r_422__53_,r_422__52_,r_422__51_,r_422__50_,r_422__49_,r_422__48_,
  r_422__47_,r_422__46_,r_422__45_,r_422__44_,r_422__43_,r_422__42_,r_422__41_,
  r_422__40_,r_422__39_,r_422__38_,r_422__37_,r_422__36_,r_422__35_,r_422__34_,
  r_422__33_,r_422__32_,r_422__31_,r_422__30_,r_422__29_,r_422__28_,r_422__27_,r_422__26_,
  r_422__25_,r_422__24_,r_422__23_,r_422__22_,r_422__21_,r_422__20_,r_422__19_,
  r_422__18_,r_422__17_,r_422__16_,r_422__15_,r_422__14_,r_422__13_,r_422__12_,
  r_422__11_,r_422__10_,r_422__9_,r_422__8_,r_422__7_,r_422__6_,r_422__5_,r_422__4_,
  r_422__3_,r_422__2_,r_422__1_,r_422__0_,r_423__63_,r_423__62_,r_423__61_,r_423__60_,
  r_423__59_,r_423__58_,r_423__57_,r_423__56_,r_423__55_,r_423__54_,r_423__53_,
  r_423__52_,r_423__51_,r_423__50_,r_423__49_,r_423__48_,r_423__47_,r_423__46_,
  r_423__45_,r_423__44_,r_423__43_,r_423__42_,r_423__41_,r_423__40_,r_423__39_,
  r_423__38_,r_423__37_,r_423__36_,r_423__35_,r_423__34_,r_423__33_,r_423__32_,r_423__31_,
  r_423__30_,r_423__29_,r_423__28_,r_423__27_,r_423__26_,r_423__25_,r_423__24_,
  r_423__23_,r_423__22_,r_423__21_,r_423__20_,r_423__19_,r_423__18_,r_423__17_,
  r_423__16_,r_423__15_,r_423__14_,r_423__13_,r_423__12_,r_423__11_,r_423__10_,r_423__9_,
  r_423__8_,r_423__7_,r_423__6_,r_423__5_,r_423__4_,r_423__3_,r_423__2_,r_423__1_,
  r_423__0_,r_424__63_,r_424__62_,r_424__61_,r_424__60_,r_424__59_,r_424__58_,
  r_424__57_,r_424__56_,r_424__55_,r_424__54_,r_424__53_,r_424__52_,r_424__51_,
  r_424__50_,r_424__49_,r_424__48_,r_424__47_,r_424__46_,r_424__45_,r_424__44_,
  r_424__43_,r_424__42_,r_424__41_,r_424__40_,r_424__39_,r_424__38_,r_424__37_,r_424__36_,
  r_424__35_,r_424__34_,r_424__33_,r_424__32_,r_424__31_,r_424__30_,r_424__29_,
  r_424__28_,r_424__27_,r_424__26_,r_424__25_,r_424__24_,r_424__23_,r_424__22_,
  r_424__21_,r_424__20_,r_424__19_,r_424__18_,r_424__17_,r_424__16_,r_424__15_,r_424__14_,
  r_424__13_,r_424__12_,r_424__11_,r_424__10_,r_424__9_,r_424__8_,r_424__7_,
  r_424__6_,r_424__5_,r_424__4_,r_424__3_,r_424__2_,r_424__1_,r_424__0_,r_425__63_,
  r_425__62_,r_425__61_,r_425__60_,r_425__59_,r_425__58_,r_425__57_,r_425__56_,
  r_425__55_,r_425__54_,r_425__53_,r_425__52_,r_425__51_,r_425__50_,r_425__49_,r_425__48_,
  r_425__47_,r_425__46_,r_425__45_,r_425__44_,r_425__43_,r_425__42_,r_425__41_,
  r_425__40_,r_425__39_,r_425__38_,r_425__37_,r_425__36_,r_425__35_,r_425__34_,
  r_425__33_,r_425__32_,r_425__31_,r_425__30_,r_425__29_,r_425__28_,r_425__27_,
  r_425__26_,r_425__25_,r_425__24_,r_425__23_,r_425__22_,r_425__21_,r_425__20_,r_425__19_,
  r_425__18_,r_425__17_,r_425__16_,r_425__15_,r_425__14_,r_425__13_,r_425__12_,
  r_425__11_,r_425__10_,r_425__9_,r_425__8_,r_425__7_,r_425__6_,r_425__5_,r_425__4_,
  r_425__3_,r_425__2_,r_425__1_,r_425__0_,r_426__63_,r_426__62_,r_426__61_,
  r_426__60_,r_426__59_,r_426__58_,r_426__57_,r_426__56_,r_426__55_,r_426__54_,r_426__53_,
  r_426__52_,r_426__51_,r_426__50_,r_426__49_,r_426__48_,r_426__47_,r_426__46_,
  r_426__45_,r_426__44_,r_426__43_,r_426__42_,r_426__41_,r_426__40_,r_426__39_,
  r_426__38_,r_426__37_,r_426__36_,r_426__35_,r_426__34_,r_426__33_,r_426__32_,
  r_426__31_,r_426__30_,r_426__29_,r_426__28_,r_426__27_,r_426__26_,r_426__25_,r_426__24_,
  r_426__23_,r_426__22_,r_426__21_,r_426__20_,r_426__19_,r_426__18_,r_426__17_,
  r_426__16_,r_426__15_,r_426__14_,r_426__13_,r_426__12_,r_426__11_,r_426__10_,
  r_426__9_,r_426__8_,r_426__7_,r_426__6_,r_426__5_,r_426__4_,r_426__3_,r_426__2_,
  r_426__1_,r_426__0_,r_427__63_,r_427__62_,r_427__61_,r_427__60_,r_427__59_,r_427__58_,
  r_427__57_,r_427__56_,r_427__55_,r_427__54_,r_427__53_,r_427__52_,r_427__51_,
  r_427__50_,r_427__49_,r_427__48_,r_427__47_,r_427__46_,r_427__45_,r_427__44_,
  r_427__43_,r_427__42_,r_427__41_,r_427__40_,r_427__39_,r_427__38_,r_427__37_,r_427__36_,
  r_427__35_,r_427__34_,r_427__33_,r_427__32_,r_427__31_,r_427__30_,r_427__29_,
  r_427__28_,r_427__27_,r_427__26_,r_427__25_,r_427__24_,r_427__23_,r_427__22_,
  r_427__21_,r_427__20_,r_427__19_,r_427__18_,r_427__17_,r_427__16_,r_427__15_,
  r_427__14_,r_427__13_,r_427__12_,r_427__11_,r_427__10_,r_427__9_,r_427__8_,r_427__7_,
  r_427__6_,r_427__5_,r_427__4_,r_427__3_,r_427__2_,r_427__1_,r_427__0_,r_428__63_,
  r_428__62_,r_428__61_,r_428__60_,r_428__59_,r_428__58_,r_428__57_,r_428__56_,
  r_428__55_,r_428__54_,r_428__53_,r_428__52_,r_428__51_,r_428__50_,r_428__49_,
  r_428__48_,r_428__47_,r_428__46_,r_428__45_,r_428__44_,r_428__43_,r_428__42_,r_428__41_,
  r_428__40_,r_428__39_,r_428__38_,r_428__37_,r_428__36_,r_428__35_,r_428__34_,
  r_428__33_,r_428__32_,r_428__31_,r_428__30_,r_428__29_,r_428__28_,r_428__27_,
  r_428__26_,r_428__25_,r_428__24_,r_428__23_,r_428__22_,r_428__21_,r_428__20_,
  r_428__19_,r_428__18_,r_428__17_,r_428__16_,r_428__15_,r_428__14_,r_428__13_,r_428__12_,
  r_428__11_,r_428__10_,r_428__9_,r_428__8_,r_428__7_,r_428__6_,r_428__5_,r_428__4_,
  r_428__3_,r_428__2_,r_428__1_,r_428__0_,r_429__63_,r_429__62_,r_429__61_,
  r_429__60_,r_429__59_,r_429__58_,r_429__57_,r_429__56_,r_429__55_,r_429__54_,
  r_429__53_,r_429__52_,r_429__51_,r_429__50_,r_429__49_,r_429__48_,r_429__47_,r_429__46_,
  r_429__45_,r_429__44_,r_429__43_,r_429__42_,r_429__41_,r_429__40_,r_429__39_,
  r_429__38_,r_429__37_,r_429__36_,r_429__35_,r_429__34_,r_429__33_,r_429__32_,
  r_429__31_,r_429__30_,r_429__29_,r_429__28_,r_429__27_,r_429__26_,r_429__25_,r_429__24_,
  r_429__23_,r_429__22_,r_429__21_,r_429__20_,r_429__19_,r_429__18_,r_429__17_,
  r_429__16_,r_429__15_,r_429__14_,r_429__13_,r_429__12_,r_429__11_,r_429__10_,
  r_429__9_,r_429__8_,r_429__7_,r_429__6_,r_429__5_,r_429__4_,r_429__3_,r_429__2_,
  r_429__1_,r_429__0_,r_430__63_,r_430__62_,r_430__61_,r_430__60_,r_430__59_,r_430__58_,
  r_430__57_,r_430__56_,r_430__55_,r_430__54_,r_430__53_,r_430__52_,r_430__51_,
  r_430__50_,r_430__49_,r_430__48_,r_430__47_,r_430__46_,r_430__45_,r_430__44_,
  r_430__43_,r_430__42_,r_430__41_,r_430__40_,r_430__39_,r_430__38_,r_430__37_,
  r_430__36_,r_430__35_,r_430__34_,r_430__33_,r_430__32_,r_430__31_,r_430__30_,r_430__29_,
  r_430__28_,r_430__27_,r_430__26_,r_430__25_,r_430__24_,r_430__23_,r_430__22_,
  r_430__21_,r_430__20_,r_430__19_,r_430__18_,r_430__17_,r_430__16_,r_430__15_,
  r_430__14_,r_430__13_,r_430__12_,r_430__11_,r_430__10_,r_430__9_,r_430__8_,r_430__7_,
  r_430__6_,r_430__5_,r_430__4_,r_430__3_,r_430__2_,r_430__1_,r_430__0_,r_431__63_,
  r_431__62_,r_431__61_,r_431__60_,r_431__59_,r_431__58_,r_431__57_,r_431__56_,
  r_431__55_,r_431__54_,r_431__53_,r_431__52_,r_431__51_,r_431__50_,r_431__49_,
  r_431__48_,r_431__47_,r_431__46_,r_431__45_,r_431__44_,r_431__43_,r_431__42_,
  r_431__41_,r_431__40_,r_431__39_,r_431__38_,r_431__37_,r_431__36_,r_431__35_,r_431__34_,
  r_431__33_,r_431__32_,r_431__31_,r_431__30_,r_431__29_,r_431__28_,r_431__27_,
  r_431__26_,r_431__25_,r_431__24_,r_431__23_,r_431__22_,r_431__21_,r_431__20_,
  r_431__19_,r_431__18_,r_431__17_,r_431__16_,r_431__15_,r_431__14_,r_431__13_,r_431__12_,
  r_431__11_,r_431__10_,r_431__9_,r_431__8_,r_431__7_,r_431__6_,r_431__5_,
  r_431__4_,r_431__3_,r_431__2_,r_431__1_,r_431__0_,r_432__63_,r_432__62_,r_432__61_,
  r_432__60_,r_432__59_,r_432__58_,r_432__57_,r_432__56_,r_432__55_,r_432__54_,
  r_432__53_,r_432__52_,r_432__51_,r_432__50_,r_432__49_,r_432__48_,r_432__47_,r_432__46_,
  r_432__45_,r_432__44_,r_432__43_,r_432__42_,r_432__41_,r_432__40_,r_432__39_,
  r_432__38_,r_432__37_,r_432__36_,r_432__35_,r_432__34_,r_432__33_,r_432__32_,
  r_432__31_,r_432__30_,r_432__29_,r_432__28_,r_432__27_,r_432__26_,r_432__25_,
  r_432__24_,r_432__23_,r_432__22_,r_432__21_,r_432__20_,r_432__19_,r_432__18_,r_432__17_,
  r_432__16_,r_432__15_,r_432__14_,r_432__13_,r_432__12_,r_432__11_,r_432__10_,
  r_432__9_,r_432__8_,r_432__7_,r_432__6_,r_432__5_,r_432__4_,r_432__3_,r_432__2_,
  r_432__1_,r_432__0_,r_433__63_,r_433__62_,r_433__61_,r_433__60_,r_433__59_,
  r_433__58_,r_433__57_,r_433__56_,r_433__55_,r_433__54_,r_433__53_,r_433__52_,r_433__51_,
  r_433__50_,r_433__49_,r_433__48_,r_433__47_,r_433__46_,r_433__45_,r_433__44_,
  r_433__43_,r_433__42_,r_433__41_,r_433__40_,r_433__39_,r_433__38_,r_433__37_,
  r_433__36_,r_433__35_,r_433__34_,r_433__33_,r_433__32_,r_433__31_,r_433__30_,
  r_433__29_,r_433__28_,r_433__27_,r_433__26_,r_433__25_,r_433__24_,r_433__23_,r_433__22_,
  r_433__21_,r_433__20_,r_433__19_,r_433__18_,r_433__17_,r_433__16_,r_433__15_,
  r_433__14_,r_433__13_,r_433__12_,r_433__11_,r_433__10_,r_433__9_,r_433__8_,r_433__7_,
  r_433__6_,r_433__5_,r_433__4_,r_433__3_,r_433__2_,r_433__1_,r_433__0_,
  r_434__63_,r_434__62_,r_434__61_,r_434__60_,r_434__59_,r_434__58_,r_434__57_,r_434__56_,
  r_434__55_,r_434__54_,r_434__53_,r_434__52_,r_434__51_,r_434__50_,r_434__49_,
  r_434__48_,r_434__47_,r_434__46_,r_434__45_,r_434__44_,r_434__43_,r_434__42_,
  r_434__41_,r_434__40_,r_434__39_,r_434__38_,r_434__37_,r_434__36_,r_434__35_,r_434__34_,
  r_434__33_,r_434__32_,r_434__31_,r_434__30_,r_434__29_,r_434__28_,r_434__27_,
  r_434__26_,r_434__25_,r_434__24_,r_434__23_,r_434__22_,r_434__21_,r_434__20_,
  r_434__19_,r_434__18_,r_434__17_,r_434__16_,r_434__15_,r_434__14_,r_434__13_,
  r_434__12_,r_434__11_,r_434__10_,r_434__9_,r_434__8_,r_434__7_,r_434__6_,r_434__5_,
  r_434__4_,r_434__3_,r_434__2_,r_434__1_,r_434__0_,r_435__63_,r_435__62_,r_435__61_,
  r_435__60_,r_435__59_,r_435__58_,r_435__57_,r_435__56_,r_435__55_,r_435__54_,
  r_435__53_,r_435__52_,r_435__51_,r_435__50_,r_435__49_,r_435__48_,r_435__47_,
  r_435__46_,r_435__45_,r_435__44_,r_435__43_,r_435__42_,r_435__41_,r_435__40_,r_435__39_,
  r_435__38_,r_435__37_,r_435__36_,r_435__35_,r_435__34_,r_435__33_,r_435__32_,
  r_435__31_,r_435__30_,r_435__29_,r_435__28_,r_435__27_,r_435__26_,r_435__25_,
  r_435__24_,r_435__23_,r_435__22_,r_435__21_,r_435__20_,r_435__19_,r_435__18_,
  r_435__17_,r_435__16_,r_435__15_,r_435__14_,r_435__13_,r_435__12_,r_435__11_,r_435__10_,
  r_435__9_,r_435__8_,r_435__7_,r_435__6_,r_435__5_,r_435__4_,r_435__3_,r_435__2_,
  r_435__1_,r_435__0_,r_436__63_,r_436__62_,r_436__61_,r_436__60_,r_436__59_,
  r_436__58_,r_436__57_,r_436__56_,r_436__55_,r_436__54_,r_436__53_,r_436__52_,
  r_436__51_,r_436__50_,r_436__49_,r_436__48_,r_436__47_,r_436__46_,r_436__45_,r_436__44_,
  r_436__43_,r_436__42_,r_436__41_,r_436__40_,r_436__39_,r_436__38_,r_436__37_,
  r_436__36_,r_436__35_,r_436__34_,r_436__33_,r_436__32_,r_436__31_,r_436__30_,
  r_436__29_,r_436__28_,r_436__27_,r_436__26_,r_436__25_,r_436__24_,r_436__23_,r_436__22_,
  r_436__21_,r_436__20_,r_436__19_,r_436__18_,r_436__17_,r_436__16_,r_436__15_,
  r_436__14_,r_436__13_,r_436__12_,r_436__11_,r_436__10_,r_436__9_,r_436__8_,
  r_436__7_,r_436__6_,r_436__5_,r_436__4_,r_436__3_,r_436__2_,r_436__1_,r_436__0_,
  r_437__63_,r_437__62_,r_437__61_,r_437__60_,r_437__59_,r_437__58_,r_437__57_,r_437__56_,
  r_437__55_,r_437__54_,r_437__53_,r_437__52_,r_437__51_,r_437__50_,r_437__49_,
  r_437__48_,r_437__47_,r_437__46_,r_437__45_,r_437__44_,r_437__43_,r_437__42_,
  r_437__41_,r_437__40_,r_437__39_,r_437__38_,r_437__37_,r_437__36_,r_437__35_,
  r_437__34_,r_437__33_,r_437__32_,r_437__31_,r_437__30_,r_437__29_,r_437__28_,r_437__27_,
  r_437__26_,r_437__25_,r_437__24_,r_437__23_,r_437__22_,r_437__21_,r_437__20_,
  r_437__19_,r_437__18_,r_437__17_,r_437__16_,r_437__15_,r_437__14_,r_437__13_,
  r_437__12_,r_437__11_,r_437__10_,r_437__9_,r_437__8_,r_437__7_,r_437__6_,r_437__5_,
  r_437__4_,r_437__3_,r_437__2_,r_437__1_,r_437__0_,r_438__63_,r_438__62_,r_438__61_,
  r_438__60_,r_438__59_,r_438__58_,r_438__57_,r_438__56_,r_438__55_,r_438__54_,
  r_438__53_,r_438__52_,r_438__51_,r_438__50_,r_438__49_,r_438__48_,r_438__47_,
  r_438__46_,r_438__45_,r_438__44_,r_438__43_,r_438__42_,r_438__41_,r_438__40_,
  r_438__39_,r_438__38_,r_438__37_,r_438__36_,r_438__35_,r_438__34_,r_438__33_,r_438__32_,
  r_438__31_,r_438__30_,r_438__29_,r_438__28_,r_438__27_,r_438__26_,r_438__25_,
  r_438__24_,r_438__23_,r_438__22_,r_438__21_,r_438__20_,r_438__19_,r_438__18_,
  r_438__17_,r_438__16_,r_438__15_,r_438__14_,r_438__13_,r_438__12_,r_438__11_,r_438__10_,
  r_438__9_,r_438__8_,r_438__7_,r_438__6_,r_438__5_,r_438__4_,r_438__3_,r_438__2_,
  r_438__1_,r_438__0_,r_439__63_,r_439__62_,r_439__61_,r_439__60_,r_439__59_,
  r_439__58_,r_439__57_,r_439__56_,r_439__55_,r_439__54_,r_439__53_,r_439__52_,
  r_439__51_,r_439__50_,r_439__49_,r_439__48_,r_439__47_,r_439__46_,r_439__45_,r_439__44_,
  r_439__43_,r_439__42_,r_439__41_,r_439__40_,r_439__39_,r_439__38_,r_439__37_,
  r_439__36_,r_439__35_,r_439__34_,r_439__33_,r_439__32_,r_439__31_,r_439__30_,
  r_439__29_,r_439__28_,r_439__27_,r_439__26_,r_439__25_,r_439__24_,r_439__23_,
  r_439__22_,r_439__21_,r_439__20_,r_439__19_,r_439__18_,r_439__17_,r_439__16_,r_439__15_,
  r_439__14_,r_439__13_,r_439__12_,r_439__11_,r_439__10_,r_439__9_,r_439__8_,
  r_439__7_,r_439__6_,r_439__5_,r_439__4_,r_439__3_,r_439__2_,r_439__1_,r_439__0_,
  r_440__63_,r_440__62_,r_440__61_,r_440__60_,r_440__59_,r_440__58_,r_440__57_,
  r_440__56_,r_440__55_,r_440__54_,r_440__53_,r_440__52_,r_440__51_,r_440__50_,r_440__49_,
  r_440__48_,r_440__47_,r_440__46_,r_440__45_,r_440__44_,r_440__43_,r_440__42_,
  r_440__41_,r_440__40_,r_440__39_,r_440__38_,r_440__37_,r_440__36_,r_440__35_,
  r_440__34_,r_440__33_,r_440__32_,r_440__31_,r_440__30_,r_440__29_,r_440__28_,
  r_440__27_,r_440__26_,r_440__25_,r_440__24_,r_440__23_,r_440__22_,r_440__21_,r_440__20_,
  r_440__19_,r_440__18_,r_440__17_,r_440__16_,r_440__15_,r_440__14_,r_440__13_,
  r_440__12_,r_440__11_,r_440__10_,r_440__9_,r_440__8_,r_440__7_,r_440__6_,r_440__5_,
  r_440__4_,r_440__3_,r_440__2_,r_440__1_,r_440__0_,r_441__63_,r_441__62_,
  r_441__61_,r_441__60_,r_441__59_,r_441__58_,r_441__57_,r_441__56_,r_441__55_,r_441__54_,
  r_441__53_,r_441__52_,r_441__51_,r_441__50_,r_441__49_,r_441__48_,r_441__47_,
  r_441__46_,r_441__45_,r_441__44_,r_441__43_,r_441__42_,r_441__41_,r_441__40_,
  r_441__39_,r_441__38_,r_441__37_,r_441__36_,r_441__35_,r_441__34_,r_441__33_,r_441__32_,
  r_441__31_,r_441__30_,r_441__29_,r_441__28_,r_441__27_,r_441__26_,r_441__25_,
  r_441__24_,r_441__23_,r_441__22_,r_441__21_,r_441__20_,r_441__19_,r_441__18_,
  r_441__17_,r_441__16_,r_441__15_,r_441__14_,r_441__13_,r_441__12_,r_441__11_,
  r_441__10_,r_441__9_,r_441__8_,r_441__7_,r_441__6_,r_441__5_,r_441__4_,r_441__3_,
  r_441__2_,r_441__1_,r_441__0_,r_442__63_,r_442__62_,r_442__61_,r_442__60_,r_442__59_,
  r_442__58_,r_442__57_,r_442__56_,r_442__55_,r_442__54_,r_442__53_,r_442__52_,
  r_442__51_,r_442__50_,r_442__49_,r_442__48_,r_442__47_,r_442__46_,r_442__45_,
  r_442__44_,r_442__43_,r_442__42_,r_442__41_,r_442__40_,r_442__39_,r_442__38_,r_442__37_,
  r_442__36_,r_442__35_,r_442__34_,r_442__33_,r_442__32_,r_442__31_,r_442__30_,
  r_442__29_,r_442__28_,r_442__27_,r_442__26_,r_442__25_,r_442__24_,r_442__23_,
  r_442__22_,r_442__21_,r_442__20_,r_442__19_,r_442__18_,r_442__17_,r_442__16_,
  r_442__15_,r_442__14_,r_442__13_,r_442__12_,r_442__11_,r_442__10_,r_442__9_,r_442__8_,
  r_442__7_,r_442__6_,r_442__5_,r_442__4_,r_442__3_,r_442__2_,r_442__1_,r_442__0_,
  r_443__63_,r_443__62_,r_443__61_,r_443__60_,r_443__59_,r_443__58_,r_443__57_,
  r_443__56_,r_443__55_,r_443__54_,r_443__53_,r_443__52_,r_443__51_,r_443__50_,
  r_443__49_,r_443__48_,r_443__47_,r_443__46_,r_443__45_,r_443__44_,r_443__43_,r_443__42_,
  r_443__41_,r_443__40_,r_443__39_,r_443__38_,r_443__37_,r_443__36_,r_443__35_,
  r_443__34_,r_443__33_,r_443__32_,r_443__31_,r_443__30_,r_443__29_,r_443__28_,
  r_443__27_,r_443__26_,r_443__25_,r_443__24_,r_443__23_,r_443__22_,r_443__21_,r_443__20_,
  r_443__19_,r_443__18_,r_443__17_,r_443__16_,r_443__15_,r_443__14_,r_443__13_,
  r_443__12_,r_443__11_,r_443__10_,r_443__9_,r_443__8_,r_443__7_,r_443__6_,r_443__5_,
  r_443__4_,r_443__3_,r_443__2_,r_443__1_,r_443__0_,r_444__63_,r_444__62_,
  r_444__61_,r_444__60_,r_444__59_,r_444__58_,r_444__57_,r_444__56_,r_444__55_,r_444__54_,
  r_444__53_,r_444__52_,r_444__51_,r_444__50_,r_444__49_,r_444__48_,r_444__47_,
  r_444__46_,r_444__45_,r_444__44_,r_444__43_,r_444__42_,r_444__41_,r_444__40_,
  r_444__39_,r_444__38_,r_444__37_,r_444__36_,r_444__35_,r_444__34_,r_444__33_,
  r_444__32_,r_444__31_,r_444__30_,r_444__29_,r_444__28_,r_444__27_,r_444__26_,r_444__25_,
  r_444__24_,r_444__23_,r_444__22_,r_444__21_,r_444__20_,r_444__19_,r_444__18_,
  r_444__17_,r_444__16_,r_444__15_,r_444__14_,r_444__13_,r_444__12_,r_444__11_,
  r_444__10_,r_444__9_,r_444__8_,r_444__7_,r_444__6_,r_444__5_,r_444__4_,r_444__3_,
  r_444__2_,r_444__1_,r_444__0_,r_445__63_,r_445__62_,r_445__61_,r_445__60_,r_445__59_,
  r_445__58_,r_445__57_,r_445__56_,r_445__55_,r_445__54_,r_445__53_,r_445__52_,
  r_445__51_,r_445__50_,r_445__49_,r_445__48_,r_445__47_,r_445__46_,r_445__45_,
  r_445__44_,r_445__43_,r_445__42_,r_445__41_,r_445__40_,r_445__39_,r_445__38_,
  r_445__37_,r_445__36_,r_445__35_,r_445__34_,r_445__33_,r_445__32_,r_445__31_,r_445__30_,
  r_445__29_,r_445__28_,r_445__27_,r_445__26_,r_445__25_,r_445__24_,r_445__23_,
  r_445__22_,r_445__21_,r_445__20_,r_445__19_,r_445__18_,r_445__17_,r_445__16_,
  r_445__15_,r_445__14_,r_445__13_,r_445__12_,r_445__11_,r_445__10_,r_445__9_,r_445__8_,
  r_445__7_,r_445__6_,r_445__5_,r_445__4_,r_445__3_,r_445__2_,r_445__1_,r_445__0_,
  r_446__63_,r_446__62_,r_446__61_,r_446__60_,r_446__59_,r_446__58_,r_446__57_,
  r_446__56_,r_446__55_,r_446__54_,r_446__53_,r_446__52_,r_446__51_,r_446__50_,
  r_446__49_,r_446__48_,r_446__47_,r_446__46_,r_446__45_,r_446__44_,r_446__43_,r_446__42_,
  r_446__41_,r_446__40_,r_446__39_,r_446__38_,r_446__37_,r_446__36_,r_446__35_,
  r_446__34_,r_446__33_,r_446__32_,r_446__31_,r_446__30_,r_446__29_,r_446__28_,
  r_446__27_,r_446__26_,r_446__25_,r_446__24_,r_446__23_,r_446__22_,r_446__21_,
  r_446__20_,r_446__19_,r_446__18_,r_446__17_,r_446__16_,r_446__15_,r_446__14_,r_446__13_,
  r_446__12_,r_446__11_,r_446__10_,r_446__9_,r_446__8_,r_446__7_,r_446__6_,
  r_446__5_,r_446__4_,r_446__3_,r_446__2_,r_446__1_,r_446__0_,r_447__63_,r_447__62_,
  r_447__61_,r_447__60_,r_447__59_,r_447__58_,r_447__57_,r_447__56_,r_447__55_,
  r_447__54_,r_447__53_,r_447__52_,r_447__51_,r_447__50_,r_447__49_,r_447__48_,r_447__47_,
  r_447__46_,r_447__45_,r_447__44_,r_447__43_,r_447__42_,r_447__41_,r_447__40_,
  r_447__39_,r_447__38_,r_447__37_,r_447__36_,r_447__35_,r_447__34_,r_447__33_,
  r_447__32_,r_447__31_,r_447__30_,r_447__29_,r_447__28_,r_447__27_,r_447__26_,
  r_447__25_,r_447__24_,r_447__23_,r_447__22_,r_447__21_,r_447__20_,r_447__19_,r_447__18_,
  r_447__17_,r_447__16_,r_447__15_,r_447__14_,r_447__13_,r_447__12_,r_447__11_,
  r_447__10_,r_447__9_,r_447__8_,r_447__7_,r_447__6_,r_447__5_,r_447__4_,r_447__3_,
  r_447__2_,r_447__1_,r_447__0_,r_448__63_,r_448__62_,r_448__61_,r_448__60_,
  r_448__59_,r_448__58_,r_448__57_,r_448__56_,r_448__55_,r_448__54_,r_448__53_,r_448__52_,
  r_448__51_,r_448__50_,r_448__49_,r_448__48_,r_448__47_,r_448__46_,r_448__45_,
  r_448__44_,r_448__43_,r_448__42_,r_448__41_,r_448__40_,r_448__39_,r_448__38_,
  r_448__37_,r_448__36_,r_448__35_,r_448__34_,r_448__33_,r_448__32_,r_448__31_,r_448__30_,
  r_448__29_,r_448__28_,r_448__27_,r_448__26_,r_448__25_,r_448__24_,r_448__23_,
  r_448__22_,r_448__21_,r_448__20_,r_448__19_,r_448__18_,r_448__17_,r_448__16_,
  r_448__15_,r_448__14_,r_448__13_,r_448__12_,r_448__11_,r_448__10_,r_448__9_,r_448__8_,
  r_448__7_,r_448__6_,r_448__5_,r_448__4_,r_448__3_,r_448__2_,r_448__1_,r_448__0_,
  r_449__63_,r_449__62_,r_449__61_,r_449__60_,r_449__59_,r_449__58_,r_449__57_,
  r_449__56_,r_449__55_,r_449__54_,r_449__53_,r_449__52_,r_449__51_,r_449__50_,
  r_449__49_,r_449__48_,r_449__47_,r_449__46_,r_449__45_,r_449__44_,r_449__43_,
  r_449__42_,r_449__41_,r_449__40_,r_449__39_,r_449__38_,r_449__37_,r_449__36_,r_449__35_,
  r_449__34_,r_449__33_,r_449__32_,r_449__31_,r_449__30_,r_449__29_,r_449__28_,
  r_449__27_,r_449__26_,r_449__25_,r_449__24_,r_449__23_,r_449__22_,r_449__21_,
  r_449__20_,r_449__19_,r_449__18_,r_449__17_,r_449__16_,r_449__15_,r_449__14_,
  r_449__13_,r_449__12_,r_449__11_,r_449__10_,r_449__9_,r_449__8_,r_449__7_,r_449__6_,
  r_449__5_,r_449__4_,r_449__3_,r_449__2_,r_449__1_,r_449__0_,r_450__63_,r_450__62_,
  r_450__61_,r_450__60_,r_450__59_,r_450__58_,r_450__57_,r_450__56_,r_450__55_,
  r_450__54_,r_450__53_,r_450__52_,r_450__51_,r_450__50_,r_450__49_,r_450__48_,
  r_450__47_,r_450__46_,r_450__45_,r_450__44_,r_450__43_,r_450__42_,r_450__41_,r_450__40_,
  r_450__39_,r_450__38_,r_450__37_,r_450__36_,r_450__35_,r_450__34_,r_450__33_,
  r_450__32_,r_450__31_,r_450__30_,r_450__29_,r_450__28_,r_450__27_,r_450__26_,
  r_450__25_,r_450__24_,r_450__23_,r_450__22_,r_450__21_,r_450__20_,r_450__19_,r_450__18_,
  r_450__17_,r_450__16_,r_450__15_,r_450__14_,r_450__13_,r_450__12_,r_450__11_,
  r_450__10_,r_450__9_,r_450__8_,r_450__7_,r_450__6_,r_450__5_,r_450__4_,r_450__3_,
  r_450__2_,r_450__1_,r_450__0_,r_451__63_,r_451__62_,r_451__61_,r_451__60_,
  r_451__59_,r_451__58_,r_451__57_,r_451__56_,r_451__55_,r_451__54_,r_451__53_,r_451__52_,
  r_451__51_,r_451__50_,r_451__49_,r_451__48_,r_451__47_,r_451__46_,r_451__45_,
  r_451__44_,r_451__43_,r_451__42_,r_451__41_,r_451__40_,r_451__39_,r_451__38_,
  r_451__37_,r_451__36_,r_451__35_,r_451__34_,r_451__33_,r_451__32_,r_451__31_,
  r_451__30_,r_451__29_,r_451__28_,r_451__27_,r_451__26_,r_451__25_,r_451__24_,r_451__23_,
  r_451__22_,r_451__21_,r_451__20_,r_451__19_,r_451__18_,r_451__17_,r_451__16_,
  r_451__15_,r_451__14_,r_451__13_,r_451__12_,r_451__11_,r_451__10_,r_451__9_,
  r_451__8_,r_451__7_,r_451__6_,r_451__5_,r_451__4_,r_451__3_,r_451__2_,r_451__1_,
  r_451__0_,r_452__63_,r_452__62_,r_452__61_,r_452__60_,r_452__59_,r_452__58_,r_452__57_,
  r_452__56_,r_452__55_,r_452__54_,r_452__53_,r_452__52_,r_452__51_,r_452__50_,
  r_452__49_,r_452__48_,r_452__47_,r_452__46_,r_452__45_,r_452__44_,r_452__43_,
  r_452__42_,r_452__41_,r_452__40_,r_452__39_,r_452__38_,r_452__37_,r_452__36_,
  r_452__35_,r_452__34_,r_452__33_,r_452__32_,r_452__31_,r_452__30_,r_452__29_,r_452__28_,
  r_452__27_,r_452__26_,r_452__25_,r_452__24_,r_452__23_,r_452__22_,r_452__21_,
  r_452__20_,r_452__19_,r_452__18_,r_452__17_,r_452__16_,r_452__15_,r_452__14_,
  r_452__13_,r_452__12_,r_452__11_,r_452__10_,r_452__9_,r_452__8_,r_452__7_,r_452__6_,
  r_452__5_,r_452__4_,r_452__3_,r_452__2_,r_452__1_,r_452__0_,r_453__63_,r_453__62_,
  r_453__61_,r_453__60_,r_453__59_,r_453__58_,r_453__57_,r_453__56_,r_453__55_,
  r_453__54_,r_453__53_,r_453__52_,r_453__51_,r_453__50_,r_453__49_,r_453__48_,
  r_453__47_,r_453__46_,r_453__45_,r_453__44_,r_453__43_,r_453__42_,r_453__41_,r_453__40_,
  r_453__39_,r_453__38_,r_453__37_,r_453__36_,r_453__35_,r_453__34_,r_453__33_,
  r_453__32_,r_453__31_,r_453__30_,r_453__29_,r_453__28_,r_453__27_,r_453__26_,
  r_453__25_,r_453__24_,r_453__23_,r_453__22_,r_453__21_,r_453__20_,r_453__19_,
  r_453__18_,r_453__17_,r_453__16_,r_453__15_,r_453__14_,r_453__13_,r_453__12_,r_453__11_,
  r_453__10_,r_453__9_,r_453__8_,r_453__7_,r_453__6_,r_453__5_,r_453__4_,r_453__3_,
  r_453__2_,r_453__1_,r_453__0_,r_454__63_,r_454__62_,r_454__61_,r_454__60_,
  r_454__59_,r_454__58_,r_454__57_,r_454__56_,r_454__55_,r_454__54_,r_454__53_,
  r_454__52_,r_454__51_,r_454__50_,r_454__49_,r_454__48_,r_454__47_,r_454__46_,r_454__45_,
  r_454__44_,r_454__43_,r_454__42_,r_454__41_,r_454__40_,r_454__39_,r_454__38_,
  r_454__37_,r_454__36_,r_454__35_,r_454__34_,r_454__33_,r_454__32_,r_454__31_,
  r_454__30_,r_454__29_,r_454__28_,r_454__27_,r_454__26_,r_454__25_,r_454__24_,
  r_454__23_,r_454__22_,r_454__21_,r_454__20_,r_454__19_,r_454__18_,r_454__17_,r_454__16_,
  r_454__15_,r_454__14_,r_454__13_,r_454__12_,r_454__11_,r_454__10_,r_454__9_,
  r_454__8_,r_454__7_,r_454__6_,r_454__5_,r_454__4_,r_454__3_,r_454__2_,r_454__1_,
  r_454__0_,r_455__63_,r_455__62_,r_455__61_,r_455__60_,r_455__59_,r_455__58_,
  r_455__57_,r_455__56_,r_455__55_,r_455__54_,r_455__53_,r_455__52_,r_455__51_,r_455__50_,
  r_455__49_,r_455__48_,r_455__47_,r_455__46_,r_455__45_,r_455__44_,r_455__43_,
  r_455__42_,r_455__41_,r_455__40_,r_455__39_,r_455__38_,r_455__37_,r_455__36_,
  r_455__35_,r_455__34_,r_455__33_,r_455__32_,r_455__31_,r_455__30_,r_455__29_,r_455__28_,
  r_455__27_,r_455__26_,r_455__25_,r_455__24_,r_455__23_,r_455__22_,r_455__21_,
  r_455__20_,r_455__19_,r_455__18_,r_455__17_,r_455__16_,r_455__15_,r_455__14_,
  r_455__13_,r_455__12_,r_455__11_,r_455__10_,r_455__9_,r_455__8_,r_455__7_,r_455__6_,
  r_455__5_,r_455__4_,r_455__3_,r_455__2_,r_455__1_,r_455__0_,r_456__63_,r_456__62_,
  r_456__61_,r_456__60_,r_456__59_,r_456__58_,r_456__57_,r_456__56_,r_456__55_,
  r_456__54_,r_456__53_,r_456__52_,r_456__51_,r_456__50_,r_456__49_,r_456__48_,
  r_456__47_,r_456__46_,r_456__45_,r_456__44_,r_456__43_,r_456__42_,r_456__41_,
  r_456__40_,r_456__39_,r_456__38_,r_456__37_,r_456__36_,r_456__35_,r_456__34_,r_456__33_,
  r_456__32_,r_456__31_,r_456__30_,r_456__29_,r_456__28_,r_456__27_,r_456__26_,
  r_456__25_,r_456__24_,r_456__23_,r_456__22_,r_456__21_,r_456__20_,r_456__19_,
  r_456__18_,r_456__17_,r_456__16_,r_456__15_,r_456__14_,r_456__13_,r_456__12_,
  r_456__11_,r_456__10_,r_456__9_,r_456__8_,r_456__7_,r_456__6_,r_456__5_,r_456__4_,
  r_456__3_,r_456__2_,r_456__1_,r_456__0_,r_457__63_,r_457__62_,r_457__61_,r_457__60_,
  r_457__59_,r_457__58_,r_457__57_,r_457__56_,r_457__55_,r_457__54_,r_457__53_,
  r_457__52_,r_457__51_,r_457__50_,r_457__49_,r_457__48_,r_457__47_,r_457__46_,
  r_457__45_,r_457__44_,r_457__43_,r_457__42_,r_457__41_,r_457__40_,r_457__39_,r_457__38_,
  r_457__37_,r_457__36_,r_457__35_,r_457__34_,r_457__33_,r_457__32_,r_457__31_,
  r_457__30_,r_457__29_,r_457__28_,r_457__27_,r_457__26_,r_457__25_,r_457__24_,
  r_457__23_,r_457__22_,r_457__21_,r_457__20_,r_457__19_,r_457__18_,r_457__17_,r_457__16_,
  r_457__15_,r_457__14_,r_457__13_,r_457__12_,r_457__11_,r_457__10_,r_457__9_,
  r_457__8_,r_457__7_,r_457__6_,r_457__5_,r_457__4_,r_457__3_,r_457__2_,r_457__1_,
  r_457__0_,r_458__63_,r_458__62_,r_458__61_,r_458__60_,r_458__59_,r_458__58_,
  r_458__57_,r_458__56_,r_458__55_,r_458__54_,r_458__53_,r_458__52_,r_458__51_,r_458__50_,
  r_458__49_,r_458__48_,r_458__47_,r_458__46_,r_458__45_,r_458__44_,r_458__43_,
  r_458__42_,r_458__41_,r_458__40_,r_458__39_,r_458__38_,r_458__37_,r_458__36_,
  r_458__35_,r_458__34_,r_458__33_,r_458__32_,r_458__31_,r_458__30_,r_458__29_,
  r_458__28_,r_458__27_,r_458__26_,r_458__25_,r_458__24_,r_458__23_,r_458__22_,r_458__21_,
  r_458__20_,r_458__19_,r_458__18_,r_458__17_,r_458__16_,r_458__15_,r_458__14_,
  r_458__13_,r_458__12_,r_458__11_,r_458__10_,r_458__9_,r_458__8_,r_458__7_,r_458__6_,
  r_458__5_,r_458__4_,r_458__3_,r_458__2_,r_458__1_,r_458__0_,r_459__63_,
  r_459__62_,r_459__61_,r_459__60_,r_459__59_,r_459__58_,r_459__57_,r_459__56_,r_459__55_,
  r_459__54_,r_459__53_,r_459__52_,r_459__51_,r_459__50_,r_459__49_,r_459__48_,
  r_459__47_,r_459__46_,r_459__45_,r_459__44_,r_459__43_,r_459__42_,r_459__41_,
  r_459__40_,r_459__39_,r_459__38_,r_459__37_,r_459__36_,r_459__35_,r_459__34_,
  r_459__33_,r_459__32_,r_459__31_,r_459__30_,r_459__29_,r_459__28_,r_459__27_,r_459__26_,
  r_459__25_,r_459__24_,r_459__23_,r_459__22_,r_459__21_,r_459__20_,r_459__19_,
  r_459__18_,r_459__17_,r_459__16_,r_459__15_,r_459__14_,r_459__13_,r_459__12_,
  r_459__11_,r_459__10_,r_459__9_,r_459__8_,r_459__7_,r_459__6_,r_459__5_,r_459__4_,
  r_459__3_,r_459__2_,r_459__1_,r_459__0_,r_460__63_,r_460__62_,r_460__61_,r_460__60_,
  r_460__59_,r_460__58_,r_460__57_,r_460__56_,r_460__55_,r_460__54_,r_460__53_,
  r_460__52_,r_460__51_,r_460__50_,r_460__49_,r_460__48_,r_460__47_,r_460__46_,
  r_460__45_,r_460__44_,r_460__43_,r_460__42_,r_460__41_,r_460__40_,r_460__39_,r_460__38_,
  r_460__37_,r_460__36_,r_460__35_,r_460__34_,r_460__33_,r_460__32_,r_460__31_,
  r_460__30_,r_460__29_,r_460__28_,r_460__27_,r_460__26_,r_460__25_,r_460__24_,
  r_460__23_,r_460__22_,r_460__21_,r_460__20_,r_460__19_,r_460__18_,r_460__17_,
  r_460__16_,r_460__15_,r_460__14_,r_460__13_,r_460__12_,r_460__11_,r_460__10_,r_460__9_,
  r_460__8_,r_460__7_,r_460__6_,r_460__5_,r_460__4_,r_460__3_,r_460__2_,r_460__1_,
  r_460__0_,r_461__63_,r_461__62_,r_461__61_,r_461__60_,r_461__59_,r_461__58_,
  r_461__57_,r_461__56_,r_461__55_,r_461__54_,r_461__53_,r_461__52_,r_461__51_,
  r_461__50_,r_461__49_,r_461__48_,r_461__47_,r_461__46_,r_461__45_,r_461__44_,r_461__43_,
  r_461__42_,r_461__41_,r_461__40_,r_461__39_,r_461__38_,r_461__37_,r_461__36_,
  r_461__35_,r_461__34_,r_461__33_,r_461__32_,r_461__31_,r_461__30_,r_461__29_,
  r_461__28_,r_461__27_,r_461__26_,r_461__25_,r_461__24_,r_461__23_,r_461__22_,
  r_461__21_,r_461__20_,r_461__19_,r_461__18_,r_461__17_,r_461__16_,r_461__15_,r_461__14_,
  r_461__13_,r_461__12_,r_461__11_,r_461__10_,r_461__9_,r_461__8_,r_461__7_,
  r_461__6_,r_461__5_,r_461__4_,r_461__3_,r_461__2_,r_461__1_,r_461__0_,r_462__63_,
  r_462__62_,r_462__61_,r_462__60_,r_462__59_,r_462__58_,r_462__57_,r_462__56_,
  r_462__55_,r_462__54_,r_462__53_,r_462__52_,r_462__51_,r_462__50_,r_462__49_,r_462__48_,
  r_462__47_,r_462__46_,r_462__45_,r_462__44_,r_462__43_,r_462__42_,r_462__41_,
  r_462__40_,r_462__39_,r_462__38_,r_462__37_,r_462__36_,r_462__35_,r_462__34_,
  r_462__33_,r_462__32_,r_462__31_,r_462__30_,r_462__29_,r_462__28_,r_462__27_,r_462__26_,
  r_462__25_,r_462__24_,r_462__23_,r_462__22_,r_462__21_,r_462__20_,r_462__19_,
  r_462__18_,r_462__17_,r_462__16_,r_462__15_,r_462__14_,r_462__13_,r_462__12_,
  r_462__11_,r_462__10_,r_462__9_,r_462__8_,r_462__7_,r_462__6_,r_462__5_,r_462__4_,
  r_462__3_,r_462__2_,r_462__1_,r_462__0_,r_463__63_,r_463__62_,r_463__61_,r_463__60_,
  r_463__59_,r_463__58_,r_463__57_,r_463__56_,r_463__55_,r_463__54_,r_463__53_,
  r_463__52_,r_463__51_,r_463__50_,r_463__49_,r_463__48_,r_463__47_,r_463__46_,
  r_463__45_,r_463__44_,r_463__43_,r_463__42_,r_463__41_,r_463__40_,r_463__39_,
  r_463__38_,r_463__37_,r_463__36_,r_463__35_,r_463__34_,r_463__33_,r_463__32_,r_463__31_,
  r_463__30_,r_463__29_,r_463__28_,r_463__27_,r_463__26_,r_463__25_,r_463__24_,
  r_463__23_,r_463__22_,r_463__21_,r_463__20_,r_463__19_,r_463__18_,r_463__17_,
  r_463__16_,r_463__15_,r_463__14_,r_463__13_,r_463__12_,r_463__11_,r_463__10_,r_463__9_,
  r_463__8_,r_463__7_,r_463__6_,r_463__5_,r_463__4_,r_463__3_,r_463__2_,r_463__1_,
  r_463__0_,r_464__63_,r_464__62_,r_464__61_,r_464__60_,r_464__59_,r_464__58_,
  r_464__57_,r_464__56_,r_464__55_,r_464__54_,r_464__53_,r_464__52_,r_464__51_,
  r_464__50_,r_464__49_,r_464__48_,r_464__47_,r_464__46_,r_464__45_,r_464__44_,
  r_464__43_,r_464__42_,r_464__41_,r_464__40_,r_464__39_,r_464__38_,r_464__37_,r_464__36_,
  r_464__35_,r_464__34_,r_464__33_,r_464__32_,r_464__31_,r_464__30_,r_464__29_,
  r_464__28_,r_464__27_,r_464__26_,r_464__25_,r_464__24_,r_464__23_,r_464__22_,
  r_464__21_,r_464__20_,r_464__19_,r_464__18_,r_464__17_,r_464__16_,r_464__15_,r_464__14_,
  r_464__13_,r_464__12_,r_464__11_,r_464__10_,r_464__9_,r_464__8_,r_464__7_,
  r_464__6_,r_464__5_,r_464__4_,r_464__3_,r_464__2_,r_464__1_,r_464__0_,r_465__63_,
  r_465__62_,r_465__61_,r_465__60_,r_465__59_,r_465__58_,r_465__57_,r_465__56_,
  r_465__55_,r_465__54_,r_465__53_,r_465__52_,r_465__51_,r_465__50_,r_465__49_,r_465__48_,
  r_465__47_,r_465__46_,r_465__45_,r_465__44_,r_465__43_,r_465__42_,r_465__41_,
  r_465__40_,r_465__39_,r_465__38_,r_465__37_,r_465__36_,r_465__35_,r_465__34_,
  r_465__33_,r_465__32_,r_465__31_,r_465__30_,r_465__29_,r_465__28_,r_465__27_,
  r_465__26_,r_465__25_,r_465__24_,r_465__23_,r_465__22_,r_465__21_,r_465__20_,r_465__19_,
  r_465__18_,r_465__17_,r_465__16_,r_465__15_,r_465__14_,r_465__13_,r_465__12_,
  r_465__11_,r_465__10_,r_465__9_,r_465__8_,r_465__7_,r_465__6_,r_465__5_,r_465__4_,
  r_465__3_,r_465__2_,r_465__1_,r_465__0_,r_466__63_,r_466__62_,r_466__61_,
  r_466__60_,r_466__59_,r_466__58_,r_466__57_,r_466__56_,r_466__55_,r_466__54_,r_466__53_,
  r_466__52_,r_466__51_,r_466__50_,r_466__49_,r_466__48_,r_466__47_,r_466__46_,
  r_466__45_,r_466__44_,r_466__43_,r_466__42_,r_466__41_,r_466__40_,r_466__39_,
  r_466__38_,r_466__37_,r_466__36_,r_466__35_,r_466__34_,r_466__33_,r_466__32_,
  r_466__31_,r_466__30_,r_466__29_,r_466__28_,r_466__27_,r_466__26_,r_466__25_,r_466__24_,
  r_466__23_,r_466__22_,r_466__21_,r_466__20_,r_466__19_,r_466__18_,r_466__17_,
  r_466__16_,r_466__15_,r_466__14_,r_466__13_,r_466__12_,r_466__11_,r_466__10_,
  r_466__9_,r_466__8_,r_466__7_,r_466__6_,r_466__5_,r_466__4_,r_466__3_,r_466__2_,
  r_466__1_,r_466__0_,r_467__63_,r_467__62_,r_467__61_,r_467__60_,r_467__59_,r_467__58_,
  r_467__57_,r_467__56_,r_467__55_,r_467__54_,r_467__53_,r_467__52_,r_467__51_,
  r_467__50_,r_467__49_,r_467__48_,r_467__47_,r_467__46_,r_467__45_,r_467__44_,
  r_467__43_,r_467__42_,r_467__41_,r_467__40_,r_467__39_,r_467__38_,r_467__37_,r_467__36_,
  r_467__35_,r_467__34_,r_467__33_,r_467__32_,r_467__31_,r_467__30_,r_467__29_,
  r_467__28_,r_467__27_,r_467__26_,r_467__25_,r_467__24_,r_467__23_,r_467__22_,
  r_467__21_,r_467__20_,r_467__19_,r_467__18_,r_467__17_,r_467__16_,r_467__15_,
  r_467__14_,r_467__13_,r_467__12_,r_467__11_,r_467__10_,r_467__9_,r_467__8_,r_467__7_,
  r_467__6_,r_467__5_,r_467__4_,r_467__3_,r_467__2_,r_467__1_,r_467__0_,r_468__63_,
  r_468__62_,r_468__61_,r_468__60_,r_468__59_,r_468__58_,r_468__57_,r_468__56_,
  r_468__55_,r_468__54_,r_468__53_,r_468__52_,r_468__51_,r_468__50_,r_468__49_,
  r_468__48_,r_468__47_,r_468__46_,r_468__45_,r_468__44_,r_468__43_,r_468__42_,r_468__41_,
  r_468__40_,r_468__39_,r_468__38_,r_468__37_,r_468__36_,r_468__35_,r_468__34_,
  r_468__33_,r_468__32_,r_468__31_,r_468__30_,r_468__29_,r_468__28_,r_468__27_,
  r_468__26_,r_468__25_,r_468__24_,r_468__23_,r_468__22_,r_468__21_,r_468__20_,
  r_468__19_,r_468__18_,r_468__17_,r_468__16_,r_468__15_,r_468__14_,r_468__13_,r_468__12_,
  r_468__11_,r_468__10_,r_468__9_,r_468__8_,r_468__7_,r_468__6_,r_468__5_,r_468__4_,
  r_468__3_,r_468__2_,r_468__1_,r_468__0_,r_469__63_,r_469__62_,r_469__61_,
  r_469__60_,r_469__59_,r_469__58_,r_469__57_,r_469__56_,r_469__55_,r_469__54_,
  r_469__53_,r_469__52_,r_469__51_,r_469__50_,r_469__49_,r_469__48_,r_469__47_,r_469__46_,
  r_469__45_,r_469__44_,r_469__43_,r_469__42_,r_469__41_,r_469__40_,r_469__39_,
  r_469__38_,r_469__37_,r_469__36_,r_469__35_,r_469__34_,r_469__33_,r_469__32_,
  r_469__31_,r_469__30_,r_469__29_,r_469__28_,r_469__27_,r_469__26_,r_469__25_,r_469__24_,
  r_469__23_,r_469__22_,r_469__21_,r_469__20_,r_469__19_,r_469__18_,r_469__17_,
  r_469__16_,r_469__15_,r_469__14_,r_469__13_,r_469__12_,r_469__11_,r_469__10_,
  r_469__9_,r_469__8_,r_469__7_,r_469__6_,r_469__5_,r_469__4_,r_469__3_,r_469__2_,
  r_469__1_,r_469__0_,r_470__63_,r_470__62_,r_470__61_,r_470__60_,r_470__59_,r_470__58_,
  r_470__57_,r_470__56_,r_470__55_,r_470__54_,r_470__53_,r_470__52_,r_470__51_,
  r_470__50_,r_470__49_,r_470__48_,r_470__47_,r_470__46_,r_470__45_,r_470__44_,
  r_470__43_,r_470__42_,r_470__41_,r_470__40_,r_470__39_,r_470__38_,r_470__37_,
  r_470__36_,r_470__35_,r_470__34_,r_470__33_,r_470__32_,r_470__31_,r_470__30_,r_470__29_,
  r_470__28_,r_470__27_,r_470__26_,r_470__25_,r_470__24_,r_470__23_,r_470__22_,
  r_470__21_,r_470__20_,r_470__19_,r_470__18_,r_470__17_,r_470__16_,r_470__15_,
  r_470__14_,r_470__13_,r_470__12_,r_470__11_,r_470__10_,r_470__9_,r_470__8_,r_470__7_,
  r_470__6_,r_470__5_,r_470__4_,r_470__3_,r_470__2_,r_470__1_,r_470__0_,r_471__63_,
  r_471__62_,r_471__61_,r_471__60_,r_471__59_,r_471__58_,r_471__57_,r_471__56_,
  r_471__55_,r_471__54_,r_471__53_,r_471__52_,r_471__51_,r_471__50_,r_471__49_,
  r_471__48_,r_471__47_,r_471__46_,r_471__45_,r_471__44_,r_471__43_,r_471__42_,
  r_471__41_,r_471__40_,r_471__39_,r_471__38_,r_471__37_,r_471__36_,r_471__35_,r_471__34_,
  r_471__33_,r_471__32_,r_471__31_,r_471__30_,r_471__29_,r_471__28_,r_471__27_,
  r_471__26_,r_471__25_,r_471__24_,r_471__23_,r_471__22_,r_471__21_,r_471__20_,
  r_471__19_,r_471__18_,r_471__17_,r_471__16_,r_471__15_,r_471__14_,r_471__13_,r_471__12_,
  r_471__11_,r_471__10_,r_471__9_,r_471__8_,r_471__7_,r_471__6_,r_471__5_,
  r_471__4_,r_471__3_,r_471__2_,r_471__1_,r_471__0_,r_472__63_,r_472__62_,r_472__61_,
  r_472__60_,r_472__59_,r_472__58_,r_472__57_,r_472__56_,r_472__55_,r_472__54_,
  r_472__53_,r_472__52_,r_472__51_,r_472__50_,r_472__49_,r_472__48_,r_472__47_,r_472__46_,
  r_472__45_,r_472__44_,r_472__43_,r_472__42_,r_472__41_,r_472__40_,r_472__39_,
  r_472__38_,r_472__37_,r_472__36_,r_472__35_,r_472__34_,r_472__33_,r_472__32_,
  r_472__31_,r_472__30_,r_472__29_,r_472__28_,r_472__27_,r_472__26_,r_472__25_,
  r_472__24_,r_472__23_,r_472__22_,r_472__21_,r_472__20_,r_472__19_,r_472__18_,r_472__17_,
  r_472__16_,r_472__15_,r_472__14_,r_472__13_,r_472__12_,r_472__11_,r_472__10_,
  r_472__9_,r_472__8_,r_472__7_,r_472__6_,r_472__5_,r_472__4_,r_472__3_,r_472__2_,
  r_472__1_,r_472__0_,r_473__63_,r_473__62_,r_473__61_,r_473__60_,r_473__59_,
  r_473__58_,r_473__57_,r_473__56_,r_473__55_,r_473__54_,r_473__53_,r_473__52_,r_473__51_,
  r_473__50_,r_473__49_,r_473__48_,r_473__47_,r_473__46_,r_473__45_,r_473__44_,
  r_473__43_,r_473__42_,r_473__41_,r_473__40_,r_473__39_,r_473__38_,r_473__37_,
  r_473__36_,r_473__35_,r_473__34_,r_473__33_,r_473__32_,r_473__31_,r_473__30_,
  r_473__29_,r_473__28_,r_473__27_,r_473__26_,r_473__25_,r_473__24_,r_473__23_,r_473__22_,
  r_473__21_,r_473__20_,r_473__19_,r_473__18_,r_473__17_,r_473__16_,r_473__15_,
  r_473__14_,r_473__13_,r_473__12_,r_473__11_,r_473__10_,r_473__9_,r_473__8_,r_473__7_,
  r_473__6_,r_473__5_,r_473__4_,r_473__3_,r_473__2_,r_473__1_,r_473__0_,
  r_474__63_,r_474__62_,r_474__61_,r_474__60_,r_474__59_,r_474__58_,r_474__57_,r_474__56_,
  r_474__55_,r_474__54_,r_474__53_,r_474__52_,r_474__51_,r_474__50_,r_474__49_,
  r_474__48_,r_474__47_,r_474__46_,r_474__45_,r_474__44_,r_474__43_,r_474__42_,
  r_474__41_,r_474__40_,r_474__39_,r_474__38_,r_474__37_,r_474__36_,r_474__35_,r_474__34_,
  r_474__33_,r_474__32_,r_474__31_,r_474__30_,r_474__29_,r_474__28_,r_474__27_,
  r_474__26_,r_474__25_,r_474__24_,r_474__23_,r_474__22_,r_474__21_,r_474__20_,
  r_474__19_,r_474__18_,r_474__17_,r_474__16_,r_474__15_,r_474__14_,r_474__13_,
  r_474__12_,r_474__11_,r_474__10_,r_474__9_,r_474__8_,r_474__7_,r_474__6_,r_474__5_,
  r_474__4_,r_474__3_,r_474__2_,r_474__1_,r_474__0_,r_475__63_,r_475__62_,r_475__61_,
  r_475__60_,r_475__59_,r_475__58_,r_475__57_,r_475__56_,r_475__55_,r_475__54_,
  r_475__53_,r_475__52_,r_475__51_,r_475__50_,r_475__49_,r_475__48_,r_475__47_,
  r_475__46_,r_475__45_,r_475__44_,r_475__43_,r_475__42_,r_475__41_,r_475__40_,r_475__39_,
  r_475__38_,r_475__37_,r_475__36_,r_475__35_,r_475__34_,r_475__33_,r_475__32_,
  r_475__31_,r_475__30_,r_475__29_,r_475__28_,r_475__27_,r_475__26_,r_475__25_,
  r_475__24_,r_475__23_,r_475__22_,r_475__21_,r_475__20_,r_475__19_,r_475__18_,
  r_475__17_,r_475__16_,r_475__15_,r_475__14_,r_475__13_,r_475__12_,r_475__11_,r_475__10_,
  r_475__9_,r_475__8_,r_475__7_,r_475__6_,r_475__5_,r_475__4_,r_475__3_,r_475__2_,
  r_475__1_,r_475__0_,r_476__63_,r_476__62_,r_476__61_,r_476__60_,r_476__59_,
  r_476__58_,r_476__57_,r_476__56_,r_476__55_,r_476__54_,r_476__53_,r_476__52_,
  r_476__51_,r_476__50_,r_476__49_,r_476__48_,r_476__47_,r_476__46_,r_476__45_,r_476__44_,
  r_476__43_,r_476__42_,r_476__41_,r_476__40_,r_476__39_,r_476__38_,r_476__37_,
  r_476__36_,r_476__35_,r_476__34_,r_476__33_,r_476__32_,r_476__31_,r_476__30_,
  r_476__29_,r_476__28_,r_476__27_,r_476__26_,r_476__25_,r_476__24_,r_476__23_,r_476__22_,
  r_476__21_,r_476__20_,r_476__19_,r_476__18_,r_476__17_,r_476__16_,r_476__15_,
  r_476__14_,r_476__13_,r_476__12_,r_476__11_,r_476__10_,r_476__9_,r_476__8_,
  r_476__7_,r_476__6_,r_476__5_,r_476__4_,r_476__3_,r_476__2_,r_476__1_,r_476__0_,
  r_477__63_,r_477__62_,r_477__61_,r_477__60_,r_477__59_,r_477__58_,r_477__57_,r_477__56_,
  r_477__55_,r_477__54_,r_477__53_,r_477__52_,r_477__51_,r_477__50_,r_477__49_,
  r_477__48_,r_477__47_,r_477__46_,r_477__45_,r_477__44_,r_477__43_,r_477__42_,
  r_477__41_,r_477__40_,r_477__39_,r_477__38_,r_477__37_,r_477__36_,r_477__35_,
  r_477__34_,r_477__33_,r_477__32_,r_477__31_,r_477__30_,r_477__29_,r_477__28_,r_477__27_,
  r_477__26_,r_477__25_,r_477__24_,r_477__23_,r_477__22_,r_477__21_,r_477__20_,
  r_477__19_,r_477__18_,r_477__17_,r_477__16_,r_477__15_,r_477__14_,r_477__13_,
  r_477__12_,r_477__11_,r_477__10_,r_477__9_,r_477__8_,r_477__7_,r_477__6_,r_477__5_,
  r_477__4_,r_477__3_,r_477__2_,r_477__1_,r_477__0_,r_478__63_,r_478__62_,r_478__61_,
  r_478__60_,r_478__59_,r_478__58_,r_478__57_,r_478__56_,r_478__55_,r_478__54_,
  r_478__53_,r_478__52_,r_478__51_,r_478__50_,r_478__49_,r_478__48_,r_478__47_,
  r_478__46_,r_478__45_,r_478__44_,r_478__43_,r_478__42_,r_478__41_,r_478__40_,
  r_478__39_,r_478__38_,r_478__37_,r_478__36_,r_478__35_,r_478__34_,r_478__33_,r_478__32_,
  r_478__31_,r_478__30_,r_478__29_,r_478__28_,r_478__27_,r_478__26_,r_478__25_,
  r_478__24_,r_478__23_,r_478__22_,r_478__21_,r_478__20_,r_478__19_,r_478__18_,
  r_478__17_,r_478__16_,r_478__15_,r_478__14_,r_478__13_,r_478__12_,r_478__11_,r_478__10_,
  r_478__9_,r_478__8_,r_478__7_,r_478__6_,r_478__5_,r_478__4_,r_478__3_,r_478__2_,
  r_478__1_,r_478__0_,r_479__63_,r_479__62_,r_479__61_,r_479__60_,r_479__59_,
  r_479__58_,r_479__57_,r_479__56_,r_479__55_,r_479__54_,r_479__53_,r_479__52_,
  r_479__51_,r_479__50_,r_479__49_,r_479__48_,r_479__47_,r_479__46_,r_479__45_,r_479__44_,
  r_479__43_,r_479__42_,r_479__41_,r_479__40_,r_479__39_,r_479__38_,r_479__37_,
  r_479__36_,r_479__35_,r_479__34_,r_479__33_,r_479__32_,r_479__31_,r_479__30_,
  r_479__29_,r_479__28_,r_479__27_,r_479__26_,r_479__25_,r_479__24_,r_479__23_,
  r_479__22_,r_479__21_,r_479__20_,r_479__19_,r_479__18_,r_479__17_,r_479__16_,r_479__15_,
  r_479__14_,r_479__13_,r_479__12_,r_479__11_,r_479__10_,r_479__9_,r_479__8_,
  r_479__7_,r_479__6_,r_479__5_,r_479__4_,r_479__3_,r_479__2_,r_479__1_,r_479__0_,
  r_480__63_,r_480__62_,r_480__61_,r_480__60_,r_480__59_,r_480__58_,r_480__57_,
  r_480__56_,r_480__55_,r_480__54_,r_480__53_,r_480__52_,r_480__51_,r_480__50_,r_480__49_,
  r_480__48_,r_480__47_,r_480__46_,r_480__45_,r_480__44_,r_480__43_,r_480__42_,
  r_480__41_,r_480__40_,r_480__39_,r_480__38_,r_480__37_,r_480__36_,r_480__35_,
  r_480__34_,r_480__33_,r_480__32_,r_480__31_,r_480__30_,r_480__29_,r_480__28_,
  r_480__27_,r_480__26_,r_480__25_,r_480__24_,r_480__23_,r_480__22_,r_480__21_,r_480__20_,
  r_480__19_,r_480__18_,r_480__17_,r_480__16_,r_480__15_,r_480__14_,r_480__13_,
  r_480__12_,r_480__11_,r_480__10_,r_480__9_,r_480__8_,r_480__7_,r_480__6_,r_480__5_,
  r_480__4_,r_480__3_,r_480__2_,r_480__1_,r_480__0_,r_481__63_,r_481__62_,
  r_481__61_,r_481__60_,r_481__59_,r_481__58_,r_481__57_,r_481__56_,r_481__55_,r_481__54_,
  r_481__53_,r_481__52_,r_481__51_,r_481__50_,r_481__49_,r_481__48_,r_481__47_,
  r_481__46_,r_481__45_,r_481__44_,r_481__43_,r_481__42_,r_481__41_,r_481__40_,
  r_481__39_,r_481__38_,r_481__37_,r_481__36_,r_481__35_,r_481__34_,r_481__33_,r_481__32_,
  r_481__31_,r_481__30_,r_481__29_,r_481__28_,r_481__27_,r_481__26_,r_481__25_,
  r_481__24_,r_481__23_,r_481__22_,r_481__21_,r_481__20_,r_481__19_,r_481__18_,
  r_481__17_,r_481__16_,r_481__15_,r_481__14_,r_481__13_,r_481__12_,r_481__11_,
  r_481__10_,r_481__9_,r_481__8_,r_481__7_,r_481__6_,r_481__5_,r_481__4_,r_481__3_,
  r_481__2_,r_481__1_,r_481__0_,r_482__63_,r_482__62_,r_482__61_,r_482__60_,r_482__59_,
  r_482__58_,r_482__57_,r_482__56_,r_482__55_,r_482__54_,r_482__53_,r_482__52_,
  r_482__51_,r_482__50_,r_482__49_,r_482__48_,r_482__47_,r_482__46_,r_482__45_,
  r_482__44_,r_482__43_,r_482__42_,r_482__41_,r_482__40_,r_482__39_,r_482__38_,r_482__37_,
  r_482__36_,r_482__35_,r_482__34_,r_482__33_,r_482__32_,r_482__31_,r_482__30_,
  r_482__29_,r_482__28_,r_482__27_,r_482__26_,r_482__25_,r_482__24_,r_482__23_,
  r_482__22_,r_482__21_,r_482__20_,r_482__19_,r_482__18_,r_482__17_,r_482__16_,
  r_482__15_,r_482__14_,r_482__13_,r_482__12_,r_482__11_,r_482__10_,r_482__9_,r_482__8_,
  r_482__7_,r_482__6_,r_482__5_,r_482__4_,r_482__3_,r_482__2_,r_482__1_,r_482__0_,
  r_483__63_,r_483__62_,r_483__61_,r_483__60_,r_483__59_,r_483__58_,r_483__57_,
  r_483__56_,r_483__55_,r_483__54_,r_483__53_,r_483__52_,r_483__51_,r_483__50_,
  r_483__49_,r_483__48_,r_483__47_,r_483__46_,r_483__45_,r_483__44_,r_483__43_,r_483__42_,
  r_483__41_,r_483__40_,r_483__39_,r_483__38_,r_483__37_,r_483__36_,r_483__35_,
  r_483__34_,r_483__33_,r_483__32_,r_483__31_,r_483__30_,r_483__29_,r_483__28_,
  r_483__27_,r_483__26_,r_483__25_,r_483__24_,r_483__23_,r_483__22_,r_483__21_,r_483__20_,
  r_483__19_,r_483__18_,r_483__17_,r_483__16_,r_483__15_,r_483__14_,r_483__13_,
  r_483__12_,r_483__11_,r_483__10_,r_483__9_,r_483__8_,r_483__7_,r_483__6_,r_483__5_,
  r_483__4_,r_483__3_,r_483__2_,r_483__1_,r_483__0_,r_484__63_,r_484__62_,
  r_484__61_,r_484__60_,r_484__59_,r_484__58_,r_484__57_,r_484__56_,r_484__55_,r_484__54_,
  r_484__53_,r_484__52_,r_484__51_,r_484__50_,r_484__49_,r_484__48_,r_484__47_,
  r_484__46_,r_484__45_,r_484__44_,r_484__43_,r_484__42_,r_484__41_,r_484__40_,
  r_484__39_,r_484__38_,r_484__37_,r_484__36_,r_484__35_,r_484__34_,r_484__33_,
  r_484__32_,r_484__31_,r_484__30_,r_484__29_,r_484__28_,r_484__27_,r_484__26_,r_484__25_,
  r_484__24_,r_484__23_,r_484__22_,r_484__21_,r_484__20_,r_484__19_,r_484__18_,
  r_484__17_,r_484__16_,r_484__15_,r_484__14_,r_484__13_,r_484__12_,r_484__11_,
  r_484__10_,r_484__9_,r_484__8_,r_484__7_,r_484__6_,r_484__5_,r_484__4_,r_484__3_,
  r_484__2_,r_484__1_,r_484__0_,r_485__63_,r_485__62_,r_485__61_,r_485__60_,r_485__59_,
  r_485__58_,r_485__57_,r_485__56_,r_485__55_,r_485__54_,r_485__53_,r_485__52_,
  r_485__51_,r_485__50_,r_485__49_,r_485__48_,r_485__47_,r_485__46_,r_485__45_,
  r_485__44_,r_485__43_,r_485__42_,r_485__41_,r_485__40_,r_485__39_,r_485__38_,
  r_485__37_,r_485__36_,r_485__35_,r_485__34_,r_485__33_,r_485__32_,r_485__31_,r_485__30_,
  r_485__29_,r_485__28_,r_485__27_,r_485__26_,r_485__25_,r_485__24_,r_485__23_,
  r_485__22_,r_485__21_,r_485__20_,r_485__19_,r_485__18_,r_485__17_,r_485__16_,
  r_485__15_,r_485__14_,r_485__13_,r_485__12_,r_485__11_,r_485__10_,r_485__9_,r_485__8_,
  r_485__7_,r_485__6_,r_485__5_,r_485__4_,r_485__3_,r_485__2_,r_485__1_,r_485__0_,
  r_486__63_,r_486__62_,r_486__61_,r_486__60_,r_486__59_,r_486__58_,r_486__57_,
  r_486__56_,r_486__55_,r_486__54_,r_486__53_,r_486__52_,r_486__51_,r_486__50_,
  r_486__49_,r_486__48_,r_486__47_,r_486__46_,r_486__45_,r_486__44_,r_486__43_,r_486__42_,
  r_486__41_,r_486__40_,r_486__39_,r_486__38_,r_486__37_,r_486__36_,r_486__35_,
  r_486__34_,r_486__33_,r_486__32_,r_486__31_,r_486__30_,r_486__29_,r_486__28_,
  r_486__27_,r_486__26_,r_486__25_,r_486__24_,r_486__23_,r_486__22_,r_486__21_,
  r_486__20_,r_486__19_,r_486__18_,r_486__17_,r_486__16_,r_486__15_,r_486__14_,r_486__13_,
  r_486__12_,r_486__11_,r_486__10_,r_486__9_,r_486__8_,r_486__7_,r_486__6_,
  r_486__5_,r_486__4_,r_486__3_,r_486__2_,r_486__1_,r_486__0_,r_487__63_,r_487__62_,
  r_487__61_,r_487__60_,r_487__59_,r_487__58_,r_487__57_,r_487__56_,r_487__55_,
  r_487__54_,r_487__53_,r_487__52_,r_487__51_,r_487__50_,r_487__49_,r_487__48_,r_487__47_,
  r_487__46_,r_487__45_,r_487__44_,r_487__43_,r_487__42_,r_487__41_,r_487__40_,
  r_487__39_,r_487__38_,r_487__37_,r_487__36_,r_487__35_,r_487__34_,r_487__33_,
  r_487__32_,r_487__31_,r_487__30_,r_487__29_,r_487__28_,r_487__27_,r_487__26_,
  r_487__25_,r_487__24_,r_487__23_,r_487__22_,r_487__21_,r_487__20_,r_487__19_,r_487__18_,
  r_487__17_,r_487__16_,r_487__15_,r_487__14_,r_487__13_,r_487__12_,r_487__11_,
  r_487__10_,r_487__9_,r_487__8_,r_487__7_,r_487__6_,r_487__5_,r_487__4_,r_487__3_,
  r_487__2_,r_487__1_,r_487__0_,r_488__63_,r_488__62_,r_488__61_,r_488__60_,
  r_488__59_,r_488__58_,r_488__57_,r_488__56_,r_488__55_,r_488__54_,r_488__53_,r_488__52_,
  r_488__51_,r_488__50_,r_488__49_,r_488__48_,r_488__47_,r_488__46_,r_488__45_,
  r_488__44_,r_488__43_,r_488__42_,r_488__41_,r_488__40_,r_488__39_,r_488__38_,
  r_488__37_,r_488__36_,r_488__35_,r_488__34_,r_488__33_,r_488__32_,r_488__31_,r_488__30_,
  r_488__29_,r_488__28_,r_488__27_,r_488__26_,r_488__25_,r_488__24_,r_488__23_,
  r_488__22_,r_488__21_,r_488__20_,r_488__19_,r_488__18_,r_488__17_,r_488__16_,
  r_488__15_,r_488__14_,r_488__13_,r_488__12_,r_488__11_,r_488__10_,r_488__9_,r_488__8_,
  r_488__7_,r_488__6_,r_488__5_,r_488__4_,r_488__3_,r_488__2_,r_488__1_,r_488__0_,
  r_489__63_,r_489__62_,r_489__61_,r_489__60_,r_489__59_,r_489__58_,r_489__57_,
  r_489__56_,r_489__55_,r_489__54_,r_489__53_,r_489__52_,r_489__51_,r_489__50_,
  r_489__49_,r_489__48_,r_489__47_,r_489__46_,r_489__45_,r_489__44_,r_489__43_,
  r_489__42_,r_489__41_,r_489__40_,r_489__39_,r_489__38_,r_489__37_,r_489__36_,r_489__35_,
  r_489__34_,r_489__33_,r_489__32_,r_489__31_,r_489__30_,r_489__29_,r_489__28_,
  r_489__27_,r_489__26_,r_489__25_,r_489__24_,r_489__23_,r_489__22_,r_489__21_,
  r_489__20_,r_489__19_,r_489__18_,r_489__17_,r_489__16_,r_489__15_,r_489__14_,
  r_489__13_,r_489__12_,r_489__11_,r_489__10_,r_489__9_,r_489__8_,r_489__7_,r_489__6_,
  r_489__5_,r_489__4_,r_489__3_,r_489__2_,r_489__1_,r_489__0_,r_490__63_,r_490__62_,
  r_490__61_,r_490__60_,r_490__59_,r_490__58_,r_490__57_,r_490__56_,r_490__55_,
  r_490__54_,r_490__53_,r_490__52_,r_490__51_,r_490__50_,r_490__49_,r_490__48_,
  r_490__47_,r_490__46_,r_490__45_,r_490__44_,r_490__43_,r_490__42_,r_490__41_,r_490__40_,
  r_490__39_,r_490__38_,r_490__37_,r_490__36_,r_490__35_,r_490__34_,r_490__33_,
  r_490__32_,r_490__31_,r_490__30_,r_490__29_,r_490__28_,r_490__27_,r_490__26_,
  r_490__25_,r_490__24_,r_490__23_,r_490__22_,r_490__21_,r_490__20_,r_490__19_,r_490__18_,
  r_490__17_,r_490__16_,r_490__15_,r_490__14_,r_490__13_,r_490__12_,r_490__11_,
  r_490__10_,r_490__9_,r_490__8_,r_490__7_,r_490__6_,r_490__5_,r_490__4_,r_490__3_,
  r_490__2_,r_490__1_,r_490__0_,r_491__63_,r_491__62_,r_491__61_,r_491__60_,
  r_491__59_,r_491__58_,r_491__57_,r_491__56_,r_491__55_,r_491__54_,r_491__53_,r_491__52_,
  r_491__51_,r_491__50_,r_491__49_,r_491__48_,r_491__47_,r_491__46_,r_491__45_,
  r_491__44_,r_491__43_,r_491__42_,r_491__41_,r_491__40_,r_491__39_,r_491__38_,
  r_491__37_,r_491__36_,r_491__35_,r_491__34_,r_491__33_,r_491__32_,r_491__31_,
  r_491__30_,r_491__29_,r_491__28_,r_491__27_,r_491__26_,r_491__25_,r_491__24_,r_491__23_,
  r_491__22_,r_491__21_,r_491__20_,r_491__19_,r_491__18_,r_491__17_,r_491__16_,
  r_491__15_,r_491__14_,r_491__13_,r_491__12_,r_491__11_,r_491__10_,r_491__9_,
  r_491__8_,r_491__7_,r_491__6_,r_491__5_,r_491__4_,r_491__3_,r_491__2_,r_491__1_,
  r_491__0_,r_492__63_,r_492__62_,r_492__61_,r_492__60_,r_492__59_,r_492__58_,r_492__57_,
  r_492__56_,r_492__55_,r_492__54_,r_492__53_,r_492__52_,r_492__51_,r_492__50_,
  r_492__49_,r_492__48_,r_492__47_,r_492__46_,r_492__45_,r_492__44_,r_492__43_,
  r_492__42_,r_492__41_,r_492__40_,r_492__39_,r_492__38_,r_492__37_,r_492__36_,
  r_492__35_,r_492__34_,r_492__33_,r_492__32_,r_492__31_,r_492__30_,r_492__29_,r_492__28_,
  r_492__27_,r_492__26_,r_492__25_,r_492__24_,r_492__23_,r_492__22_,r_492__21_,
  r_492__20_,r_492__19_,r_492__18_,r_492__17_,r_492__16_,r_492__15_,r_492__14_,
  r_492__13_,r_492__12_,r_492__11_,r_492__10_,r_492__9_,r_492__8_,r_492__7_,r_492__6_,
  r_492__5_,r_492__4_,r_492__3_,r_492__2_,r_492__1_,r_492__0_,r_493__63_,r_493__62_,
  r_493__61_,r_493__60_,r_493__59_,r_493__58_,r_493__57_,r_493__56_,r_493__55_,
  r_493__54_,r_493__53_,r_493__52_,r_493__51_,r_493__50_,r_493__49_,r_493__48_,
  r_493__47_,r_493__46_,r_493__45_,r_493__44_,r_493__43_,r_493__42_,r_493__41_,r_493__40_,
  r_493__39_,r_493__38_,r_493__37_,r_493__36_,r_493__35_,r_493__34_,r_493__33_,
  r_493__32_,r_493__31_,r_493__30_,r_493__29_,r_493__28_,r_493__27_,r_493__26_,
  r_493__25_,r_493__24_,r_493__23_,r_493__22_,r_493__21_,r_493__20_,r_493__19_,
  r_493__18_,r_493__17_,r_493__16_,r_493__15_,r_493__14_,r_493__13_,r_493__12_,r_493__11_,
  r_493__10_,r_493__9_,r_493__8_,r_493__7_,r_493__6_,r_493__5_,r_493__4_,r_493__3_,
  r_493__2_,r_493__1_,r_493__0_,r_494__63_,r_494__62_,r_494__61_,r_494__60_,
  r_494__59_,r_494__58_,r_494__57_,r_494__56_,r_494__55_,r_494__54_,r_494__53_,
  r_494__52_,r_494__51_,r_494__50_,r_494__49_,r_494__48_,r_494__47_,r_494__46_,r_494__45_,
  r_494__44_,r_494__43_,r_494__42_,r_494__41_,r_494__40_,r_494__39_,r_494__38_,
  r_494__37_,r_494__36_,r_494__35_,r_494__34_,r_494__33_,r_494__32_,r_494__31_,
  r_494__30_,r_494__29_,r_494__28_,r_494__27_,r_494__26_,r_494__25_,r_494__24_,
  r_494__23_,r_494__22_,r_494__21_,r_494__20_,r_494__19_,r_494__18_,r_494__17_,r_494__16_,
  r_494__15_,r_494__14_,r_494__13_,r_494__12_,r_494__11_,r_494__10_,r_494__9_,
  r_494__8_,r_494__7_,r_494__6_,r_494__5_,r_494__4_,r_494__3_,r_494__2_,r_494__1_,
  r_494__0_,r_495__63_,r_495__62_,r_495__61_,r_495__60_,r_495__59_,r_495__58_,
  r_495__57_,r_495__56_,r_495__55_,r_495__54_,r_495__53_,r_495__52_,r_495__51_,r_495__50_,
  r_495__49_,r_495__48_,r_495__47_,r_495__46_,r_495__45_,r_495__44_,r_495__43_,
  r_495__42_,r_495__41_,r_495__40_,r_495__39_,r_495__38_,r_495__37_,r_495__36_,
  r_495__35_,r_495__34_,r_495__33_,r_495__32_,r_495__31_,r_495__30_,r_495__29_,r_495__28_,
  r_495__27_,r_495__26_,r_495__25_,r_495__24_,r_495__23_,r_495__22_,r_495__21_,
  r_495__20_,r_495__19_,r_495__18_,r_495__17_,r_495__16_,r_495__15_,r_495__14_,
  r_495__13_,r_495__12_,r_495__11_,r_495__10_,r_495__9_,r_495__8_,r_495__7_,r_495__6_,
  r_495__5_,r_495__4_,r_495__3_,r_495__2_,r_495__1_,r_495__0_,r_496__63_,r_496__62_,
  r_496__61_,r_496__60_,r_496__59_,r_496__58_,r_496__57_,r_496__56_,r_496__55_,
  r_496__54_,r_496__53_,r_496__52_,r_496__51_,r_496__50_,r_496__49_,r_496__48_,
  r_496__47_,r_496__46_,r_496__45_,r_496__44_,r_496__43_,r_496__42_,r_496__41_,
  r_496__40_,r_496__39_,r_496__38_,r_496__37_,r_496__36_,r_496__35_,r_496__34_,r_496__33_,
  r_496__32_,r_496__31_,r_496__30_,r_496__29_,r_496__28_,r_496__27_,r_496__26_,
  r_496__25_,r_496__24_,r_496__23_,r_496__22_,r_496__21_,r_496__20_,r_496__19_,
  r_496__18_,r_496__17_,r_496__16_,r_496__15_,r_496__14_,r_496__13_,r_496__12_,
  r_496__11_,r_496__10_,r_496__9_,r_496__8_,r_496__7_,r_496__6_,r_496__5_,r_496__4_,
  r_496__3_,r_496__2_,r_496__1_,r_496__0_,r_497__63_,r_497__62_,r_497__61_,r_497__60_,
  r_497__59_,r_497__58_,r_497__57_,r_497__56_,r_497__55_,r_497__54_,r_497__53_,
  r_497__52_,r_497__51_,r_497__50_,r_497__49_,r_497__48_,r_497__47_,r_497__46_,
  r_497__45_,r_497__44_,r_497__43_,r_497__42_,r_497__41_,r_497__40_,r_497__39_,r_497__38_,
  r_497__37_,r_497__36_,r_497__35_,r_497__34_,r_497__33_,r_497__32_,r_497__31_,
  r_497__30_,r_497__29_,r_497__28_,r_497__27_,r_497__26_,r_497__25_,r_497__24_,
  r_497__23_,r_497__22_,r_497__21_,r_497__20_,r_497__19_,r_497__18_,r_497__17_,r_497__16_,
  r_497__15_,r_497__14_,r_497__13_,r_497__12_,r_497__11_,r_497__10_,r_497__9_,
  r_497__8_,r_497__7_,r_497__6_,r_497__5_,r_497__4_,r_497__3_,r_497__2_,r_497__1_,
  r_497__0_,r_498__63_,r_498__62_,r_498__61_,r_498__60_,r_498__59_,r_498__58_,
  r_498__57_,r_498__56_,r_498__55_,r_498__54_,r_498__53_,r_498__52_,r_498__51_,r_498__50_,
  r_498__49_,r_498__48_,r_498__47_,r_498__46_,r_498__45_,r_498__44_,r_498__43_,
  r_498__42_,r_498__41_,r_498__40_,r_498__39_,r_498__38_,r_498__37_,r_498__36_,
  r_498__35_,r_498__34_,r_498__33_,r_498__32_,r_498__31_,r_498__30_,r_498__29_,
  r_498__28_,r_498__27_,r_498__26_,r_498__25_,r_498__24_,r_498__23_,r_498__22_,r_498__21_,
  r_498__20_,r_498__19_,r_498__18_,r_498__17_,r_498__16_,r_498__15_,r_498__14_,
  r_498__13_,r_498__12_,r_498__11_,r_498__10_,r_498__9_,r_498__8_,r_498__7_,r_498__6_,
  r_498__5_,r_498__4_,r_498__3_,r_498__2_,r_498__1_,r_498__0_,r_499__63_,
  r_499__62_,r_499__61_,r_499__60_,r_499__59_,r_499__58_,r_499__57_,r_499__56_,r_499__55_,
  r_499__54_,r_499__53_,r_499__52_,r_499__51_,r_499__50_,r_499__49_,r_499__48_,
  r_499__47_,r_499__46_,r_499__45_,r_499__44_,r_499__43_,r_499__42_,r_499__41_,
  r_499__40_,r_499__39_,r_499__38_,r_499__37_,r_499__36_,r_499__35_,r_499__34_,
  r_499__33_,r_499__32_,r_499__31_,r_499__30_,r_499__29_,r_499__28_,r_499__27_,r_499__26_,
  r_499__25_,r_499__24_,r_499__23_,r_499__22_,r_499__21_,r_499__20_,r_499__19_,
  r_499__18_,r_499__17_,r_499__16_,r_499__15_,r_499__14_,r_499__13_,r_499__12_,
  r_499__11_,r_499__10_,r_499__9_,r_499__8_,r_499__7_,r_499__6_,r_499__5_,r_499__4_,
  r_499__3_,r_499__2_,r_499__1_,r_499__0_,r_500__63_,r_500__62_,r_500__61_,r_500__60_,
  r_500__59_,r_500__58_,r_500__57_,r_500__56_,r_500__55_,r_500__54_,r_500__53_,
  r_500__52_,r_500__51_,r_500__50_,r_500__49_,r_500__48_,r_500__47_,r_500__46_,
  r_500__45_,r_500__44_,r_500__43_,r_500__42_,r_500__41_,r_500__40_,r_500__39_,r_500__38_,
  r_500__37_,r_500__36_,r_500__35_,r_500__34_,r_500__33_,r_500__32_,r_500__31_,
  r_500__30_,r_500__29_,r_500__28_,r_500__27_,r_500__26_,r_500__25_,r_500__24_,
  r_500__23_,r_500__22_,r_500__21_,r_500__20_,r_500__19_,r_500__18_,r_500__17_,
  r_500__16_,r_500__15_,r_500__14_,r_500__13_,r_500__12_,r_500__11_,r_500__10_,r_500__9_,
  r_500__8_,r_500__7_,r_500__6_,r_500__5_,r_500__4_,r_500__3_,r_500__2_,r_500__1_,
  r_500__0_,r_501__63_,r_501__62_,r_501__61_,r_501__60_,r_501__59_,r_501__58_,
  r_501__57_,r_501__56_,r_501__55_,r_501__54_,r_501__53_,r_501__52_,r_501__51_,
  r_501__50_,r_501__49_,r_501__48_,r_501__47_,r_501__46_,r_501__45_,r_501__44_,r_501__43_,
  r_501__42_,r_501__41_,r_501__40_,r_501__39_,r_501__38_,r_501__37_,r_501__36_,
  r_501__35_,r_501__34_,r_501__33_,r_501__32_,r_501__31_,r_501__30_,r_501__29_,
  r_501__28_,r_501__27_,r_501__26_,r_501__25_,r_501__24_,r_501__23_,r_501__22_,
  r_501__21_,r_501__20_,r_501__19_,r_501__18_,r_501__17_,r_501__16_,r_501__15_,r_501__14_,
  r_501__13_,r_501__12_,r_501__11_,r_501__10_,r_501__9_,r_501__8_,r_501__7_,
  r_501__6_,r_501__5_,r_501__4_,r_501__3_,r_501__2_,r_501__1_,r_501__0_,r_502__63_,
  r_502__62_,r_502__61_,r_502__60_,r_502__59_,r_502__58_,r_502__57_,r_502__56_,
  r_502__55_,r_502__54_,r_502__53_,r_502__52_,r_502__51_,r_502__50_,r_502__49_,r_502__48_,
  r_502__47_,r_502__46_,r_502__45_,r_502__44_,r_502__43_,r_502__42_,r_502__41_,
  r_502__40_,r_502__39_,r_502__38_,r_502__37_,r_502__36_,r_502__35_,r_502__34_,
  r_502__33_,r_502__32_,r_502__31_,r_502__30_,r_502__29_,r_502__28_,r_502__27_,r_502__26_,
  r_502__25_,r_502__24_,r_502__23_,r_502__22_,r_502__21_,r_502__20_,r_502__19_,
  r_502__18_,r_502__17_,r_502__16_,r_502__15_,r_502__14_,r_502__13_,r_502__12_,
  r_502__11_,r_502__10_,r_502__9_,r_502__8_,r_502__7_,r_502__6_,r_502__5_,r_502__4_,
  r_502__3_,r_502__2_,r_502__1_,r_502__0_,r_503__63_,r_503__62_,r_503__61_,r_503__60_,
  r_503__59_,r_503__58_,r_503__57_,r_503__56_,r_503__55_,r_503__54_,r_503__53_,
  r_503__52_,r_503__51_,r_503__50_,r_503__49_,r_503__48_,r_503__47_,r_503__46_,
  r_503__45_,r_503__44_,r_503__43_,r_503__42_,r_503__41_,r_503__40_,r_503__39_,
  r_503__38_,r_503__37_,r_503__36_,r_503__35_,r_503__34_,r_503__33_,r_503__32_,r_503__31_,
  r_503__30_,r_503__29_,r_503__28_,r_503__27_,r_503__26_,r_503__25_,r_503__24_,
  r_503__23_,r_503__22_,r_503__21_,r_503__20_,r_503__19_,r_503__18_,r_503__17_,
  r_503__16_,r_503__15_,r_503__14_,r_503__13_,r_503__12_,r_503__11_,r_503__10_,r_503__9_,
  r_503__8_,r_503__7_,r_503__6_,r_503__5_,r_503__4_,r_503__3_,r_503__2_,r_503__1_,
  r_503__0_,r_504__63_,r_504__62_,r_504__61_,r_504__60_,r_504__59_,r_504__58_,
  r_504__57_,r_504__56_,r_504__55_,r_504__54_,r_504__53_,r_504__52_,r_504__51_,
  r_504__50_,r_504__49_,r_504__48_,r_504__47_,r_504__46_,r_504__45_,r_504__44_,
  r_504__43_,r_504__42_,r_504__41_,r_504__40_,r_504__39_,r_504__38_,r_504__37_,r_504__36_,
  r_504__35_,r_504__34_,r_504__33_,r_504__32_,r_504__31_,r_504__30_,r_504__29_,
  r_504__28_,r_504__27_,r_504__26_,r_504__25_,r_504__24_,r_504__23_,r_504__22_,
  r_504__21_,r_504__20_,r_504__19_,r_504__18_,r_504__17_,r_504__16_,r_504__15_,r_504__14_,
  r_504__13_,r_504__12_,r_504__11_,r_504__10_,r_504__9_,r_504__8_,r_504__7_,
  r_504__6_,r_504__5_,r_504__4_,r_504__3_,r_504__2_,r_504__1_,r_504__0_,r_505__63_,
  r_505__62_,r_505__61_,r_505__60_,r_505__59_,r_505__58_,r_505__57_,r_505__56_,
  r_505__55_,r_505__54_,r_505__53_,r_505__52_,r_505__51_,r_505__50_,r_505__49_,r_505__48_,
  r_505__47_,r_505__46_,r_505__45_,r_505__44_,r_505__43_,r_505__42_,r_505__41_,
  r_505__40_,r_505__39_,r_505__38_,r_505__37_,r_505__36_,r_505__35_,r_505__34_,
  r_505__33_,r_505__32_,r_505__31_,r_505__30_,r_505__29_,r_505__28_,r_505__27_,
  r_505__26_,r_505__25_,r_505__24_,r_505__23_,r_505__22_,r_505__21_,r_505__20_,r_505__19_,
  r_505__18_,r_505__17_,r_505__16_,r_505__15_,r_505__14_,r_505__13_,r_505__12_,
  r_505__11_,r_505__10_,r_505__9_,r_505__8_,r_505__7_,r_505__6_,r_505__5_,r_505__4_,
  r_505__3_,r_505__2_,r_505__1_,r_505__0_,r_506__63_,r_506__62_,r_506__61_,
  r_506__60_,r_506__59_,r_506__58_,r_506__57_,r_506__56_,r_506__55_,r_506__54_,r_506__53_,
  r_506__52_,r_506__51_,r_506__50_,r_506__49_,r_506__48_,r_506__47_,r_506__46_,
  r_506__45_,r_506__44_,r_506__43_,r_506__42_,r_506__41_,r_506__40_,r_506__39_,
  r_506__38_,r_506__37_,r_506__36_,r_506__35_,r_506__34_,r_506__33_,r_506__32_,
  r_506__31_,r_506__30_,r_506__29_,r_506__28_,r_506__27_,r_506__26_,r_506__25_,r_506__24_,
  r_506__23_,r_506__22_,r_506__21_,r_506__20_,r_506__19_,r_506__18_,r_506__17_,
  r_506__16_,r_506__15_,r_506__14_,r_506__13_,r_506__12_,r_506__11_,r_506__10_,
  r_506__9_,r_506__8_,r_506__7_,r_506__6_,r_506__5_,r_506__4_,r_506__3_,r_506__2_,
  r_506__1_,r_506__0_,r_507__63_,r_507__62_,r_507__61_,r_507__60_,r_507__59_,r_507__58_,
  r_507__57_,r_507__56_,r_507__55_,r_507__54_,r_507__53_,r_507__52_,r_507__51_,
  r_507__50_,r_507__49_,r_507__48_,r_507__47_,r_507__46_,r_507__45_,r_507__44_,
  r_507__43_,r_507__42_,r_507__41_,r_507__40_,r_507__39_,r_507__38_,r_507__37_,r_507__36_,
  r_507__35_,r_507__34_,r_507__33_,r_507__32_,r_507__31_,r_507__30_,r_507__29_,
  r_507__28_,r_507__27_,r_507__26_,r_507__25_,r_507__24_,r_507__23_,r_507__22_,
  r_507__21_,r_507__20_,r_507__19_,r_507__18_,r_507__17_,r_507__16_,r_507__15_,
  r_507__14_,r_507__13_,r_507__12_,r_507__11_,r_507__10_,r_507__9_,r_507__8_,r_507__7_,
  r_507__6_,r_507__5_,r_507__4_,r_507__3_,r_507__2_,r_507__1_,r_507__0_,r_508__63_,
  r_508__62_,r_508__61_,r_508__60_,r_508__59_,r_508__58_,r_508__57_,r_508__56_,
  r_508__55_,r_508__54_,r_508__53_,r_508__52_,r_508__51_,r_508__50_,r_508__49_,
  r_508__48_,r_508__47_,r_508__46_,r_508__45_,r_508__44_,r_508__43_,r_508__42_,r_508__41_,
  r_508__40_,r_508__39_,r_508__38_,r_508__37_,r_508__36_,r_508__35_,r_508__34_,
  r_508__33_,r_508__32_,r_508__31_,r_508__30_,r_508__29_,r_508__28_,r_508__27_,
  r_508__26_,r_508__25_,r_508__24_,r_508__23_,r_508__22_,r_508__21_,r_508__20_,
  r_508__19_,r_508__18_,r_508__17_,r_508__16_,r_508__15_,r_508__14_,r_508__13_,r_508__12_,
  r_508__11_,r_508__10_,r_508__9_,r_508__8_,r_508__7_,r_508__6_,r_508__5_,r_508__4_,
  r_508__3_,r_508__2_,r_508__1_,r_508__0_,r_509__63_,r_509__62_,r_509__61_,
  r_509__60_,r_509__59_,r_509__58_,r_509__57_,r_509__56_,r_509__55_,r_509__54_,
  r_509__53_,r_509__52_,r_509__51_,r_509__50_,r_509__49_,r_509__48_,r_509__47_,r_509__46_,
  r_509__45_,r_509__44_,r_509__43_,r_509__42_,r_509__41_,r_509__40_,r_509__39_,
  r_509__38_,r_509__37_,r_509__36_,r_509__35_,r_509__34_,r_509__33_,r_509__32_,
  r_509__31_,r_509__30_,r_509__29_,r_509__28_,r_509__27_,r_509__26_,r_509__25_,r_509__24_,
  r_509__23_,r_509__22_,r_509__21_,r_509__20_,r_509__19_,r_509__18_,r_509__17_,
  r_509__16_,r_509__15_,r_509__14_,r_509__13_,r_509__12_,r_509__11_,r_509__10_,
  r_509__9_,r_509__8_,r_509__7_,r_509__6_,r_509__5_,r_509__4_,r_509__3_,r_509__2_,
  r_509__1_,r_509__0_,r_510__63_,r_510__62_,r_510__61_,r_510__60_,r_510__59_,r_510__58_,
  r_510__57_,r_510__56_,r_510__55_,r_510__54_,r_510__53_,r_510__52_,r_510__51_,
  r_510__50_,r_510__49_,r_510__48_,r_510__47_,r_510__46_,r_510__45_,r_510__44_,
  r_510__43_,r_510__42_,r_510__41_,r_510__40_,r_510__39_,r_510__38_,r_510__37_,
  r_510__36_,r_510__35_,r_510__34_,r_510__33_,r_510__32_,r_510__31_,r_510__30_,r_510__29_,
  r_510__28_,r_510__27_,r_510__26_,r_510__25_,r_510__24_,r_510__23_,r_510__22_,
  r_510__21_,r_510__20_,r_510__19_,r_510__18_,r_510__17_,r_510__16_,r_510__15_,
  r_510__14_,r_510__13_,r_510__12_,r_510__11_,r_510__10_,r_510__9_,r_510__8_,r_510__7_,
  r_510__6_,r_510__5_,r_510__4_,r_510__3_,r_510__2_,r_510__1_,r_510__0_,r_511__63_,
  r_511__62_,r_511__61_,r_511__60_,r_511__59_,r_511__58_,r_511__57_,r_511__56_,
  r_511__55_,r_511__54_,r_511__53_,r_511__52_,r_511__51_,r_511__50_,r_511__49_,
  r_511__48_,r_511__47_,r_511__46_,r_511__45_,r_511__44_,r_511__43_,r_511__42_,
  r_511__41_,r_511__40_,r_511__39_,r_511__38_,r_511__37_,r_511__36_,r_511__35_,r_511__34_,
  r_511__33_,r_511__32_,r_511__31_,r_511__30_,r_511__29_,r_511__28_,r_511__27_,
  r_511__26_,r_511__25_,r_511__24_,r_511__23_,r_511__22_,r_511__21_,r_511__20_,
  r_511__19_,r_511__18_,r_511__17_,r_511__16_,r_511__15_,r_511__14_,r_511__13_,r_511__12_,
  r_511__11_,r_511__10_,r_511__9_,r_511__8_,r_511__7_,r_511__6_,r_511__5_,
  r_511__4_,r_511__3_,r_511__2_,r_511__1_,r_511__0_;
  assign N1024 = sel_i[1] & sel_i[0];
  assign N1026 = N1025 & N1028;
  assign N1029 = sel_i[3] & sel_i[2];
  assign N1031 = N1030 & N1033;
  assign N1034 = sel_i[5] & sel_i[4];
  assign N1036 = N1035 & N1038;
  assign N1039 = sel_i[7] & sel_i[6];
  assign N1041 = N1040 & N1043;
  assign N1044 = sel_i[9] & sel_i[8];
  assign N1046 = N1045 & N1048;
  assign N1049 = sel_i[11] & sel_i[10];
  assign N1051 = N1050 & N1053;
  assign N1054 = sel_i[13] & sel_i[12];
  assign N1056 = N1055 & N1058;
  assign N1059 = sel_i[15] & sel_i[14];
  assign N1061 = N1060 & N1063;
  assign N1064 = sel_i[17] & sel_i[16];
  assign N1066 = N1065 & N1068;
  assign N1069 = sel_i[19] & sel_i[18];
  assign N1071 = N1070 & N1073;
  assign N1074 = sel_i[21] & sel_i[20];
  assign N1076 = N1075 & N1078;
  assign N1079 = sel_i[23] & sel_i[22];
  assign N1081 = N1080 & N1083;
  assign N1084 = sel_i[25] & sel_i[24];
  assign N1086 = N1085 & N1088;
  assign N1089 = sel_i[27] & sel_i[26];
  assign N1091 = N1090 & N1093;
  assign N1094 = sel_i[29] & sel_i[28];
  assign N1096 = N1095 & N1098;
  assign N1099 = sel_i[31] & sel_i[30];
  assign N1101 = N1100 & N1103;
  assign N1104 = sel_i[33] & sel_i[32];
  assign N1106 = N1105 & N1108;
  assign N1109 = sel_i[35] & sel_i[34];
  assign N1111 = N1110 & N1113;
  assign N1114 = sel_i[37] & sel_i[36];
  assign N1116 = N1115 & N1118;
  assign N1119 = sel_i[39] & sel_i[38];
  assign N1121 = N1120 & N1123;
  assign N1124 = sel_i[41] & sel_i[40];
  assign N1126 = N1125 & N1128;
  assign N1129 = sel_i[43] & sel_i[42];
  assign N1131 = N1130 & N1133;
  assign N1134 = sel_i[45] & sel_i[44];
  assign N1136 = N1135 & N1138;
  assign N1139 = sel_i[47] & sel_i[46];
  assign N1141 = N1140 & N1143;
  assign N1144 = sel_i[49] & sel_i[48];
  assign N1146 = N1145 & N1148;
  assign N1149 = sel_i[51] & sel_i[50];
  assign N1151 = N1150 & N1153;
  assign N1154 = sel_i[53] & sel_i[52];
  assign N1156 = N1155 & N1158;
  assign N1159 = sel_i[55] & sel_i[54];
  assign N1161 = N1160 & N1163;
  assign N1164 = sel_i[57] & sel_i[56];
  assign N1166 = N1165 & N1168;
  assign N1169 = sel_i[59] & sel_i[58];
  assign N1171 = N1170 & N1173;
  assign N1174 = sel_i[61] & sel_i[60];
  assign N1176 = N1175 & N1178;
  assign N1179 = sel_i[63] & sel_i[62];
  assign N1181 = N1180 & N1183;
  assign N1184 = sel_i[65] & sel_i[64];
  assign N1186 = N1185 & N1188;
  assign N1189 = sel_i[67] & sel_i[66];
  assign N1191 = N1190 & N1193;
  assign N1194 = sel_i[69] & sel_i[68];
  assign N1196 = N1195 & N1198;
  assign N1199 = sel_i[71] & sel_i[70];
  assign N1201 = N1200 & N1203;
  assign N1204 = sel_i[73] & sel_i[72];
  assign N1206 = N1205 & N1208;
  assign N1209 = sel_i[75] & sel_i[74];
  assign N1211 = N1210 & N1213;
  assign N1214 = sel_i[77] & sel_i[76];
  assign N1216 = N1215 & N1218;
  assign N1219 = sel_i[79] & sel_i[78];
  assign N1221 = N1220 & N1223;
  assign N1224 = sel_i[81] & sel_i[80];
  assign N1226 = N1225 & N1228;
  assign N1229 = sel_i[83] & sel_i[82];
  assign N1231 = N1230 & N1233;
  assign N1234 = sel_i[85] & sel_i[84];
  assign N1236 = N1235 & N1238;
  assign N1239 = sel_i[87] & sel_i[86];
  assign N1241 = N1240 & N1243;
  assign N1244 = sel_i[89] & sel_i[88];
  assign N1246 = N1245 & N1248;
  assign N1249 = sel_i[91] & sel_i[90];
  assign N1251 = N1250 & N1253;
  assign N1254 = sel_i[93] & sel_i[92];
  assign N1256 = N1255 & N1258;
  assign N1259 = sel_i[95] & sel_i[94];
  assign N1261 = N1260 & N1263;
  assign N1264 = sel_i[97] & sel_i[96];
  assign N1266 = N1265 & N1268;
  assign N1269 = sel_i[99] & sel_i[98];
  assign N1271 = N1270 & N1273;
  assign N1274 = sel_i[101] & sel_i[100];
  assign N1276 = N1275 & N1278;
  assign N1279 = sel_i[103] & sel_i[102];
  assign N1281 = N1280 & N1283;
  assign N1284 = sel_i[105] & sel_i[104];
  assign N1286 = N1285 & N1288;
  assign N1289 = sel_i[107] & sel_i[106];
  assign N1291 = N1290 & N1293;
  assign N1294 = sel_i[109] & sel_i[108];
  assign N1296 = N1295 & N1298;
  assign N1299 = sel_i[111] & sel_i[110];
  assign N1301 = N1300 & N1303;
  assign N1304 = sel_i[113] & sel_i[112];
  assign N1306 = N1305 & N1308;
  assign N1309 = sel_i[115] & sel_i[114];
  assign N1311 = N1310 & N1313;
  assign N1314 = sel_i[117] & sel_i[116];
  assign N1316 = N1315 & N1318;
  assign N1319 = sel_i[119] & sel_i[118];
  assign N1321 = N1320 & N1323;
  assign N1324 = sel_i[121] & sel_i[120];
  assign N1326 = N1325 & N1328;
  assign N1329 = sel_i[123] & sel_i[122];
  assign N1331 = N1330 & N1333;
  assign N1334 = sel_i[125] & sel_i[124];
  assign N1336 = N1335 & N1338;
  assign N1339 = sel_i[127] & sel_i[126];
  assign N1341 = N1340 & N1343;
  assign N1344 = sel_i[129] & sel_i[128];
  assign N1346 = N1345 & N1348;
  assign N1349 = sel_i[131] & sel_i[130];
  assign N1351 = N1350 & N1353;
  assign N1354 = sel_i[133] & sel_i[132];
  assign N1356 = N1355 & N1358;
  assign N1359 = sel_i[135] & sel_i[134];
  assign N1361 = N1360 & N1363;
  assign N1364 = sel_i[137] & sel_i[136];
  assign N1366 = N1365 & N1368;
  assign N1369 = sel_i[139] & sel_i[138];
  assign N1371 = N1370 & N1373;
  assign N1374 = sel_i[141] & sel_i[140];
  assign N1376 = N1375 & N1378;
  assign N1379 = sel_i[143] & sel_i[142];
  assign N1381 = N1380 & N1383;
  assign N1384 = sel_i[145] & sel_i[144];
  assign N1386 = N1385 & N1388;
  assign N1389 = sel_i[147] & sel_i[146];
  assign N1391 = N1390 & N1393;
  assign N1394 = sel_i[149] & sel_i[148];
  assign N1396 = N1395 & N1398;
  assign N1399 = sel_i[151] & sel_i[150];
  assign N1401 = N1400 & N1403;
  assign N1404 = sel_i[153] & sel_i[152];
  assign N1406 = N1405 & N1408;
  assign N1409 = sel_i[155] & sel_i[154];
  assign N1411 = N1410 & N1413;
  assign N1414 = sel_i[157] & sel_i[156];
  assign N1416 = N1415 & N1418;
  assign N1419 = sel_i[159] & sel_i[158];
  assign N1421 = N1420 & N1423;
  assign N1424 = sel_i[161] & sel_i[160];
  assign N1426 = N1425 & N1428;
  assign N1429 = sel_i[163] & sel_i[162];
  assign N1431 = N1430 & N1433;
  assign N1434 = sel_i[165] & sel_i[164];
  assign N1436 = N1435 & N1438;
  assign N1439 = sel_i[167] & sel_i[166];
  assign N1441 = N1440 & N1443;
  assign N1444 = sel_i[169] & sel_i[168];
  assign N1446 = N1445 & N1448;
  assign N1449 = sel_i[171] & sel_i[170];
  assign N1451 = N1450 & N1453;
  assign N1454 = sel_i[173] & sel_i[172];
  assign N1456 = N1455 & N1458;
  assign N1459 = sel_i[175] & sel_i[174];
  assign N1461 = N1460 & N1463;
  assign N1464 = sel_i[177] & sel_i[176];
  assign N1466 = N1465 & N1468;
  assign N1469 = sel_i[179] & sel_i[178];
  assign N1471 = N1470 & N1473;
  assign N1474 = sel_i[181] & sel_i[180];
  assign N1476 = N1475 & N1478;
  assign N1479 = sel_i[183] & sel_i[182];
  assign N1481 = N1480 & N1483;
  assign N1484 = sel_i[185] & sel_i[184];
  assign N1486 = N1485 & N1488;
  assign N1489 = sel_i[187] & sel_i[186];
  assign N1491 = N1490 & N1493;
  assign N1494 = sel_i[189] & sel_i[188];
  assign N1496 = N1495 & N1498;
  assign N1499 = sel_i[191] & sel_i[190];
  assign N1501 = N1500 & N1503;
  assign N1504 = sel_i[193] & sel_i[192];
  assign N1506 = N1505 & N1508;
  assign N1509 = sel_i[195] & sel_i[194];
  assign N1511 = N1510 & N1513;
  assign N1514 = sel_i[197] & sel_i[196];
  assign N1516 = N1515 & N1518;
  assign N1519 = sel_i[199] & sel_i[198];
  assign N1521 = N1520 & N1523;
  assign N1524 = sel_i[201] & sel_i[200];
  assign N1526 = N1525 & N1528;
  assign N1529 = sel_i[203] & sel_i[202];
  assign N1531 = N1530 & N1533;
  assign N1534 = sel_i[205] & sel_i[204];
  assign N1536 = N1535 & N1538;
  assign N1539 = sel_i[207] & sel_i[206];
  assign N1541 = N1540 & N1543;
  assign N1544 = sel_i[209] & sel_i[208];
  assign N1546 = N1545 & N1548;
  assign N1549 = sel_i[211] & sel_i[210];
  assign N1551 = N1550 & N1553;
  assign N1554 = sel_i[213] & sel_i[212];
  assign N1556 = N1555 & N1558;
  assign N1559 = sel_i[215] & sel_i[214];
  assign N1561 = N1560 & N1563;
  assign N1564 = sel_i[217] & sel_i[216];
  assign N1566 = N1565 & N1568;
  assign N1569 = sel_i[219] & sel_i[218];
  assign N1571 = N1570 & N1573;
  assign N1574 = sel_i[221] & sel_i[220];
  assign N1576 = N1575 & N1578;
  assign N1579 = sel_i[223] & sel_i[222];
  assign N1581 = N1580 & N1583;
  assign N1584 = sel_i[225] & sel_i[224];
  assign N1586 = N1585 & N1588;
  assign N1589 = sel_i[227] & sel_i[226];
  assign N1591 = N1590 & N1593;
  assign N1594 = sel_i[229] & sel_i[228];
  assign N1596 = N1595 & N1598;
  assign N1599 = sel_i[231] & sel_i[230];
  assign N1601 = N1600 & N1603;
  assign N1604 = sel_i[233] & sel_i[232];
  assign N1606 = N1605 & N1608;
  assign N1609 = sel_i[235] & sel_i[234];
  assign N1611 = N1610 & N1613;
  assign N1614 = sel_i[237] & sel_i[236];
  assign N1616 = N1615 & N1618;
  assign N1619 = sel_i[239] & sel_i[238];
  assign N1621 = N1620 & N1623;
  assign N1624 = sel_i[241] & sel_i[240];
  assign N1626 = N1625 & N1628;
  assign N1629 = sel_i[243] & sel_i[242];
  assign N1631 = N1630 & N1633;
  assign N1634 = sel_i[245] & sel_i[244];
  assign N1636 = N1635 & N1638;
  assign N1639 = sel_i[247] & sel_i[246];
  assign N1641 = N1640 & N1643;
  assign N1644 = sel_i[249] & sel_i[248];
  assign N1646 = N1645 & N1648;
  assign N1649 = sel_i[251] & sel_i[250];
  assign N1651 = N1650 & N1653;
  assign N1654 = sel_i[253] & sel_i[252];
  assign N1656 = N1655 & N1658;
  assign N1659 = sel_i[255] & sel_i[254];
  assign N1661 = N1660 & N1663;
  assign N1664 = sel_i[257] & sel_i[256];
  assign N1666 = N1665 & N1668;
  assign N1669 = sel_i[259] & sel_i[258];
  assign N1671 = N1670 & N1673;
  assign N1674 = sel_i[261] & sel_i[260];
  assign N1676 = N1675 & N1678;
  assign N1679 = sel_i[263] & sel_i[262];
  assign N1681 = N1680 & N1683;
  assign N1684 = sel_i[265] & sel_i[264];
  assign N1686 = N1685 & N1688;
  assign N1689 = sel_i[267] & sel_i[266];
  assign N1691 = N1690 & N1693;
  assign N1694 = sel_i[269] & sel_i[268];
  assign N1696 = N1695 & N1698;
  assign N1699 = sel_i[271] & sel_i[270];
  assign N1701 = N1700 & N1703;
  assign N1704 = sel_i[273] & sel_i[272];
  assign N1706 = N1705 & N1708;
  assign N1709 = sel_i[275] & sel_i[274];
  assign N1711 = N1710 & N1713;
  assign N1714 = sel_i[277] & sel_i[276];
  assign N1716 = N1715 & N1718;
  assign N1719 = sel_i[279] & sel_i[278];
  assign N1721 = N1720 & N1723;
  assign N1724 = sel_i[281] & sel_i[280];
  assign N1726 = N1725 & N1728;
  assign N1729 = sel_i[283] & sel_i[282];
  assign N1731 = N1730 & N1733;
  assign N1734 = sel_i[285] & sel_i[284];
  assign N1736 = N1735 & N1738;
  assign N1739 = sel_i[287] & sel_i[286];
  assign N1741 = N1740 & N1743;
  assign N1744 = sel_i[289] & sel_i[288];
  assign N1746 = N1745 & N1748;
  assign N1749 = sel_i[291] & sel_i[290];
  assign N1751 = N1750 & N1753;
  assign N1754 = sel_i[293] & sel_i[292];
  assign N1756 = N1755 & N1758;
  assign N1759 = sel_i[295] & sel_i[294];
  assign N1761 = N1760 & N1763;
  assign N1764 = sel_i[297] & sel_i[296];
  assign N1766 = N1765 & N1768;
  assign N1769 = sel_i[299] & sel_i[298];
  assign N1771 = N1770 & N1773;
  assign N1774 = sel_i[301] & sel_i[300];
  assign N1776 = N1775 & N1778;
  assign N1779 = sel_i[303] & sel_i[302];
  assign N1781 = N1780 & N1783;
  assign N1784 = sel_i[305] & sel_i[304];
  assign N1786 = N1785 & N1788;
  assign N1789 = sel_i[307] & sel_i[306];
  assign N1791 = N1790 & N1793;
  assign N1794 = sel_i[309] & sel_i[308];
  assign N1796 = N1795 & N1798;
  assign N1799 = sel_i[311] & sel_i[310];
  assign N1801 = N1800 & N1803;
  assign N1804 = sel_i[313] & sel_i[312];
  assign N1806 = N1805 & N1808;
  assign N1809 = sel_i[315] & sel_i[314];
  assign N1811 = N1810 & N1813;
  assign N1814 = sel_i[317] & sel_i[316];
  assign N1816 = N1815 & N1818;
  assign N1819 = sel_i[319] & sel_i[318];
  assign N1821 = N1820 & N1823;
  assign N1824 = sel_i[321] & sel_i[320];
  assign N1826 = N1825 & N1828;
  assign N1829 = sel_i[323] & sel_i[322];
  assign N1831 = N1830 & N1833;
  assign N1834 = sel_i[325] & sel_i[324];
  assign N1836 = N1835 & N1838;
  assign N1839 = sel_i[327] & sel_i[326];
  assign N1841 = N1840 & N1843;
  assign N1844 = sel_i[329] & sel_i[328];
  assign N1846 = N1845 & N1848;
  assign N1849 = sel_i[331] & sel_i[330];
  assign N1851 = N1850 & N1853;
  assign N1854 = sel_i[333] & sel_i[332];
  assign N1856 = N1855 & N1858;
  assign N1859 = sel_i[335] & sel_i[334];
  assign N1861 = N1860 & N1863;
  assign N1864 = sel_i[337] & sel_i[336];
  assign N1866 = N1865 & N1868;
  assign N1869 = sel_i[339] & sel_i[338];
  assign N1871 = N1870 & N1873;
  assign N1874 = sel_i[341] & sel_i[340];
  assign N1876 = N1875 & N1878;
  assign N1879 = sel_i[343] & sel_i[342];
  assign N1881 = N1880 & N1883;
  assign N1884 = sel_i[345] & sel_i[344];
  assign N1886 = N1885 & N1888;
  assign N1889 = sel_i[347] & sel_i[346];
  assign N1891 = N1890 & N1893;
  assign N1894 = sel_i[349] & sel_i[348];
  assign N1896 = N1895 & N1898;
  assign N1899 = sel_i[351] & sel_i[350];
  assign N1901 = N1900 & N1903;
  assign N1904 = sel_i[353] & sel_i[352];
  assign N1906 = N1905 & N1908;
  assign N1909 = sel_i[355] & sel_i[354];
  assign N1911 = N1910 & N1913;
  assign N1914 = sel_i[357] & sel_i[356];
  assign N1916 = N1915 & N1918;
  assign N1919 = sel_i[359] & sel_i[358];
  assign N1921 = N1920 & N1923;
  assign N1924 = sel_i[361] & sel_i[360];
  assign N1926 = N1925 & N1928;
  assign N1929 = sel_i[363] & sel_i[362];
  assign N1931 = N1930 & N1933;
  assign N1934 = sel_i[365] & sel_i[364];
  assign N1936 = N1935 & N1938;
  assign N1939 = sel_i[367] & sel_i[366];
  assign N1941 = N1940 & N1943;
  assign N1944 = sel_i[369] & sel_i[368];
  assign N1946 = N1945 & N1948;
  assign N1949 = sel_i[371] & sel_i[370];
  assign N1951 = N1950 & N1953;
  assign N1954 = sel_i[373] & sel_i[372];
  assign N1956 = N1955 & N1958;
  assign N1959 = sel_i[375] & sel_i[374];
  assign N1961 = N1960 & N1963;
  assign N1964 = sel_i[377] & sel_i[376];
  assign N1966 = N1965 & N1968;
  assign N1969 = sel_i[379] & sel_i[378];
  assign N1971 = N1970 & N1973;
  assign N1974 = sel_i[381] & sel_i[380];
  assign N1976 = N1975 & N1978;
  assign N1979 = sel_i[383] & sel_i[382];
  assign N1981 = N1980 & N1983;
  assign N1984 = sel_i[385] & sel_i[384];
  assign N1986 = N1985 & N1988;
  assign N1989 = sel_i[387] & sel_i[386];
  assign N1991 = N1990 & N1993;
  assign N1994 = sel_i[389] & sel_i[388];
  assign N1996 = N1995 & N1998;
  assign N1999 = sel_i[391] & sel_i[390];
  assign N2001 = N2000 & N2003;
  assign N2004 = sel_i[393] & sel_i[392];
  assign N2006 = N2005 & N2008;
  assign N2009 = sel_i[395] & sel_i[394];
  assign N2011 = N2010 & N2013;
  assign N2014 = sel_i[397] & sel_i[396];
  assign N2016 = N2015 & N2018;
  assign N2019 = sel_i[399] & sel_i[398];
  assign N2021 = N2020 & N2023;
  assign N2024 = sel_i[401] & sel_i[400];
  assign N2026 = N2025 & N2028;
  assign N2029 = sel_i[403] & sel_i[402];
  assign N2031 = N2030 & N2033;
  assign N2034 = sel_i[405] & sel_i[404];
  assign N2036 = N2035 & N2038;
  assign N2039 = sel_i[407] & sel_i[406];
  assign N2041 = N2040 & N2043;
  assign N2044 = sel_i[409] & sel_i[408];
  assign N2046 = N2045 & N2048;
  assign N2049 = sel_i[411] & sel_i[410];
  assign N2051 = N2050 & N2053;
  assign N2054 = sel_i[413] & sel_i[412];
  assign N2056 = N2055 & N2058;
  assign N2059 = sel_i[415] & sel_i[414];
  assign N2061 = N2060 & N2063;
  assign N2064 = sel_i[417] & sel_i[416];
  assign N2066 = N2065 & N2068;
  assign N2069 = sel_i[419] & sel_i[418];
  assign N2071 = N2070 & N2073;
  assign N2074 = sel_i[421] & sel_i[420];
  assign N2076 = N2075 & N2078;
  assign N2079 = sel_i[423] & sel_i[422];
  assign N2081 = N2080 & N2083;
  assign N2084 = sel_i[425] & sel_i[424];
  assign N2086 = N2085 & N2088;
  assign N2089 = sel_i[427] & sel_i[426];
  assign N2091 = N2090 & N2093;
  assign N2094 = sel_i[429] & sel_i[428];
  assign N2096 = N2095 & N2098;
  assign N2099 = sel_i[431] & sel_i[430];
  assign N2101 = N2100 & N2103;
  assign N2104 = sel_i[433] & sel_i[432];
  assign N2106 = N2105 & N2108;
  assign N2109 = sel_i[435] & sel_i[434];
  assign N2111 = N2110 & N2113;
  assign N2114 = sel_i[437] & sel_i[436];
  assign N2116 = N2115 & N2118;
  assign N2119 = sel_i[439] & sel_i[438];
  assign N2121 = N2120 & N2123;
  assign N2124 = sel_i[441] & sel_i[440];
  assign N2126 = N2125 & N2128;
  assign N2129 = sel_i[443] & sel_i[442];
  assign N2131 = N2130 & N2133;
  assign N2134 = sel_i[445] & sel_i[444];
  assign N2136 = N2135 & N2138;
  assign N2139 = sel_i[447] & sel_i[446];
  assign N2141 = N2140 & N2143;
  assign N2144 = sel_i[449] & sel_i[448];
  assign N2146 = N2145 & N2148;
  assign N2149 = sel_i[451] & sel_i[450];
  assign N2151 = N2150 & N2153;
  assign N2154 = sel_i[453] & sel_i[452];
  assign N2156 = N2155 & N2158;
  assign N2159 = sel_i[455] & sel_i[454];
  assign N2161 = N2160 & N2163;
  assign N2164 = sel_i[457] & sel_i[456];
  assign N2166 = N2165 & N2168;
  assign N2169 = sel_i[459] & sel_i[458];
  assign N2171 = N2170 & N2173;
  assign N2174 = sel_i[461] & sel_i[460];
  assign N2176 = N2175 & N2178;
  assign N2179 = sel_i[463] & sel_i[462];
  assign N2181 = N2180 & N2183;
  assign N2184 = sel_i[465] & sel_i[464];
  assign N2186 = N2185 & N2188;
  assign N2189 = sel_i[467] & sel_i[466];
  assign N2191 = N2190 & N2193;
  assign N2194 = sel_i[469] & sel_i[468];
  assign N2196 = N2195 & N2198;
  assign N2199 = sel_i[471] & sel_i[470];
  assign N2201 = N2200 & N2203;
  assign N2204 = sel_i[473] & sel_i[472];
  assign N2206 = N2205 & N2208;
  assign N2209 = sel_i[475] & sel_i[474];
  assign N2211 = N2210 & N2213;
  assign N2214 = sel_i[477] & sel_i[476];
  assign N2216 = N2215 & N2218;
  assign N2219 = sel_i[479] & sel_i[478];
  assign N2221 = N2220 & N2223;
  assign N2224 = sel_i[481] & sel_i[480];
  assign N2226 = N2225 & N2228;
  assign N2229 = sel_i[483] & sel_i[482];
  assign N2231 = N2230 & N2233;
  assign N2234 = sel_i[485] & sel_i[484];
  assign N2236 = N2235 & N2238;
  assign N2239 = sel_i[487] & sel_i[486];
  assign N2241 = N2240 & N2243;
  assign N2244 = sel_i[489] & sel_i[488];
  assign N2246 = N2245 & N2248;
  assign N2249 = sel_i[491] & sel_i[490];
  assign N2251 = N2250 & N2253;
  assign N2254 = sel_i[493] & sel_i[492];
  assign N2256 = N2255 & N2258;
  assign N2259 = sel_i[495] & sel_i[494];
  assign N2261 = N2260 & N2263;
  assign N2264 = sel_i[497] & sel_i[496];
  assign N2266 = N2265 & N2268;
  assign N2269 = sel_i[499] & sel_i[498];
  assign N2271 = N2270 & N2273;
  assign N2274 = sel_i[501] & sel_i[500];
  assign N2276 = N2275 & N2278;
  assign N2279 = sel_i[503] & sel_i[502];
  assign N2281 = N2280 & N2283;
  assign N2284 = sel_i[505] & sel_i[504];
  assign N2286 = N2285 & N2288;
  assign N2289 = sel_i[507] & sel_i[506];
  assign N2291 = N2290 & N2293;
  assign N2294 = sel_i[509] & sel_i[508];
  assign N2296 = N2295 & N2298;
  assign N2299 = sel_i[511] & sel_i[510];
  assign N2301 = N2300 & N2303;
  assign N2304 = sel_i[513] & sel_i[512];
  assign N2306 = N2305 & N2308;
  assign N2309 = sel_i[515] & sel_i[514];
  assign N2311 = N2310 & N2313;
  assign N2314 = sel_i[517] & sel_i[516];
  assign N2316 = N2315 & N2318;
  assign N2319 = sel_i[519] & sel_i[518];
  assign N2321 = N2320 & N2323;
  assign N2324 = sel_i[521] & sel_i[520];
  assign N2326 = N2325 & N2328;
  assign N2329 = sel_i[523] & sel_i[522];
  assign N2331 = N2330 & N2333;
  assign N2334 = sel_i[525] & sel_i[524];
  assign N2336 = N2335 & N2338;
  assign N2339 = sel_i[527] & sel_i[526];
  assign N2341 = N2340 & N2343;
  assign N2344 = sel_i[529] & sel_i[528];
  assign N2346 = N2345 & N2348;
  assign N2349 = sel_i[531] & sel_i[530];
  assign N2351 = N2350 & N2353;
  assign N2354 = sel_i[533] & sel_i[532];
  assign N2356 = N2355 & N2358;
  assign N2359 = sel_i[535] & sel_i[534];
  assign N2361 = N2360 & N2363;
  assign N2364 = sel_i[537] & sel_i[536];
  assign N2366 = N2365 & N2368;
  assign N2369 = sel_i[539] & sel_i[538];
  assign N2371 = N2370 & N2373;
  assign N2374 = sel_i[541] & sel_i[540];
  assign N2376 = N2375 & N2378;
  assign N2379 = sel_i[543] & sel_i[542];
  assign N2381 = N2380 & N2383;
  assign N2384 = sel_i[545] & sel_i[544];
  assign N2386 = N2385 & N2388;
  assign N2389 = sel_i[547] & sel_i[546];
  assign N2391 = N2390 & N2393;
  assign N2394 = sel_i[549] & sel_i[548];
  assign N2396 = N2395 & N2398;
  assign N2399 = sel_i[551] & sel_i[550];
  assign N2401 = N2400 & N2403;
  assign N2404 = sel_i[553] & sel_i[552];
  assign N2406 = N2405 & N2408;
  assign N2409 = sel_i[555] & sel_i[554];
  assign N2411 = N2410 & N2413;
  assign N2414 = sel_i[557] & sel_i[556];
  assign N2416 = N2415 & N2418;
  assign N2419 = sel_i[559] & sel_i[558];
  assign N2421 = N2420 & N2423;
  assign N2424 = sel_i[561] & sel_i[560];
  assign N2426 = N2425 & N2428;
  assign N2429 = sel_i[563] & sel_i[562];
  assign N2431 = N2430 & N2433;
  assign N2434 = sel_i[565] & sel_i[564];
  assign N2436 = N2435 & N2438;
  assign N2439 = sel_i[567] & sel_i[566];
  assign N2441 = N2440 & N2443;
  assign N2444 = sel_i[569] & sel_i[568];
  assign N2446 = N2445 & N2448;
  assign N2449 = sel_i[571] & sel_i[570];
  assign N2451 = N2450 & N2453;
  assign N2454 = sel_i[573] & sel_i[572];
  assign N2456 = N2455 & N2458;
  assign N2459 = sel_i[575] & sel_i[574];
  assign N2461 = N2460 & N2463;
  assign N2464 = sel_i[577] & sel_i[576];
  assign N2466 = N2465 & N2468;
  assign N2469 = sel_i[579] & sel_i[578];
  assign N2471 = N2470 & N2473;
  assign N2474 = sel_i[581] & sel_i[580];
  assign N2476 = N2475 & N2478;
  assign N2479 = sel_i[583] & sel_i[582];
  assign N2481 = N2480 & N2483;
  assign N2484 = sel_i[585] & sel_i[584];
  assign N2486 = N2485 & N2488;
  assign N2489 = sel_i[587] & sel_i[586];
  assign N2491 = N2490 & N2493;
  assign N2494 = sel_i[589] & sel_i[588];
  assign N2496 = N2495 & N2498;
  assign N2499 = sel_i[591] & sel_i[590];
  assign N2501 = N2500 & N2503;
  assign N2504 = sel_i[593] & sel_i[592];
  assign N2506 = N2505 & N2508;
  assign N2509 = sel_i[595] & sel_i[594];
  assign N2511 = N2510 & N2513;
  assign N2514 = sel_i[597] & sel_i[596];
  assign N2516 = N2515 & N2518;
  assign N2519 = sel_i[599] & sel_i[598];
  assign N2521 = N2520 & N2523;
  assign N2524 = sel_i[601] & sel_i[600];
  assign N2526 = N2525 & N2528;
  assign N2529 = sel_i[603] & sel_i[602];
  assign N2531 = N2530 & N2533;
  assign N2534 = sel_i[605] & sel_i[604];
  assign N2536 = N2535 & N2538;
  assign N2539 = sel_i[607] & sel_i[606];
  assign N2541 = N2540 & N2543;
  assign N2544 = sel_i[609] & sel_i[608];
  assign N2546 = N2545 & N2548;
  assign N2549 = sel_i[611] & sel_i[610];
  assign N2551 = N2550 & N2553;
  assign N2554 = sel_i[613] & sel_i[612];
  assign N2556 = N2555 & N2558;
  assign N2559 = sel_i[615] & sel_i[614];
  assign N2561 = N2560 & N2563;
  assign N2564 = sel_i[617] & sel_i[616];
  assign N2566 = N2565 & N2568;
  assign N2569 = sel_i[619] & sel_i[618];
  assign N2571 = N2570 & N2573;
  assign N2574 = sel_i[621] & sel_i[620];
  assign N2576 = N2575 & N2578;
  assign N2579 = sel_i[623] & sel_i[622];
  assign N2581 = N2580 & N2583;
  assign N2584 = sel_i[625] & sel_i[624];
  assign N2586 = N2585 & N2588;
  assign N2589 = sel_i[627] & sel_i[626];
  assign N2591 = N2590 & N2593;
  assign N2594 = sel_i[629] & sel_i[628];
  assign N2596 = N2595 & N2598;
  assign N2599 = sel_i[631] & sel_i[630];
  assign N2601 = N2600 & N2603;
  assign N2604 = sel_i[633] & sel_i[632];
  assign N2606 = N2605 & N2608;
  assign N2609 = sel_i[635] & sel_i[634];
  assign N2611 = N2610 & N2613;
  assign N2614 = sel_i[637] & sel_i[636];
  assign N2616 = N2615 & N2618;
  assign N2619 = sel_i[639] & sel_i[638];
  assign N2621 = N2620 & N2623;
  assign N2624 = sel_i[641] & sel_i[640];
  assign N2626 = N2625 & N2628;
  assign N2629 = sel_i[643] & sel_i[642];
  assign N2631 = N2630 & N2633;
  assign N2634 = sel_i[645] & sel_i[644];
  assign N2636 = N2635 & N2638;
  assign N2639 = sel_i[647] & sel_i[646];
  assign N2641 = N2640 & N2643;
  assign N2644 = sel_i[649] & sel_i[648];
  assign N2646 = N2645 & N2648;
  assign N2649 = sel_i[651] & sel_i[650];
  assign N2651 = N2650 & N2653;
  assign N2654 = sel_i[653] & sel_i[652];
  assign N2656 = N2655 & N2658;
  assign N2659 = sel_i[655] & sel_i[654];
  assign N2661 = N2660 & N2663;
  assign N2664 = sel_i[657] & sel_i[656];
  assign N2666 = N2665 & N2668;
  assign N2669 = sel_i[659] & sel_i[658];
  assign N2671 = N2670 & N2673;
  assign N2674 = sel_i[661] & sel_i[660];
  assign N2676 = N2675 & N2678;
  assign N2679 = sel_i[663] & sel_i[662];
  assign N2681 = N2680 & N2683;
  assign N2684 = sel_i[665] & sel_i[664];
  assign N2686 = N2685 & N2688;
  assign N2689 = sel_i[667] & sel_i[666];
  assign N2691 = N2690 & N2693;
  assign N2694 = sel_i[669] & sel_i[668];
  assign N2696 = N2695 & N2698;
  assign N2699 = sel_i[671] & sel_i[670];
  assign N2701 = N2700 & N2703;
  assign N2704 = sel_i[673] & sel_i[672];
  assign N2706 = N2705 & N2708;
  assign N2709 = sel_i[675] & sel_i[674];
  assign N2711 = N2710 & N2713;
  assign N2714 = sel_i[677] & sel_i[676];
  assign N2716 = N2715 & N2718;
  assign N2719 = sel_i[679] & sel_i[678];
  assign N2721 = N2720 & N2723;
  assign N2724 = sel_i[681] & sel_i[680];
  assign N2726 = N2725 & N2728;
  assign N2729 = sel_i[683] & sel_i[682];
  assign N2731 = N2730 & N2733;
  assign N2734 = sel_i[685] & sel_i[684];
  assign N2736 = N2735 & N2738;
  assign N2739 = sel_i[687] & sel_i[686];
  assign N2741 = N2740 & N2743;
  assign N2744 = sel_i[689] & sel_i[688];
  assign N2746 = N2745 & N2748;
  assign N2749 = sel_i[691] & sel_i[690];
  assign N2751 = N2750 & N2753;
  assign N2754 = sel_i[693] & sel_i[692];
  assign N2756 = N2755 & N2758;
  assign N2759 = sel_i[695] & sel_i[694];
  assign N2761 = N2760 & N2763;
  assign N2764 = sel_i[697] & sel_i[696];
  assign N2766 = N2765 & N2768;
  assign N2769 = sel_i[699] & sel_i[698];
  assign N2771 = N2770 & N2773;
  assign N2774 = sel_i[701] & sel_i[700];
  assign N2776 = N2775 & N2778;
  assign N2779 = sel_i[703] & sel_i[702];
  assign N2781 = N2780 & N2783;
  assign N2784 = sel_i[705] & sel_i[704];
  assign N2786 = N2785 & N2788;
  assign N2789 = sel_i[707] & sel_i[706];
  assign N2791 = N2790 & N2793;
  assign N2794 = sel_i[709] & sel_i[708];
  assign N2796 = N2795 & N2798;
  assign N2799 = sel_i[711] & sel_i[710];
  assign N2801 = N2800 & N2803;
  assign N2804 = sel_i[713] & sel_i[712];
  assign N2806 = N2805 & N2808;
  assign N2809 = sel_i[715] & sel_i[714];
  assign N2811 = N2810 & N2813;
  assign N2814 = sel_i[717] & sel_i[716];
  assign N2816 = N2815 & N2818;
  assign N2819 = sel_i[719] & sel_i[718];
  assign N2821 = N2820 & N2823;
  assign N2824 = sel_i[721] & sel_i[720];
  assign N2826 = N2825 & N2828;
  assign N2829 = sel_i[723] & sel_i[722];
  assign N2831 = N2830 & N2833;
  assign N2834 = sel_i[725] & sel_i[724];
  assign N2836 = N2835 & N2838;
  assign N2839 = sel_i[727] & sel_i[726];
  assign N2841 = N2840 & N2843;
  assign N2844 = sel_i[729] & sel_i[728];
  assign N2846 = N2845 & N2848;
  assign N2849 = sel_i[731] & sel_i[730];
  assign N2851 = N2850 & N2853;
  assign N2854 = sel_i[733] & sel_i[732];
  assign N2856 = N2855 & N2858;
  assign N2859 = sel_i[735] & sel_i[734];
  assign N2861 = N2860 & N2863;
  assign N2864 = sel_i[737] & sel_i[736];
  assign N2866 = N2865 & N2868;
  assign N2869 = sel_i[739] & sel_i[738];
  assign N2871 = N2870 & N2873;
  assign N2874 = sel_i[741] & sel_i[740];
  assign N2876 = N2875 & N2878;
  assign N2879 = sel_i[743] & sel_i[742];
  assign N2881 = N2880 & N2883;
  assign N2884 = sel_i[745] & sel_i[744];
  assign N2886 = N2885 & N2888;
  assign N2889 = sel_i[747] & sel_i[746];
  assign N2891 = N2890 & N2893;
  assign N2894 = sel_i[749] & sel_i[748];
  assign N2896 = N2895 & N2898;
  assign N2899 = sel_i[751] & sel_i[750];
  assign N2901 = N2900 & N2903;
  assign N2904 = sel_i[753] & sel_i[752];
  assign N2906 = N2905 & N2908;
  assign N2909 = sel_i[755] & sel_i[754];
  assign N2911 = N2910 & N2913;
  assign N2914 = sel_i[757] & sel_i[756];
  assign N2916 = N2915 & N2918;
  assign N2919 = sel_i[759] & sel_i[758];
  assign N2921 = N2920 & N2923;
  assign N2924 = sel_i[761] & sel_i[760];
  assign N2926 = N2925 & N2928;
  assign N2929 = sel_i[763] & sel_i[762];
  assign N2931 = N2930 & N2933;
  assign N2934 = sel_i[765] & sel_i[764];
  assign N2936 = N2935 & N2938;
  assign N2939 = sel_i[767] & sel_i[766];
  assign N2941 = N2940 & N2943;
  assign N2944 = sel_i[769] & sel_i[768];
  assign N2946 = N2945 & N2948;
  assign N2949 = sel_i[771] & sel_i[770];
  assign N2951 = N2950 & N2953;
  assign N2954 = sel_i[773] & sel_i[772];
  assign N2956 = N2955 & N2958;
  assign N2959 = sel_i[775] & sel_i[774];
  assign N2961 = N2960 & N2963;
  assign N2964 = sel_i[777] & sel_i[776];
  assign N2966 = N2965 & N2968;
  assign N2969 = sel_i[779] & sel_i[778];
  assign N2971 = N2970 & N2973;
  assign N2974 = sel_i[781] & sel_i[780];
  assign N2976 = N2975 & N2978;
  assign N2979 = sel_i[783] & sel_i[782];
  assign N2981 = N2980 & N2983;
  assign N2984 = sel_i[785] & sel_i[784];
  assign N2986 = N2985 & N2988;
  assign N2989 = sel_i[787] & sel_i[786];
  assign N2991 = N2990 & N2993;
  assign N2994 = sel_i[789] & sel_i[788];
  assign N2996 = N2995 & N2998;
  assign N2999 = sel_i[791] & sel_i[790];
  assign N3001 = N3000 & N3003;
  assign N3004 = sel_i[793] & sel_i[792];
  assign N3006 = N3005 & N3008;
  assign N3009 = sel_i[795] & sel_i[794];
  assign N3011 = N3010 & N3013;
  assign N3014 = sel_i[797] & sel_i[796];
  assign N3016 = N3015 & N3018;
  assign N3019 = sel_i[799] & sel_i[798];
  assign N3021 = N3020 & N3023;
  assign N3024 = sel_i[801] & sel_i[800];
  assign N3026 = N3025 & N3028;
  assign N3029 = sel_i[803] & sel_i[802];
  assign N3031 = N3030 & N3033;
  assign N3034 = sel_i[805] & sel_i[804];
  assign N3036 = N3035 & N3038;
  assign N3039 = sel_i[807] & sel_i[806];
  assign N3041 = N3040 & N3043;
  assign N3044 = sel_i[809] & sel_i[808];
  assign N3046 = N3045 & N3048;
  assign N3049 = sel_i[811] & sel_i[810];
  assign N3051 = N3050 & N3053;
  assign N3054 = sel_i[813] & sel_i[812];
  assign N3056 = N3055 & N3058;
  assign N3059 = sel_i[815] & sel_i[814];
  assign N3061 = N3060 & N3063;
  assign N3064 = sel_i[817] & sel_i[816];
  assign N3066 = N3065 & N3068;
  assign N3069 = sel_i[819] & sel_i[818];
  assign N3071 = N3070 & N3073;
  assign N3074 = sel_i[821] & sel_i[820];
  assign N3076 = N3075 & N3078;
  assign N3079 = sel_i[823] & sel_i[822];
  assign N3081 = N3080 & N3083;
  assign N3084 = sel_i[825] & sel_i[824];
  assign N3086 = N3085 & N3088;
  assign N3089 = sel_i[827] & sel_i[826];
  assign N3091 = N3090 & N3093;
  assign N3094 = sel_i[829] & sel_i[828];
  assign N3096 = N3095 & N3098;
  assign N3099 = sel_i[831] & sel_i[830];
  assign N3101 = N3100 & N3103;
  assign N3104 = sel_i[833] & sel_i[832];
  assign N3106 = N3105 & N3108;
  assign N3109 = sel_i[835] & sel_i[834];
  assign N3111 = N3110 & N3113;
  assign N3114 = sel_i[837] & sel_i[836];
  assign N3116 = N3115 & N3118;
  assign N3119 = sel_i[839] & sel_i[838];
  assign N3121 = N3120 & N3123;
  assign N3124 = sel_i[841] & sel_i[840];
  assign N3126 = N3125 & N3128;
  assign N3129 = sel_i[843] & sel_i[842];
  assign N3131 = N3130 & N3133;
  assign N3134 = sel_i[845] & sel_i[844];
  assign N3136 = N3135 & N3138;
  assign N3139 = sel_i[847] & sel_i[846];
  assign N3141 = N3140 & N3143;
  assign N3144 = sel_i[849] & sel_i[848];
  assign N3146 = N3145 & N3148;
  assign N3149 = sel_i[851] & sel_i[850];
  assign N3151 = N3150 & N3153;
  assign N3154 = sel_i[853] & sel_i[852];
  assign N3156 = N3155 & N3158;
  assign N3159 = sel_i[855] & sel_i[854];
  assign N3161 = N3160 & N3163;
  assign N3164 = sel_i[857] & sel_i[856];
  assign N3166 = N3165 & N3168;
  assign N3169 = sel_i[859] & sel_i[858];
  assign N3171 = N3170 & N3173;
  assign N3174 = sel_i[861] & sel_i[860];
  assign N3176 = N3175 & N3178;
  assign N3179 = sel_i[863] & sel_i[862];
  assign N3181 = N3180 & N3183;
  assign N3184 = sel_i[865] & sel_i[864];
  assign N3186 = N3185 & N3188;
  assign N3189 = sel_i[867] & sel_i[866];
  assign N3191 = N3190 & N3193;
  assign N3194 = sel_i[869] & sel_i[868];
  assign N3196 = N3195 & N3198;
  assign N3199 = sel_i[871] & sel_i[870];
  assign N3201 = N3200 & N3203;
  assign N3204 = sel_i[873] & sel_i[872];
  assign N3206 = N3205 & N3208;
  assign N3209 = sel_i[875] & sel_i[874];
  assign N3211 = N3210 & N3213;
  assign N3214 = sel_i[877] & sel_i[876];
  assign N3216 = N3215 & N3218;
  assign N3219 = sel_i[879] & sel_i[878];
  assign N3221 = N3220 & N3223;
  assign N3224 = sel_i[881] & sel_i[880];
  assign N3226 = N3225 & N3228;
  assign N3229 = sel_i[883] & sel_i[882];
  assign N3231 = N3230 & N3233;
  assign N3234 = sel_i[885] & sel_i[884];
  assign N3236 = N3235 & N3238;
  assign N3239 = sel_i[887] & sel_i[886];
  assign N3241 = N3240 & N3243;
  assign N3244 = sel_i[889] & sel_i[888];
  assign N3246 = N3245 & N3248;
  assign N3249 = sel_i[891] & sel_i[890];
  assign N3251 = N3250 & N3253;
  assign N3254 = sel_i[893] & sel_i[892];
  assign N3256 = N3255 & N3258;
  assign N3259 = sel_i[895] & sel_i[894];
  assign N3261 = N3260 & N3263;
  assign N3264 = sel_i[897] & sel_i[896];
  assign N3266 = N3265 & N3268;
  assign N3269 = sel_i[899] & sel_i[898];
  assign N3271 = N3270 & N3273;
  assign N3274 = sel_i[901] & sel_i[900];
  assign N3276 = N3275 & N3278;
  assign N3279 = sel_i[903] & sel_i[902];
  assign N3281 = N3280 & N3283;
  assign N3284 = sel_i[905] & sel_i[904];
  assign N3286 = N3285 & N3288;
  assign N3289 = sel_i[907] & sel_i[906];
  assign N3291 = N3290 & N3293;
  assign N3294 = sel_i[909] & sel_i[908];
  assign N3296 = N3295 & N3298;
  assign N3299 = sel_i[911] & sel_i[910];
  assign N3301 = N3300 & N3303;
  assign N3304 = sel_i[913] & sel_i[912];
  assign N3306 = N3305 & N3308;
  assign N3309 = sel_i[915] & sel_i[914];
  assign N3311 = N3310 & N3313;
  assign N3314 = sel_i[917] & sel_i[916];
  assign N3316 = N3315 & N3318;
  assign N3319 = sel_i[919] & sel_i[918];
  assign N3321 = N3320 & N3323;
  assign N3324 = sel_i[921] & sel_i[920];
  assign N3326 = N3325 & N3328;
  assign N3329 = sel_i[923] & sel_i[922];
  assign N3331 = N3330 & N3333;
  assign N3334 = sel_i[925] & sel_i[924];
  assign N3336 = N3335 & N3338;
  assign N3339 = sel_i[927] & sel_i[926];
  assign N3341 = N3340 & N3343;
  assign N3344 = sel_i[929] & sel_i[928];
  assign N3346 = N3345 & N3348;
  assign N3349 = sel_i[931] & sel_i[930];
  assign N3351 = N3350 & N3353;
  assign N3354 = sel_i[933] & sel_i[932];
  assign N3356 = N3355 & N3358;
  assign N3359 = sel_i[935] & sel_i[934];
  assign N3361 = N3360 & N3363;
  assign N3364 = sel_i[937] & sel_i[936];
  assign N3366 = N3365 & N3368;
  assign N3369 = sel_i[939] & sel_i[938];
  assign N3371 = N3370 & N3373;
  assign N3374 = sel_i[941] & sel_i[940];
  assign N3376 = N3375 & N3378;
  assign N3379 = sel_i[943] & sel_i[942];
  assign N3381 = N3380 & N3383;
  assign N3384 = sel_i[945] & sel_i[944];
  assign N3386 = N3385 & N3388;
  assign N3389 = sel_i[947] & sel_i[946];
  assign N3391 = N3390 & N3393;
  assign N3394 = sel_i[949] & sel_i[948];
  assign N3396 = N3395 & N3398;
  assign N3399 = sel_i[951] & sel_i[950];
  assign N3401 = N3400 & N3403;
  assign N3404 = sel_i[953] & sel_i[952];
  assign N3406 = N3405 & N3408;
  assign N3409 = sel_i[955] & sel_i[954];
  assign N3411 = N3410 & N3413;
  assign N3414 = sel_i[957] & sel_i[956];
  assign N3416 = N3415 & N3418;
  assign N3419 = sel_i[959] & sel_i[958];
  assign N3421 = N3420 & N3423;
  assign N3424 = sel_i[961] & sel_i[960];
  assign N3426 = N3425 & N3428;
  assign N3429 = sel_i[963] & sel_i[962];
  assign N3431 = N3430 & N3433;
  assign N3434 = sel_i[965] & sel_i[964];
  assign N3436 = N3435 & N3438;
  assign N3439 = sel_i[967] & sel_i[966];
  assign N3441 = N3440 & N3443;
  assign N3444 = sel_i[969] & sel_i[968];
  assign N3446 = N3445 & N3448;
  assign N3449 = sel_i[971] & sel_i[970];
  assign N3451 = N3450 & N3453;
  assign N3454 = sel_i[973] & sel_i[972];
  assign N3456 = N3455 & N3458;
  assign N3459 = sel_i[975] & sel_i[974];
  assign N3461 = N3460 & N3463;
  assign N3464 = sel_i[977] & sel_i[976];
  assign N3466 = N3465 & N3468;
  assign N3469 = sel_i[979] & sel_i[978];
  assign N3471 = N3470 & N3473;
  assign N3474 = sel_i[981] & sel_i[980];
  assign N3476 = N3475 & N3478;
  assign N3479 = sel_i[983] & sel_i[982];
  assign N3481 = N3480 & N3483;
  assign N3484 = sel_i[985] & sel_i[984];
  assign N3486 = N3485 & N3488;
  assign N3489 = sel_i[987] & sel_i[986];
  assign N3491 = N3490 & N3493;
  assign N3494 = sel_i[989] & sel_i[988];
  assign N3496 = N3495 & N3498;
  assign N3499 = sel_i[991] & sel_i[990];
  assign N3501 = N3500 & N3503;
  assign N3504 = sel_i[993] & sel_i[992];
  assign N3506 = N3505 & N3508;
  assign N3509 = sel_i[995] & sel_i[994];
  assign N3511 = N3510 & N3513;
  assign N3514 = sel_i[997] & sel_i[996];
  assign N3516 = N3515 & N3518;
  assign N3519 = sel_i[999] & sel_i[998];
  assign N3521 = N3520 & N3523;
  assign N3524 = sel_i[1001] & sel_i[1000];
  assign N3526 = N3525 & N3528;
  assign N3529 = sel_i[1003] & sel_i[1002];
  assign N3531 = N3530 & N3533;
  assign N3534 = sel_i[1005] & sel_i[1004];
  assign N3536 = N3535 & N3538;
  assign N3539 = sel_i[1007] & sel_i[1006];
  assign N3541 = N3540 & N3543;
  assign N3544 = sel_i[1009] & sel_i[1008];
  assign N3546 = N3545 & N3548;
  assign N3549 = sel_i[1011] & sel_i[1010];
  assign N3551 = N3550 & N3553;
  assign N3554 = sel_i[1013] & sel_i[1012];
  assign N3556 = N3555 & N3558;
  assign N3559 = sel_i[1015] & sel_i[1014];
  assign N3561 = N3560 & N3563;
  assign N3564 = sel_i[1017] & sel_i[1016];
  assign N3566 = N3565 & N3568;
  assign N3569 = sel_i[1019] & sel_i[1018];
  assign N3571 = N3570 & N3573;
  assign N3574 = sel_i[1021] & sel_i[1020];
  assign N3576 = N3575 & N3578;
  assign N3579 = sel_i[1023] & sel_i[1022];
  assign N3581 = N3580 & N3583;
  assign N1028 = ~sel_i[0];
  assign N1033 = ~sel_i[2];
  assign N1038 = ~sel_i[4];
  assign N1043 = ~sel_i[6];
  assign N1048 = ~sel_i[8];
  assign N1053 = ~sel_i[10];
  assign N1058 = ~sel_i[12];
  assign N1063 = ~sel_i[14];
  assign N1068 = ~sel_i[16];
  assign N1073 = ~sel_i[18];
  assign N1078 = ~sel_i[20];
  assign N1083 = ~sel_i[22];
  assign N1088 = ~sel_i[24];
  assign N1093 = ~sel_i[26];
  assign N1098 = ~sel_i[28];
  assign N1103 = ~sel_i[30];
  assign N1108 = ~sel_i[32];
  assign N1113 = ~sel_i[34];
  assign N1118 = ~sel_i[36];
  assign N1123 = ~sel_i[38];
  assign N1128 = ~sel_i[40];
  assign N1133 = ~sel_i[42];
  assign N1138 = ~sel_i[44];
  assign N1143 = ~sel_i[46];
  assign N1148 = ~sel_i[48];
  assign N1153 = ~sel_i[50];
  assign N1158 = ~sel_i[52];
  assign N1163 = ~sel_i[54];
  assign N1168 = ~sel_i[56];
  assign N1173 = ~sel_i[58];
  assign N1178 = ~sel_i[60];
  assign N1183 = ~sel_i[62];
  assign N1188 = ~sel_i[64];
  assign N1193 = ~sel_i[66];
  assign N1198 = ~sel_i[68];
  assign N1203 = ~sel_i[70];
  assign N1208 = ~sel_i[72];
  assign N1213 = ~sel_i[74];
  assign N1218 = ~sel_i[76];
  assign N1223 = ~sel_i[78];
  assign N1228 = ~sel_i[80];
  assign N1233 = ~sel_i[82];
  assign N1238 = ~sel_i[84];
  assign N1243 = ~sel_i[86];
  assign N1248 = ~sel_i[88];
  assign N1253 = ~sel_i[90];
  assign N1258 = ~sel_i[92];
  assign N1263 = ~sel_i[94];
  assign N1268 = ~sel_i[96];
  assign N1273 = ~sel_i[98];
  assign N1278 = ~sel_i[100];
  assign N1283 = ~sel_i[102];
  assign N1288 = ~sel_i[104];
  assign N1293 = ~sel_i[106];
  assign N1298 = ~sel_i[108];
  assign N1303 = ~sel_i[110];
  assign N1308 = ~sel_i[112];
  assign N1313 = ~sel_i[114];
  assign N1318 = ~sel_i[116];
  assign N1323 = ~sel_i[118];
  assign N1328 = ~sel_i[120];
  assign N1333 = ~sel_i[122];
  assign N1338 = ~sel_i[124];
  assign N1343 = ~sel_i[126];
  assign N1348 = ~sel_i[128];
  assign N1353 = ~sel_i[130];
  assign N1358 = ~sel_i[132];
  assign N1363 = ~sel_i[134];
  assign N1368 = ~sel_i[136];
  assign N1373 = ~sel_i[138];
  assign N1378 = ~sel_i[140];
  assign N1383 = ~sel_i[142];
  assign N1388 = ~sel_i[144];
  assign N1393 = ~sel_i[146];
  assign N1398 = ~sel_i[148];
  assign N1403 = ~sel_i[150];
  assign N1408 = ~sel_i[152];
  assign N1413 = ~sel_i[154];
  assign N1418 = ~sel_i[156];
  assign N1423 = ~sel_i[158];
  assign N1428 = ~sel_i[160];
  assign N1433 = ~sel_i[162];
  assign N1438 = ~sel_i[164];
  assign N1443 = ~sel_i[166];
  assign N1448 = ~sel_i[168];
  assign N1453 = ~sel_i[170];
  assign N1458 = ~sel_i[172];
  assign N1463 = ~sel_i[174];
  assign N1468 = ~sel_i[176];
  assign N1473 = ~sel_i[178];
  assign N1478 = ~sel_i[180];
  assign N1483 = ~sel_i[182];
  assign N1488 = ~sel_i[184];
  assign N1493 = ~sel_i[186];
  assign N1498 = ~sel_i[188];
  assign N1503 = ~sel_i[190];
  assign N1508 = ~sel_i[192];
  assign N1513 = ~sel_i[194];
  assign N1518 = ~sel_i[196];
  assign N1523 = ~sel_i[198];
  assign N1528 = ~sel_i[200];
  assign N1533 = ~sel_i[202];
  assign N1538 = ~sel_i[204];
  assign N1543 = ~sel_i[206];
  assign N1548 = ~sel_i[208];
  assign N1553 = ~sel_i[210];
  assign N1558 = ~sel_i[212];
  assign N1563 = ~sel_i[214];
  assign N1568 = ~sel_i[216];
  assign N1573 = ~sel_i[218];
  assign N1578 = ~sel_i[220];
  assign N1583 = ~sel_i[222];
  assign N1588 = ~sel_i[224];
  assign N1593 = ~sel_i[226];
  assign N1598 = ~sel_i[228];
  assign N1603 = ~sel_i[230];
  assign N1608 = ~sel_i[232];
  assign N1613 = ~sel_i[234];
  assign N1618 = ~sel_i[236];
  assign N1623 = ~sel_i[238];
  assign N1628 = ~sel_i[240];
  assign N1633 = ~sel_i[242];
  assign N1638 = ~sel_i[244];
  assign N1643 = ~sel_i[246];
  assign N1648 = ~sel_i[248];
  assign N1653 = ~sel_i[250];
  assign N1658 = ~sel_i[252];
  assign N1663 = ~sel_i[254];
  assign N1668 = ~sel_i[256];
  assign N1673 = ~sel_i[258];
  assign N1678 = ~sel_i[260];
  assign N1683 = ~sel_i[262];
  assign N1688 = ~sel_i[264];
  assign N1693 = ~sel_i[266];
  assign N1698 = ~sel_i[268];
  assign N1703 = ~sel_i[270];
  assign N1708 = ~sel_i[272];
  assign N1713 = ~sel_i[274];
  assign N1718 = ~sel_i[276];
  assign N1723 = ~sel_i[278];
  assign N1728 = ~sel_i[280];
  assign N1733 = ~sel_i[282];
  assign N1738 = ~sel_i[284];
  assign N1743 = ~sel_i[286];
  assign N1748 = ~sel_i[288];
  assign N1753 = ~sel_i[290];
  assign N1758 = ~sel_i[292];
  assign N1763 = ~sel_i[294];
  assign N1768 = ~sel_i[296];
  assign N1773 = ~sel_i[298];
  assign N1778 = ~sel_i[300];
  assign N1783 = ~sel_i[302];
  assign N1788 = ~sel_i[304];
  assign N1793 = ~sel_i[306];
  assign N1798 = ~sel_i[308];
  assign N1803 = ~sel_i[310];
  assign N1808 = ~sel_i[312];
  assign N1813 = ~sel_i[314];
  assign N1818 = ~sel_i[316];
  assign N1823 = ~sel_i[318];
  assign N1828 = ~sel_i[320];
  assign N1833 = ~sel_i[322];
  assign N1838 = ~sel_i[324];
  assign N1843 = ~sel_i[326];
  assign N1848 = ~sel_i[328];
  assign N1853 = ~sel_i[330];
  assign N1858 = ~sel_i[332];
  assign N1863 = ~sel_i[334];
  assign N1868 = ~sel_i[336];
  assign N1873 = ~sel_i[338];
  assign N1878 = ~sel_i[340];
  assign N1883 = ~sel_i[342];
  assign N1888 = ~sel_i[344];
  assign N1893 = ~sel_i[346];
  assign N1898 = ~sel_i[348];
  assign N1903 = ~sel_i[350];
  assign N1908 = ~sel_i[352];
  assign N1913 = ~sel_i[354];
  assign N1918 = ~sel_i[356];
  assign N1923 = ~sel_i[358];
  assign N1928 = ~sel_i[360];
  assign N1933 = ~sel_i[362];
  assign N1938 = ~sel_i[364];
  assign N1943 = ~sel_i[366];
  assign N1948 = ~sel_i[368];
  assign N1953 = ~sel_i[370];
  assign N1958 = ~sel_i[372];
  assign N1963 = ~sel_i[374];
  assign N1968 = ~sel_i[376];
  assign N1973 = ~sel_i[378];
  assign N1978 = ~sel_i[380];
  assign N1983 = ~sel_i[382];
  assign N1988 = ~sel_i[384];
  assign N1993 = ~sel_i[386];
  assign N1998 = ~sel_i[388];
  assign N2003 = ~sel_i[390];
  assign N2008 = ~sel_i[392];
  assign N2013 = ~sel_i[394];
  assign N2018 = ~sel_i[396];
  assign N2023 = ~sel_i[398];
  assign N2028 = ~sel_i[400];
  assign N2033 = ~sel_i[402];
  assign N2038 = ~sel_i[404];
  assign N2043 = ~sel_i[406];
  assign N2048 = ~sel_i[408];
  assign N2053 = ~sel_i[410];
  assign N2058 = ~sel_i[412];
  assign N2063 = ~sel_i[414];
  assign N2068 = ~sel_i[416];
  assign N2073 = ~sel_i[418];
  assign N2078 = ~sel_i[420];
  assign N2083 = ~sel_i[422];
  assign N2088 = ~sel_i[424];
  assign N2093 = ~sel_i[426];
  assign N2098 = ~sel_i[428];
  assign N2103 = ~sel_i[430];
  assign N2108 = ~sel_i[432];
  assign N2113 = ~sel_i[434];
  assign N2118 = ~sel_i[436];
  assign N2123 = ~sel_i[438];
  assign N2128 = ~sel_i[440];
  assign N2133 = ~sel_i[442];
  assign N2138 = ~sel_i[444];
  assign N2143 = ~sel_i[446];
  assign N2148 = ~sel_i[448];
  assign N2153 = ~sel_i[450];
  assign N2158 = ~sel_i[452];
  assign N2163 = ~sel_i[454];
  assign N2168 = ~sel_i[456];
  assign N2173 = ~sel_i[458];
  assign N2178 = ~sel_i[460];
  assign N2183 = ~sel_i[462];
  assign N2188 = ~sel_i[464];
  assign N2193 = ~sel_i[466];
  assign N2198 = ~sel_i[468];
  assign N2203 = ~sel_i[470];
  assign N2208 = ~sel_i[472];
  assign N2213 = ~sel_i[474];
  assign N2218 = ~sel_i[476];
  assign N2223 = ~sel_i[478];
  assign N2228 = ~sel_i[480];
  assign N2233 = ~sel_i[482];
  assign N2238 = ~sel_i[484];
  assign N2243 = ~sel_i[486];
  assign N2248 = ~sel_i[488];
  assign N2253 = ~sel_i[490];
  assign N2258 = ~sel_i[492];
  assign N2263 = ~sel_i[494];
  assign N2268 = ~sel_i[496];
  assign N2273 = ~sel_i[498];
  assign N2278 = ~sel_i[500];
  assign N2283 = ~sel_i[502];
  assign N2288 = ~sel_i[504];
  assign N2293 = ~sel_i[506];
  assign N2298 = ~sel_i[508];
  assign N2303 = ~sel_i[510];
  assign N2308 = ~sel_i[512];
  assign N2313 = ~sel_i[514];
  assign N2318 = ~sel_i[516];
  assign N2323 = ~sel_i[518];
  assign N2328 = ~sel_i[520];
  assign N2333 = ~sel_i[522];
  assign N2338 = ~sel_i[524];
  assign N2343 = ~sel_i[526];
  assign N2348 = ~sel_i[528];
  assign N2353 = ~sel_i[530];
  assign N2358 = ~sel_i[532];
  assign N2363 = ~sel_i[534];
  assign N2368 = ~sel_i[536];
  assign N2373 = ~sel_i[538];
  assign N2378 = ~sel_i[540];
  assign N2383 = ~sel_i[542];
  assign N2388 = ~sel_i[544];
  assign N2393 = ~sel_i[546];
  assign N2398 = ~sel_i[548];
  assign N2403 = ~sel_i[550];
  assign N2408 = ~sel_i[552];
  assign N2413 = ~sel_i[554];
  assign N2418 = ~sel_i[556];
  assign N2423 = ~sel_i[558];
  assign N2428 = ~sel_i[560];
  assign N2433 = ~sel_i[562];
  assign N2438 = ~sel_i[564];
  assign N2443 = ~sel_i[566];
  assign N2448 = ~sel_i[568];
  assign N2453 = ~sel_i[570];
  assign N2458 = ~sel_i[572];
  assign N2463 = ~sel_i[574];
  assign N2468 = ~sel_i[576];
  assign N2473 = ~sel_i[578];
  assign N2478 = ~sel_i[580];
  assign N2483 = ~sel_i[582];
  assign N2488 = ~sel_i[584];
  assign N2493 = ~sel_i[586];
  assign N2498 = ~sel_i[588];
  assign N2503 = ~sel_i[590];
  assign N2508 = ~sel_i[592];
  assign N2513 = ~sel_i[594];
  assign N2518 = ~sel_i[596];
  assign N2523 = ~sel_i[598];
  assign N2528 = ~sel_i[600];
  assign N2533 = ~sel_i[602];
  assign N2538 = ~sel_i[604];
  assign N2543 = ~sel_i[606];
  assign N2548 = ~sel_i[608];
  assign N2553 = ~sel_i[610];
  assign N2558 = ~sel_i[612];
  assign N2563 = ~sel_i[614];
  assign N2568 = ~sel_i[616];
  assign N2573 = ~sel_i[618];
  assign N2578 = ~sel_i[620];
  assign N2583 = ~sel_i[622];
  assign N2588 = ~sel_i[624];
  assign N2593 = ~sel_i[626];
  assign N2598 = ~sel_i[628];
  assign N2603 = ~sel_i[630];
  assign N2608 = ~sel_i[632];
  assign N2613 = ~sel_i[634];
  assign N2618 = ~sel_i[636];
  assign N2623 = ~sel_i[638];
  assign N2628 = ~sel_i[640];
  assign N2633 = ~sel_i[642];
  assign N2638 = ~sel_i[644];
  assign N2643 = ~sel_i[646];
  assign N2648 = ~sel_i[648];
  assign N2653 = ~sel_i[650];
  assign N2658 = ~sel_i[652];
  assign N2663 = ~sel_i[654];
  assign N2668 = ~sel_i[656];
  assign N2673 = ~sel_i[658];
  assign N2678 = ~sel_i[660];
  assign N2683 = ~sel_i[662];
  assign N2688 = ~sel_i[664];
  assign N2693 = ~sel_i[666];
  assign N2698 = ~sel_i[668];
  assign N2703 = ~sel_i[670];
  assign N2708 = ~sel_i[672];
  assign N2713 = ~sel_i[674];
  assign N2718 = ~sel_i[676];
  assign N2723 = ~sel_i[678];
  assign N2728 = ~sel_i[680];
  assign N2733 = ~sel_i[682];
  assign N2738 = ~sel_i[684];
  assign N2743 = ~sel_i[686];
  assign N2748 = ~sel_i[688];
  assign N2753 = ~sel_i[690];
  assign N2758 = ~sel_i[692];
  assign N2763 = ~sel_i[694];
  assign N2768 = ~sel_i[696];
  assign N2773 = ~sel_i[698];
  assign N2778 = ~sel_i[700];
  assign N2783 = ~sel_i[702];
  assign N2788 = ~sel_i[704];
  assign N2793 = ~sel_i[706];
  assign N2798 = ~sel_i[708];
  assign N2803 = ~sel_i[710];
  assign N2808 = ~sel_i[712];
  assign N2813 = ~sel_i[714];
  assign N2818 = ~sel_i[716];
  assign N2823 = ~sel_i[718];
  assign N2828 = ~sel_i[720];
  assign N2833 = ~sel_i[722];
  assign N2838 = ~sel_i[724];
  assign N2843 = ~sel_i[726];
  assign N2848 = ~sel_i[728];
  assign N2853 = ~sel_i[730];
  assign N2858 = ~sel_i[732];
  assign N2863 = ~sel_i[734];
  assign N2868 = ~sel_i[736];
  assign N2873 = ~sel_i[738];
  assign N2878 = ~sel_i[740];
  assign N2883 = ~sel_i[742];
  assign N2888 = ~sel_i[744];
  assign N2893 = ~sel_i[746];
  assign N2898 = ~sel_i[748];
  assign N2903 = ~sel_i[750];
  assign N2908 = ~sel_i[752];
  assign N2913 = ~sel_i[754];
  assign N2918 = ~sel_i[756];
  assign N2923 = ~sel_i[758];
  assign N2928 = ~sel_i[760];
  assign N2933 = ~sel_i[762];
  assign N2938 = ~sel_i[764];
  assign N2943 = ~sel_i[766];
  assign N2948 = ~sel_i[768];
  assign N2953 = ~sel_i[770];
  assign N2958 = ~sel_i[772];
  assign N2963 = ~sel_i[774];
  assign N2968 = ~sel_i[776];
  assign N2973 = ~sel_i[778];
  assign N2978 = ~sel_i[780];
  assign N2983 = ~sel_i[782];
  assign N2988 = ~sel_i[784];
  assign N2993 = ~sel_i[786];
  assign N2998 = ~sel_i[788];
  assign N3003 = ~sel_i[790];
  assign N3008 = ~sel_i[792];
  assign N3013 = ~sel_i[794];
  assign N3018 = ~sel_i[796];
  assign N3023 = ~sel_i[798];
  assign N3028 = ~sel_i[800];
  assign N3033 = ~sel_i[802];
  assign N3038 = ~sel_i[804];
  assign N3043 = ~sel_i[806];
  assign N3048 = ~sel_i[808];
  assign N3053 = ~sel_i[810];
  assign N3058 = ~sel_i[812];
  assign N3063 = ~sel_i[814];
  assign N3068 = ~sel_i[816];
  assign N3073 = ~sel_i[818];
  assign N3078 = ~sel_i[820];
  assign N3083 = ~sel_i[822];
  assign N3088 = ~sel_i[824];
  assign N3093 = ~sel_i[826];
  assign N3098 = ~sel_i[828];
  assign N3103 = ~sel_i[830];
  assign N3108 = ~sel_i[832];
  assign N3113 = ~sel_i[834];
  assign N3118 = ~sel_i[836];
  assign N3123 = ~sel_i[838];
  assign N3128 = ~sel_i[840];
  assign N3133 = ~sel_i[842];
  assign N3138 = ~sel_i[844];
  assign N3143 = ~sel_i[846];
  assign N3148 = ~sel_i[848];
  assign N3153 = ~sel_i[850];
  assign N3158 = ~sel_i[852];
  assign N3163 = ~sel_i[854];
  assign N3168 = ~sel_i[856];
  assign N3173 = ~sel_i[858];
  assign N3178 = ~sel_i[860];
  assign N3183 = ~sel_i[862];
  assign N3188 = ~sel_i[864];
  assign N3193 = ~sel_i[866];
  assign N3198 = ~sel_i[868];
  assign N3203 = ~sel_i[870];
  assign N3208 = ~sel_i[872];
  assign N3213 = ~sel_i[874];
  assign N3218 = ~sel_i[876];
  assign N3223 = ~sel_i[878];
  assign N3228 = ~sel_i[880];
  assign N3233 = ~sel_i[882];
  assign N3238 = ~sel_i[884];
  assign N3243 = ~sel_i[886];
  assign N3248 = ~sel_i[888];
  assign N3253 = ~sel_i[890];
  assign N3258 = ~sel_i[892];
  assign N3263 = ~sel_i[894];
  assign N3268 = ~sel_i[896];
  assign N3273 = ~sel_i[898];
  assign N3278 = ~sel_i[900];
  assign N3283 = ~sel_i[902];
  assign N3288 = ~sel_i[904];
  assign N3293 = ~sel_i[906];
  assign N3298 = ~sel_i[908];
  assign N3303 = ~sel_i[910];
  assign N3308 = ~sel_i[912];
  assign N3313 = ~sel_i[914];
  assign N3318 = ~sel_i[916];
  assign N3323 = ~sel_i[918];
  assign N3328 = ~sel_i[920];
  assign N3333 = ~sel_i[922];
  assign N3338 = ~sel_i[924];
  assign N3343 = ~sel_i[926];
  assign N3348 = ~sel_i[928];
  assign N3353 = ~sel_i[930];
  assign N3358 = ~sel_i[932];
  assign N3363 = ~sel_i[934];
  assign N3368 = ~sel_i[936];
  assign N3373 = ~sel_i[938];
  assign N3378 = ~sel_i[940];
  assign N3383 = ~sel_i[942];
  assign N3388 = ~sel_i[944];
  assign N3393 = ~sel_i[946];
  assign N3398 = ~sel_i[948];
  assign N3403 = ~sel_i[950];
  assign N3408 = ~sel_i[952];
  assign N3413 = ~sel_i[954];
  assign N3418 = ~sel_i[956];
  assign N3423 = ~sel_i[958];
  assign N3428 = ~sel_i[960];
  assign N3433 = ~sel_i[962];
  assign N3438 = ~sel_i[964];
  assign N3443 = ~sel_i[966];
  assign N3448 = ~sel_i[968];
  assign N3453 = ~sel_i[970];
  assign N3458 = ~sel_i[972];
  assign N3463 = ~sel_i[974];
  assign N3468 = ~sel_i[976];
  assign N3473 = ~sel_i[978];
  assign N3478 = ~sel_i[980];
  assign N3483 = ~sel_i[982];
  assign N3488 = ~sel_i[984];
  assign N3493 = ~sel_i[986];
  assign N3498 = ~sel_i[988];
  assign N3503 = ~sel_i[990];
  assign N3508 = ~sel_i[992];
  assign N3513 = ~sel_i[994];
  assign N3518 = ~sel_i[996];
  assign N3523 = ~sel_i[998];
  assign N3528 = ~sel_i[1000];
  assign N3533 = ~sel_i[1002];
  assign N3538 = ~sel_i[1004];
  assign N3543 = ~sel_i[1006];
  assign N3548 = ~sel_i[1008];
  assign N3553 = ~sel_i[1010];
  assign N3558 = ~sel_i[1012];
  assign N3563 = ~sel_i[1014];
  assign N3568 = ~sel_i[1016];
  assign N3573 = ~sel_i[1018];
  assign N3578 = ~sel_i[1020];
  assign N3583 = ~sel_i[1022];
  assign { r_n_0__63_, r_n_0__62_, r_n_0__61_, r_n_0__60_, r_n_0__59_, r_n_0__58_, r_n_0__57_, r_n_0__56_, r_n_0__55_, r_n_0__54_, r_n_0__53_, r_n_0__52_, r_n_0__51_, r_n_0__50_, r_n_0__49_, r_n_0__48_, r_n_0__47_, r_n_0__46_, r_n_0__45_, r_n_0__44_, r_n_0__43_, r_n_0__42_, r_n_0__41_, r_n_0__40_, r_n_0__39_, r_n_0__38_, r_n_0__37_, r_n_0__36_, r_n_0__35_, r_n_0__34_, r_n_0__33_, r_n_0__32_, r_n_0__31_, r_n_0__30_, r_n_0__29_, r_n_0__28_, r_n_0__27_, r_n_0__26_, r_n_0__25_, r_n_0__24_, r_n_0__23_, r_n_0__22_, r_n_0__21_, r_n_0__20_, r_n_0__19_, r_n_0__18_, r_n_0__17_, r_n_0__16_, r_n_0__15_, r_n_0__14_, r_n_0__13_, r_n_0__12_, r_n_0__11_, r_n_0__10_, r_n_0__9_, r_n_0__8_, r_n_0__7_, r_n_0__6_, r_n_0__5_, r_n_0__4_, r_n_0__3_, r_n_0__2_, r_n_0__1_, r_n_0__0_ } = (N0)? { r_1__63_, r_1__62_, r_1__61_, r_1__60_, r_1__59_, r_1__58_, r_1__57_, r_1__56_, r_1__55_, r_1__54_, r_1__53_, r_1__52_, r_1__51_, r_1__50_, r_1__49_, r_1__48_, r_1__47_, r_1__46_, r_1__45_, r_1__44_, r_1__43_, r_1__42_, r_1__41_, r_1__40_, r_1__39_, r_1__38_, r_1__37_, r_1__36_, r_1__35_, r_1__34_, r_1__33_, r_1__32_, r_1__31_, r_1__30_, r_1__29_, r_1__28_, r_1__27_, r_1__26_, r_1__25_, r_1__24_, r_1__23_, r_1__22_, r_1__21_, r_1__20_, r_1__19_, r_1__18_, r_1__17_, r_1__16_, r_1__15_, r_1__14_, r_1__13_, r_1__12_, r_1__11_, r_1__10_, r_1__9_, r_1__8_, r_1__7_, r_1__6_, r_1__5_, r_1__4_, r_1__3_, r_1__2_, r_1__1_, r_1__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N1)? data_i : 1'b0;
  assign N0 = sel_i[0];
  assign N1 = N1028;
  assign { r_n_1__63_, r_n_1__62_, r_n_1__61_, r_n_1__60_, r_n_1__59_, r_n_1__58_, r_n_1__57_, r_n_1__56_, r_n_1__55_, r_n_1__54_, r_n_1__53_, r_n_1__52_, r_n_1__51_, r_n_1__50_, r_n_1__49_, r_n_1__48_, r_n_1__47_, r_n_1__46_, r_n_1__45_, r_n_1__44_, r_n_1__43_, r_n_1__42_, r_n_1__41_, r_n_1__40_, r_n_1__39_, r_n_1__38_, r_n_1__37_, r_n_1__36_, r_n_1__35_, r_n_1__34_, r_n_1__33_, r_n_1__32_, r_n_1__31_, r_n_1__30_, r_n_1__29_, r_n_1__28_, r_n_1__27_, r_n_1__26_, r_n_1__25_, r_n_1__24_, r_n_1__23_, r_n_1__22_, r_n_1__21_, r_n_1__20_, r_n_1__19_, r_n_1__18_, r_n_1__17_, r_n_1__16_, r_n_1__15_, r_n_1__14_, r_n_1__13_, r_n_1__12_, r_n_1__11_, r_n_1__10_, r_n_1__9_, r_n_1__8_, r_n_1__7_, r_n_1__6_, r_n_1__5_, r_n_1__4_, r_n_1__3_, r_n_1__2_, r_n_1__1_, r_n_1__0_ } = (N2)? { r_2__63_, r_2__62_, r_2__61_, r_2__60_, r_2__59_, r_2__58_, r_2__57_, r_2__56_, r_2__55_, r_2__54_, r_2__53_, r_2__52_, r_2__51_, r_2__50_, r_2__49_, r_2__48_, r_2__47_, r_2__46_, r_2__45_, r_2__44_, r_2__43_, r_2__42_, r_2__41_, r_2__40_, r_2__39_, r_2__38_, r_2__37_, r_2__36_, r_2__35_, r_2__34_, r_2__33_, r_2__32_, r_2__31_, r_2__30_, r_2__29_, r_2__28_, r_2__27_, r_2__26_, r_2__25_, r_2__24_, r_2__23_, r_2__22_, r_2__21_, r_2__20_, r_2__19_, r_2__18_, r_2__17_, r_2__16_, r_2__15_, r_2__14_, r_2__13_, r_2__12_, r_2__11_, r_2__10_, r_2__9_, r_2__8_, r_2__7_, r_2__6_, r_2__5_, r_2__4_, r_2__3_, r_2__2_, r_2__1_, r_2__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N3)? data_i : 1'b0;
  assign N2 = sel_i[2];
  assign N3 = N1033;
  assign { r_n_2__63_, r_n_2__62_, r_n_2__61_, r_n_2__60_, r_n_2__59_, r_n_2__58_, r_n_2__57_, r_n_2__56_, r_n_2__55_, r_n_2__54_, r_n_2__53_, r_n_2__52_, r_n_2__51_, r_n_2__50_, r_n_2__49_, r_n_2__48_, r_n_2__47_, r_n_2__46_, r_n_2__45_, r_n_2__44_, r_n_2__43_, r_n_2__42_, r_n_2__41_, r_n_2__40_, r_n_2__39_, r_n_2__38_, r_n_2__37_, r_n_2__36_, r_n_2__35_, r_n_2__34_, r_n_2__33_, r_n_2__32_, r_n_2__31_, r_n_2__30_, r_n_2__29_, r_n_2__28_, r_n_2__27_, r_n_2__26_, r_n_2__25_, r_n_2__24_, r_n_2__23_, r_n_2__22_, r_n_2__21_, r_n_2__20_, r_n_2__19_, r_n_2__18_, r_n_2__17_, r_n_2__16_, r_n_2__15_, r_n_2__14_, r_n_2__13_, r_n_2__12_, r_n_2__11_, r_n_2__10_, r_n_2__9_, r_n_2__8_, r_n_2__7_, r_n_2__6_, r_n_2__5_, r_n_2__4_, r_n_2__3_, r_n_2__2_, r_n_2__1_, r_n_2__0_ } = (N4)? { r_3__63_, r_3__62_, r_3__61_, r_3__60_, r_3__59_, r_3__58_, r_3__57_, r_3__56_, r_3__55_, r_3__54_, r_3__53_, r_3__52_, r_3__51_, r_3__50_, r_3__49_, r_3__48_, r_3__47_, r_3__46_, r_3__45_, r_3__44_, r_3__43_, r_3__42_, r_3__41_, r_3__40_, r_3__39_, r_3__38_, r_3__37_, r_3__36_, r_3__35_, r_3__34_, r_3__33_, r_3__32_, r_3__31_, r_3__30_, r_3__29_, r_3__28_, r_3__27_, r_3__26_, r_3__25_, r_3__24_, r_3__23_, r_3__22_, r_3__21_, r_3__20_, r_3__19_, r_3__18_, r_3__17_, r_3__16_, r_3__15_, r_3__14_, r_3__13_, r_3__12_, r_3__11_, r_3__10_, r_3__9_, r_3__8_, r_3__7_, r_3__6_, r_3__5_, r_3__4_, r_3__3_, r_3__2_, r_3__1_, r_3__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N5)? data_i : 1'b0;
  assign N4 = sel_i[4];
  assign N5 = N1038;
  assign { r_n_3__63_, r_n_3__62_, r_n_3__61_, r_n_3__60_, r_n_3__59_, r_n_3__58_, r_n_3__57_, r_n_3__56_, r_n_3__55_, r_n_3__54_, r_n_3__53_, r_n_3__52_, r_n_3__51_, r_n_3__50_, r_n_3__49_, r_n_3__48_, r_n_3__47_, r_n_3__46_, r_n_3__45_, r_n_3__44_, r_n_3__43_, r_n_3__42_, r_n_3__41_, r_n_3__40_, r_n_3__39_, r_n_3__38_, r_n_3__37_, r_n_3__36_, r_n_3__35_, r_n_3__34_, r_n_3__33_, r_n_3__32_, r_n_3__31_, r_n_3__30_, r_n_3__29_, r_n_3__28_, r_n_3__27_, r_n_3__26_, r_n_3__25_, r_n_3__24_, r_n_3__23_, r_n_3__22_, r_n_3__21_, r_n_3__20_, r_n_3__19_, r_n_3__18_, r_n_3__17_, r_n_3__16_, r_n_3__15_, r_n_3__14_, r_n_3__13_, r_n_3__12_, r_n_3__11_, r_n_3__10_, r_n_3__9_, r_n_3__8_, r_n_3__7_, r_n_3__6_, r_n_3__5_, r_n_3__4_, r_n_3__3_, r_n_3__2_, r_n_3__1_, r_n_3__0_ } = (N6)? { r_4__63_, r_4__62_, r_4__61_, r_4__60_, r_4__59_, r_4__58_, r_4__57_, r_4__56_, r_4__55_, r_4__54_, r_4__53_, r_4__52_, r_4__51_, r_4__50_, r_4__49_, r_4__48_, r_4__47_, r_4__46_, r_4__45_, r_4__44_, r_4__43_, r_4__42_, r_4__41_, r_4__40_, r_4__39_, r_4__38_, r_4__37_, r_4__36_, r_4__35_, r_4__34_, r_4__33_, r_4__32_, r_4__31_, r_4__30_, r_4__29_, r_4__28_, r_4__27_, r_4__26_, r_4__25_, r_4__24_, r_4__23_, r_4__22_, r_4__21_, r_4__20_, r_4__19_, r_4__18_, r_4__17_, r_4__16_, r_4__15_, r_4__14_, r_4__13_, r_4__12_, r_4__11_, r_4__10_, r_4__9_, r_4__8_, r_4__7_, r_4__6_, r_4__5_, r_4__4_, r_4__3_, r_4__2_, r_4__1_, r_4__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N7)? data_i : 1'b0;
  assign N6 = sel_i[6];
  assign N7 = N1043;
  assign { r_n_4__63_, r_n_4__62_, r_n_4__61_, r_n_4__60_, r_n_4__59_, r_n_4__58_, r_n_4__57_, r_n_4__56_, r_n_4__55_, r_n_4__54_, r_n_4__53_, r_n_4__52_, r_n_4__51_, r_n_4__50_, r_n_4__49_, r_n_4__48_, r_n_4__47_, r_n_4__46_, r_n_4__45_, r_n_4__44_, r_n_4__43_, r_n_4__42_, r_n_4__41_, r_n_4__40_, r_n_4__39_, r_n_4__38_, r_n_4__37_, r_n_4__36_, r_n_4__35_, r_n_4__34_, r_n_4__33_, r_n_4__32_, r_n_4__31_, r_n_4__30_, r_n_4__29_, r_n_4__28_, r_n_4__27_, r_n_4__26_, r_n_4__25_, r_n_4__24_, r_n_4__23_, r_n_4__22_, r_n_4__21_, r_n_4__20_, r_n_4__19_, r_n_4__18_, r_n_4__17_, r_n_4__16_, r_n_4__15_, r_n_4__14_, r_n_4__13_, r_n_4__12_, r_n_4__11_, r_n_4__10_, r_n_4__9_, r_n_4__8_, r_n_4__7_, r_n_4__6_, r_n_4__5_, r_n_4__4_, r_n_4__3_, r_n_4__2_, r_n_4__1_, r_n_4__0_ } = (N8)? { r_5__63_, r_5__62_, r_5__61_, r_5__60_, r_5__59_, r_5__58_, r_5__57_, r_5__56_, r_5__55_, r_5__54_, r_5__53_, r_5__52_, r_5__51_, r_5__50_, r_5__49_, r_5__48_, r_5__47_, r_5__46_, r_5__45_, r_5__44_, r_5__43_, r_5__42_, r_5__41_, r_5__40_, r_5__39_, r_5__38_, r_5__37_, r_5__36_, r_5__35_, r_5__34_, r_5__33_, r_5__32_, r_5__31_, r_5__30_, r_5__29_, r_5__28_, r_5__27_, r_5__26_, r_5__25_, r_5__24_, r_5__23_, r_5__22_, r_5__21_, r_5__20_, r_5__19_, r_5__18_, r_5__17_, r_5__16_, r_5__15_, r_5__14_, r_5__13_, r_5__12_, r_5__11_, r_5__10_, r_5__9_, r_5__8_, r_5__7_, r_5__6_, r_5__5_, r_5__4_, r_5__3_, r_5__2_, r_5__1_, r_5__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N9)? data_i : 1'b0;
  assign N8 = sel_i[8];
  assign N9 = N1048;
  assign { r_n_5__63_, r_n_5__62_, r_n_5__61_, r_n_5__60_, r_n_5__59_, r_n_5__58_, r_n_5__57_, r_n_5__56_, r_n_5__55_, r_n_5__54_, r_n_5__53_, r_n_5__52_, r_n_5__51_, r_n_5__50_, r_n_5__49_, r_n_5__48_, r_n_5__47_, r_n_5__46_, r_n_5__45_, r_n_5__44_, r_n_5__43_, r_n_5__42_, r_n_5__41_, r_n_5__40_, r_n_5__39_, r_n_5__38_, r_n_5__37_, r_n_5__36_, r_n_5__35_, r_n_5__34_, r_n_5__33_, r_n_5__32_, r_n_5__31_, r_n_5__30_, r_n_5__29_, r_n_5__28_, r_n_5__27_, r_n_5__26_, r_n_5__25_, r_n_5__24_, r_n_5__23_, r_n_5__22_, r_n_5__21_, r_n_5__20_, r_n_5__19_, r_n_5__18_, r_n_5__17_, r_n_5__16_, r_n_5__15_, r_n_5__14_, r_n_5__13_, r_n_5__12_, r_n_5__11_, r_n_5__10_, r_n_5__9_, r_n_5__8_, r_n_5__7_, r_n_5__6_, r_n_5__5_, r_n_5__4_, r_n_5__3_, r_n_5__2_, r_n_5__1_, r_n_5__0_ } = (N10)? { r_6__63_, r_6__62_, r_6__61_, r_6__60_, r_6__59_, r_6__58_, r_6__57_, r_6__56_, r_6__55_, r_6__54_, r_6__53_, r_6__52_, r_6__51_, r_6__50_, r_6__49_, r_6__48_, r_6__47_, r_6__46_, r_6__45_, r_6__44_, r_6__43_, r_6__42_, r_6__41_, r_6__40_, r_6__39_, r_6__38_, r_6__37_, r_6__36_, r_6__35_, r_6__34_, r_6__33_, r_6__32_, r_6__31_, r_6__30_, r_6__29_, r_6__28_, r_6__27_, r_6__26_, r_6__25_, r_6__24_, r_6__23_, r_6__22_, r_6__21_, r_6__20_, r_6__19_, r_6__18_, r_6__17_, r_6__16_, r_6__15_, r_6__14_, r_6__13_, r_6__12_, r_6__11_, r_6__10_, r_6__9_, r_6__8_, r_6__7_, r_6__6_, r_6__5_, r_6__4_, r_6__3_, r_6__2_, r_6__1_, r_6__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N11)? data_i : 1'b0;
  assign N10 = sel_i[10];
  assign N11 = N1053;
  assign { r_n_6__63_, r_n_6__62_, r_n_6__61_, r_n_6__60_, r_n_6__59_, r_n_6__58_, r_n_6__57_, r_n_6__56_, r_n_6__55_, r_n_6__54_, r_n_6__53_, r_n_6__52_, r_n_6__51_, r_n_6__50_, r_n_6__49_, r_n_6__48_, r_n_6__47_, r_n_6__46_, r_n_6__45_, r_n_6__44_, r_n_6__43_, r_n_6__42_, r_n_6__41_, r_n_6__40_, r_n_6__39_, r_n_6__38_, r_n_6__37_, r_n_6__36_, r_n_6__35_, r_n_6__34_, r_n_6__33_, r_n_6__32_, r_n_6__31_, r_n_6__30_, r_n_6__29_, r_n_6__28_, r_n_6__27_, r_n_6__26_, r_n_6__25_, r_n_6__24_, r_n_6__23_, r_n_6__22_, r_n_6__21_, r_n_6__20_, r_n_6__19_, r_n_6__18_, r_n_6__17_, r_n_6__16_, r_n_6__15_, r_n_6__14_, r_n_6__13_, r_n_6__12_, r_n_6__11_, r_n_6__10_, r_n_6__9_, r_n_6__8_, r_n_6__7_, r_n_6__6_, r_n_6__5_, r_n_6__4_, r_n_6__3_, r_n_6__2_, r_n_6__1_, r_n_6__0_ } = (N12)? { r_7__63_, r_7__62_, r_7__61_, r_7__60_, r_7__59_, r_7__58_, r_7__57_, r_7__56_, r_7__55_, r_7__54_, r_7__53_, r_7__52_, r_7__51_, r_7__50_, r_7__49_, r_7__48_, r_7__47_, r_7__46_, r_7__45_, r_7__44_, r_7__43_, r_7__42_, r_7__41_, r_7__40_, r_7__39_, r_7__38_, r_7__37_, r_7__36_, r_7__35_, r_7__34_, r_7__33_, r_7__32_, r_7__31_, r_7__30_, r_7__29_, r_7__28_, r_7__27_, r_7__26_, r_7__25_, r_7__24_, r_7__23_, r_7__22_, r_7__21_, r_7__20_, r_7__19_, r_7__18_, r_7__17_, r_7__16_, r_7__15_, r_7__14_, r_7__13_, r_7__12_, r_7__11_, r_7__10_, r_7__9_, r_7__8_, r_7__7_, r_7__6_, r_7__5_, r_7__4_, r_7__3_, r_7__2_, r_7__1_, r_7__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N13)? data_i : 1'b0;
  assign N12 = sel_i[12];
  assign N13 = N1058;
  assign { r_n_7__63_, r_n_7__62_, r_n_7__61_, r_n_7__60_, r_n_7__59_, r_n_7__58_, r_n_7__57_, r_n_7__56_, r_n_7__55_, r_n_7__54_, r_n_7__53_, r_n_7__52_, r_n_7__51_, r_n_7__50_, r_n_7__49_, r_n_7__48_, r_n_7__47_, r_n_7__46_, r_n_7__45_, r_n_7__44_, r_n_7__43_, r_n_7__42_, r_n_7__41_, r_n_7__40_, r_n_7__39_, r_n_7__38_, r_n_7__37_, r_n_7__36_, r_n_7__35_, r_n_7__34_, r_n_7__33_, r_n_7__32_, r_n_7__31_, r_n_7__30_, r_n_7__29_, r_n_7__28_, r_n_7__27_, r_n_7__26_, r_n_7__25_, r_n_7__24_, r_n_7__23_, r_n_7__22_, r_n_7__21_, r_n_7__20_, r_n_7__19_, r_n_7__18_, r_n_7__17_, r_n_7__16_, r_n_7__15_, r_n_7__14_, r_n_7__13_, r_n_7__12_, r_n_7__11_, r_n_7__10_, r_n_7__9_, r_n_7__8_, r_n_7__7_, r_n_7__6_, r_n_7__5_, r_n_7__4_, r_n_7__3_, r_n_7__2_, r_n_7__1_, r_n_7__0_ } = (N14)? { r_8__63_, r_8__62_, r_8__61_, r_8__60_, r_8__59_, r_8__58_, r_8__57_, r_8__56_, r_8__55_, r_8__54_, r_8__53_, r_8__52_, r_8__51_, r_8__50_, r_8__49_, r_8__48_, r_8__47_, r_8__46_, r_8__45_, r_8__44_, r_8__43_, r_8__42_, r_8__41_, r_8__40_, r_8__39_, r_8__38_, r_8__37_, r_8__36_, r_8__35_, r_8__34_, r_8__33_, r_8__32_, r_8__31_, r_8__30_, r_8__29_, r_8__28_, r_8__27_, r_8__26_, r_8__25_, r_8__24_, r_8__23_, r_8__22_, r_8__21_, r_8__20_, r_8__19_, r_8__18_, r_8__17_, r_8__16_, r_8__15_, r_8__14_, r_8__13_, r_8__12_, r_8__11_, r_8__10_, r_8__9_, r_8__8_, r_8__7_, r_8__6_, r_8__5_, r_8__4_, r_8__3_, r_8__2_, r_8__1_, r_8__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N15)? data_i : 1'b0;
  assign N14 = sel_i[14];
  assign N15 = N1063;
  assign { r_n_8__63_, r_n_8__62_, r_n_8__61_, r_n_8__60_, r_n_8__59_, r_n_8__58_, r_n_8__57_, r_n_8__56_, r_n_8__55_, r_n_8__54_, r_n_8__53_, r_n_8__52_, r_n_8__51_, r_n_8__50_, r_n_8__49_, r_n_8__48_, r_n_8__47_, r_n_8__46_, r_n_8__45_, r_n_8__44_, r_n_8__43_, r_n_8__42_, r_n_8__41_, r_n_8__40_, r_n_8__39_, r_n_8__38_, r_n_8__37_, r_n_8__36_, r_n_8__35_, r_n_8__34_, r_n_8__33_, r_n_8__32_, r_n_8__31_, r_n_8__30_, r_n_8__29_, r_n_8__28_, r_n_8__27_, r_n_8__26_, r_n_8__25_, r_n_8__24_, r_n_8__23_, r_n_8__22_, r_n_8__21_, r_n_8__20_, r_n_8__19_, r_n_8__18_, r_n_8__17_, r_n_8__16_, r_n_8__15_, r_n_8__14_, r_n_8__13_, r_n_8__12_, r_n_8__11_, r_n_8__10_, r_n_8__9_, r_n_8__8_, r_n_8__7_, r_n_8__6_, r_n_8__5_, r_n_8__4_, r_n_8__3_, r_n_8__2_, r_n_8__1_, r_n_8__0_ } = (N16)? { r_9__63_, r_9__62_, r_9__61_, r_9__60_, r_9__59_, r_9__58_, r_9__57_, r_9__56_, r_9__55_, r_9__54_, r_9__53_, r_9__52_, r_9__51_, r_9__50_, r_9__49_, r_9__48_, r_9__47_, r_9__46_, r_9__45_, r_9__44_, r_9__43_, r_9__42_, r_9__41_, r_9__40_, r_9__39_, r_9__38_, r_9__37_, r_9__36_, r_9__35_, r_9__34_, r_9__33_, r_9__32_, r_9__31_, r_9__30_, r_9__29_, r_9__28_, r_9__27_, r_9__26_, r_9__25_, r_9__24_, r_9__23_, r_9__22_, r_9__21_, r_9__20_, r_9__19_, r_9__18_, r_9__17_, r_9__16_, r_9__15_, r_9__14_, r_9__13_, r_9__12_, r_9__11_, r_9__10_, r_9__9_, r_9__8_, r_9__7_, r_9__6_, r_9__5_, r_9__4_, r_9__3_, r_9__2_, r_9__1_, r_9__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N17)? data_i : 1'b0;
  assign N16 = sel_i[16];
  assign N17 = N1068;
  assign { r_n_9__63_, r_n_9__62_, r_n_9__61_, r_n_9__60_, r_n_9__59_, r_n_9__58_, r_n_9__57_, r_n_9__56_, r_n_9__55_, r_n_9__54_, r_n_9__53_, r_n_9__52_, r_n_9__51_, r_n_9__50_, r_n_9__49_, r_n_9__48_, r_n_9__47_, r_n_9__46_, r_n_9__45_, r_n_9__44_, r_n_9__43_, r_n_9__42_, r_n_9__41_, r_n_9__40_, r_n_9__39_, r_n_9__38_, r_n_9__37_, r_n_9__36_, r_n_9__35_, r_n_9__34_, r_n_9__33_, r_n_9__32_, r_n_9__31_, r_n_9__30_, r_n_9__29_, r_n_9__28_, r_n_9__27_, r_n_9__26_, r_n_9__25_, r_n_9__24_, r_n_9__23_, r_n_9__22_, r_n_9__21_, r_n_9__20_, r_n_9__19_, r_n_9__18_, r_n_9__17_, r_n_9__16_, r_n_9__15_, r_n_9__14_, r_n_9__13_, r_n_9__12_, r_n_9__11_, r_n_9__10_, r_n_9__9_, r_n_9__8_, r_n_9__7_, r_n_9__6_, r_n_9__5_, r_n_9__4_, r_n_9__3_, r_n_9__2_, r_n_9__1_, r_n_9__0_ } = (N18)? { r_10__63_, r_10__62_, r_10__61_, r_10__60_, r_10__59_, r_10__58_, r_10__57_, r_10__56_, r_10__55_, r_10__54_, r_10__53_, r_10__52_, r_10__51_, r_10__50_, r_10__49_, r_10__48_, r_10__47_, r_10__46_, r_10__45_, r_10__44_, r_10__43_, r_10__42_, r_10__41_, r_10__40_, r_10__39_, r_10__38_, r_10__37_, r_10__36_, r_10__35_, r_10__34_, r_10__33_, r_10__32_, r_10__31_, r_10__30_, r_10__29_, r_10__28_, r_10__27_, r_10__26_, r_10__25_, r_10__24_, r_10__23_, r_10__22_, r_10__21_, r_10__20_, r_10__19_, r_10__18_, r_10__17_, r_10__16_, r_10__15_, r_10__14_, r_10__13_, r_10__12_, r_10__11_, r_10__10_, r_10__9_, r_10__8_, r_10__7_, r_10__6_, r_10__5_, r_10__4_, r_10__3_, r_10__2_, r_10__1_, r_10__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N19)? data_i : 1'b0;
  assign N18 = sel_i[18];
  assign N19 = N1073;
  assign { r_n_10__63_, r_n_10__62_, r_n_10__61_, r_n_10__60_, r_n_10__59_, r_n_10__58_, r_n_10__57_, r_n_10__56_, r_n_10__55_, r_n_10__54_, r_n_10__53_, r_n_10__52_, r_n_10__51_, r_n_10__50_, r_n_10__49_, r_n_10__48_, r_n_10__47_, r_n_10__46_, r_n_10__45_, r_n_10__44_, r_n_10__43_, r_n_10__42_, r_n_10__41_, r_n_10__40_, r_n_10__39_, r_n_10__38_, r_n_10__37_, r_n_10__36_, r_n_10__35_, r_n_10__34_, r_n_10__33_, r_n_10__32_, r_n_10__31_, r_n_10__30_, r_n_10__29_, r_n_10__28_, r_n_10__27_, r_n_10__26_, r_n_10__25_, r_n_10__24_, r_n_10__23_, r_n_10__22_, r_n_10__21_, r_n_10__20_, r_n_10__19_, r_n_10__18_, r_n_10__17_, r_n_10__16_, r_n_10__15_, r_n_10__14_, r_n_10__13_, r_n_10__12_, r_n_10__11_, r_n_10__10_, r_n_10__9_, r_n_10__8_, r_n_10__7_, r_n_10__6_, r_n_10__5_, r_n_10__4_, r_n_10__3_, r_n_10__2_, r_n_10__1_, r_n_10__0_ } = (N20)? { r_11__63_, r_11__62_, r_11__61_, r_11__60_, r_11__59_, r_11__58_, r_11__57_, r_11__56_, r_11__55_, r_11__54_, r_11__53_, r_11__52_, r_11__51_, r_11__50_, r_11__49_, r_11__48_, r_11__47_, r_11__46_, r_11__45_, r_11__44_, r_11__43_, r_11__42_, r_11__41_, r_11__40_, r_11__39_, r_11__38_, r_11__37_, r_11__36_, r_11__35_, r_11__34_, r_11__33_, r_11__32_, r_11__31_, r_11__30_, r_11__29_, r_11__28_, r_11__27_, r_11__26_, r_11__25_, r_11__24_, r_11__23_, r_11__22_, r_11__21_, r_11__20_, r_11__19_, r_11__18_, r_11__17_, r_11__16_, r_11__15_, r_11__14_, r_11__13_, r_11__12_, r_11__11_, r_11__10_, r_11__9_, r_11__8_, r_11__7_, r_11__6_, r_11__5_, r_11__4_, r_11__3_, r_11__2_, r_11__1_, r_11__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N21)? data_i : 1'b0;
  assign N20 = sel_i[20];
  assign N21 = N1078;
  assign { r_n_11__63_, r_n_11__62_, r_n_11__61_, r_n_11__60_, r_n_11__59_, r_n_11__58_, r_n_11__57_, r_n_11__56_, r_n_11__55_, r_n_11__54_, r_n_11__53_, r_n_11__52_, r_n_11__51_, r_n_11__50_, r_n_11__49_, r_n_11__48_, r_n_11__47_, r_n_11__46_, r_n_11__45_, r_n_11__44_, r_n_11__43_, r_n_11__42_, r_n_11__41_, r_n_11__40_, r_n_11__39_, r_n_11__38_, r_n_11__37_, r_n_11__36_, r_n_11__35_, r_n_11__34_, r_n_11__33_, r_n_11__32_, r_n_11__31_, r_n_11__30_, r_n_11__29_, r_n_11__28_, r_n_11__27_, r_n_11__26_, r_n_11__25_, r_n_11__24_, r_n_11__23_, r_n_11__22_, r_n_11__21_, r_n_11__20_, r_n_11__19_, r_n_11__18_, r_n_11__17_, r_n_11__16_, r_n_11__15_, r_n_11__14_, r_n_11__13_, r_n_11__12_, r_n_11__11_, r_n_11__10_, r_n_11__9_, r_n_11__8_, r_n_11__7_, r_n_11__6_, r_n_11__5_, r_n_11__4_, r_n_11__3_, r_n_11__2_, r_n_11__1_, r_n_11__0_ } = (N22)? { r_12__63_, r_12__62_, r_12__61_, r_12__60_, r_12__59_, r_12__58_, r_12__57_, r_12__56_, r_12__55_, r_12__54_, r_12__53_, r_12__52_, r_12__51_, r_12__50_, r_12__49_, r_12__48_, r_12__47_, r_12__46_, r_12__45_, r_12__44_, r_12__43_, r_12__42_, r_12__41_, r_12__40_, r_12__39_, r_12__38_, r_12__37_, r_12__36_, r_12__35_, r_12__34_, r_12__33_, r_12__32_, r_12__31_, r_12__30_, r_12__29_, r_12__28_, r_12__27_, r_12__26_, r_12__25_, r_12__24_, r_12__23_, r_12__22_, r_12__21_, r_12__20_, r_12__19_, r_12__18_, r_12__17_, r_12__16_, r_12__15_, r_12__14_, r_12__13_, r_12__12_, r_12__11_, r_12__10_, r_12__9_, r_12__8_, r_12__7_, r_12__6_, r_12__5_, r_12__4_, r_12__3_, r_12__2_, r_12__1_, r_12__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N23)? data_i : 1'b0;
  assign N22 = sel_i[22];
  assign N23 = N1083;
  assign { r_n_12__63_, r_n_12__62_, r_n_12__61_, r_n_12__60_, r_n_12__59_, r_n_12__58_, r_n_12__57_, r_n_12__56_, r_n_12__55_, r_n_12__54_, r_n_12__53_, r_n_12__52_, r_n_12__51_, r_n_12__50_, r_n_12__49_, r_n_12__48_, r_n_12__47_, r_n_12__46_, r_n_12__45_, r_n_12__44_, r_n_12__43_, r_n_12__42_, r_n_12__41_, r_n_12__40_, r_n_12__39_, r_n_12__38_, r_n_12__37_, r_n_12__36_, r_n_12__35_, r_n_12__34_, r_n_12__33_, r_n_12__32_, r_n_12__31_, r_n_12__30_, r_n_12__29_, r_n_12__28_, r_n_12__27_, r_n_12__26_, r_n_12__25_, r_n_12__24_, r_n_12__23_, r_n_12__22_, r_n_12__21_, r_n_12__20_, r_n_12__19_, r_n_12__18_, r_n_12__17_, r_n_12__16_, r_n_12__15_, r_n_12__14_, r_n_12__13_, r_n_12__12_, r_n_12__11_, r_n_12__10_, r_n_12__9_, r_n_12__8_, r_n_12__7_, r_n_12__6_, r_n_12__5_, r_n_12__4_, r_n_12__3_, r_n_12__2_, r_n_12__1_, r_n_12__0_ } = (N24)? { r_13__63_, r_13__62_, r_13__61_, r_13__60_, r_13__59_, r_13__58_, r_13__57_, r_13__56_, r_13__55_, r_13__54_, r_13__53_, r_13__52_, r_13__51_, r_13__50_, r_13__49_, r_13__48_, r_13__47_, r_13__46_, r_13__45_, r_13__44_, r_13__43_, r_13__42_, r_13__41_, r_13__40_, r_13__39_, r_13__38_, r_13__37_, r_13__36_, r_13__35_, r_13__34_, r_13__33_, r_13__32_, r_13__31_, r_13__30_, r_13__29_, r_13__28_, r_13__27_, r_13__26_, r_13__25_, r_13__24_, r_13__23_, r_13__22_, r_13__21_, r_13__20_, r_13__19_, r_13__18_, r_13__17_, r_13__16_, r_13__15_, r_13__14_, r_13__13_, r_13__12_, r_13__11_, r_13__10_, r_13__9_, r_13__8_, r_13__7_, r_13__6_, r_13__5_, r_13__4_, r_13__3_, r_13__2_, r_13__1_, r_13__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N25)? data_i : 1'b0;
  assign N24 = sel_i[24];
  assign N25 = N1088;
  assign { r_n_13__63_, r_n_13__62_, r_n_13__61_, r_n_13__60_, r_n_13__59_, r_n_13__58_, r_n_13__57_, r_n_13__56_, r_n_13__55_, r_n_13__54_, r_n_13__53_, r_n_13__52_, r_n_13__51_, r_n_13__50_, r_n_13__49_, r_n_13__48_, r_n_13__47_, r_n_13__46_, r_n_13__45_, r_n_13__44_, r_n_13__43_, r_n_13__42_, r_n_13__41_, r_n_13__40_, r_n_13__39_, r_n_13__38_, r_n_13__37_, r_n_13__36_, r_n_13__35_, r_n_13__34_, r_n_13__33_, r_n_13__32_, r_n_13__31_, r_n_13__30_, r_n_13__29_, r_n_13__28_, r_n_13__27_, r_n_13__26_, r_n_13__25_, r_n_13__24_, r_n_13__23_, r_n_13__22_, r_n_13__21_, r_n_13__20_, r_n_13__19_, r_n_13__18_, r_n_13__17_, r_n_13__16_, r_n_13__15_, r_n_13__14_, r_n_13__13_, r_n_13__12_, r_n_13__11_, r_n_13__10_, r_n_13__9_, r_n_13__8_, r_n_13__7_, r_n_13__6_, r_n_13__5_, r_n_13__4_, r_n_13__3_, r_n_13__2_, r_n_13__1_, r_n_13__0_ } = (N26)? { r_14__63_, r_14__62_, r_14__61_, r_14__60_, r_14__59_, r_14__58_, r_14__57_, r_14__56_, r_14__55_, r_14__54_, r_14__53_, r_14__52_, r_14__51_, r_14__50_, r_14__49_, r_14__48_, r_14__47_, r_14__46_, r_14__45_, r_14__44_, r_14__43_, r_14__42_, r_14__41_, r_14__40_, r_14__39_, r_14__38_, r_14__37_, r_14__36_, r_14__35_, r_14__34_, r_14__33_, r_14__32_, r_14__31_, r_14__30_, r_14__29_, r_14__28_, r_14__27_, r_14__26_, r_14__25_, r_14__24_, r_14__23_, r_14__22_, r_14__21_, r_14__20_, r_14__19_, r_14__18_, r_14__17_, r_14__16_, r_14__15_, r_14__14_, r_14__13_, r_14__12_, r_14__11_, r_14__10_, r_14__9_, r_14__8_, r_14__7_, r_14__6_, r_14__5_, r_14__4_, r_14__3_, r_14__2_, r_14__1_, r_14__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N27)? data_i : 1'b0;
  assign N26 = sel_i[26];
  assign N27 = N1093;
  assign { r_n_14__63_, r_n_14__62_, r_n_14__61_, r_n_14__60_, r_n_14__59_, r_n_14__58_, r_n_14__57_, r_n_14__56_, r_n_14__55_, r_n_14__54_, r_n_14__53_, r_n_14__52_, r_n_14__51_, r_n_14__50_, r_n_14__49_, r_n_14__48_, r_n_14__47_, r_n_14__46_, r_n_14__45_, r_n_14__44_, r_n_14__43_, r_n_14__42_, r_n_14__41_, r_n_14__40_, r_n_14__39_, r_n_14__38_, r_n_14__37_, r_n_14__36_, r_n_14__35_, r_n_14__34_, r_n_14__33_, r_n_14__32_, r_n_14__31_, r_n_14__30_, r_n_14__29_, r_n_14__28_, r_n_14__27_, r_n_14__26_, r_n_14__25_, r_n_14__24_, r_n_14__23_, r_n_14__22_, r_n_14__21_, r_n_14__20_, r_n_14__19_, r_n_14__18_, r_n_14__17_, r_n_14__16_, r_n_14__15_, r_n_14__14_, r_n_14__13_, r_n_14__12_, r_n_14__11_, r_n_14__10_, r_n_14__9_, r_n_14__8_, r_n_14__7_, r_n_14__6_, r_n_14__5_, r_n_14__4_, r_n_14__3_, r_n_14__2_, r_n_14__1_, r_n_14__0_ } = (N28)? { r_15__63_, r_15__62_, r_15__61_, r_15__60_, r_15__59_, r_15__58_, r_15__57_, r_15__56_, r_15__55_, r_15__54_, r_15__53_, r_15__52_, r_15__51_, r_15__50_, r_15__49_, r_15__48_, r_15__47_, r_15__46_, r_15__45_, r_15__44_, r_15__43_, r_15__42_, r_15__41_, r_15__40_, r_15__39_, r_15__38_, r_15__37_, r_15__36_, r_15__35_, r_15__34_, r_15__33_, r_15__32_, r_15__31_, r_15__30_, r_15__29_, r_15__28_, r_15__27_, r_15__26_, r_15__25_, r_15__24_, r_15__23_, r_15__22_, r_15__21_, r_15__20_, r_15__19_, r_15__18_, r_15__17_, r_15__16_, r_15__15_, r_15__14_, r_15__13_, r_15__12_, r_15__11_, r_15__10_, r_15__9_, r_15__8_, r_15__7_, r_15__6_, r_15__5_, r_15__4_, r_15__3_, r_15__2_, r_15__1_, r_15__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N29)? data_i : 1'b0;
  assign N28 = sel_i[28];
  assign N29 = N1098;
  assign { r_n_15__63_, r_n_15__62_, r_n_15__61_, r_n_15__60_, r_n_15__59_, r_n_15__58_, r_n_15__57_, r_n_15__56_, r_n_15__55_, r_n_15__54_, r_n_15__53_, r_n_15__52_, r_n_15__51_, r_n_15__50_, r_n_15__49_, r_n_15__48_, r_n_15__47_, r_n_15__46_, r_n_15__45_, r_n_15__44_, r_n_15__43_, r_n_15__42_, r_n_15__41_, r_n_15__40_, r_n_15__39_, r_n_15__38_, r_n_15__37_, r_n_15__36_, r_n_15__35_, r_n_15__34_, r_n_15__33_, r_n_15__32_, r_n_15__31_, r_n_15__30_, r_n_15__29_, r_n_15__28_, r_n_15__27_, r_n_15__26_, r_n_15__25_, r_n_15__24_, r_n_15__23_, r_n_15__22_, r_n_15__21_, r_n_15__20_, r_n_15__19_, r_n_15__18_, r_n_15__17_, r_n_15__16_, r_n_15__15_, r_n_15__14_, r_n_15__13_, r_n_15__12_, r_n_15__11_, r_n_15__10_, r_n_15__9_, r_n_15__8_, r_n_15__7_, r_n_15__6_, r_n_15__5_, r_n_15__4_, r_n_15__3_, r_n_15__2_, r_n_15__1_, r_n_15__0_ } = (N30)? { r_16__63_, r_16__62_, r_16__61_, r_16__60_, r_16__59_, r_16__58_, r_16__57_, r_16__56_, r_16__55_, r_16__54_, r_16__53_, r_16__52_, r_16__51_, r_16__50_, r_16__49_, r_16__48_, r_16__47_, r_16__46_, r_16__45_, r_16__44_, r_16__43_, r_16__42_, r_16__41_, r_16__40_, r_16__39_, r_16__38_, r_16__37_, r_16__36_, r_16__35_, r_16__34_, r_16__33_, r_16__32_, r_16__31_, r_16__30_, r_16__29_, r_16__28_, r_16__27_, r_16__26_, r_16__25_, r_16__24_, r_16__23_, r_16__22_, r_16__21_, r_16__20_, r_16__19_, r_16__18_, r_16__17_, r_16__16_, r_16__15_, r_16__14_, r_16__13_, r_16__12_, r_16__11_, r_16__10_, r_16__9_, r_16__8_, r_16__7_, r_16__6_, r_16__5_, r_16__4_, r_16__3_, r_16__2_, r_16__1_, r_16__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N31)? data_i : 1'b0;
  assign N30 = sel_i[30];
  assign N31 = N1103;
  assign { r_n_16__63_, r_n_16__62_, r_n_16__61_, r_n_16__60_, r_n_16__59_, r_n_16__58_, r_n_16__57_, r_n_16__56_, r_n_16__55_, r_n_16__54_, r_n_16__53_, r_n_16__52_, r_n_16__51_, r_n_16__50_, r_n_16__49_, r_n_16__48_, r_n_16__47_, r_n_16__46_, r_n_16__45_, r_n_16__44_, r_n_16__43_, r_n_16__42_, r_n_16__41_, r_n_16__40_, r_n_16__39_, r_n_16__38_, r_n_16__37_, r_n_16__36_, r_n_16__35_, r_n_16__34_, r_n_16__33_, r_n_16__32_, r_n_16__31_, r_n_16__30_, r_n_16__29_, r_n_16__28_, r_n_16__27_, r_n_16__26_, r_n_16__25_, r_n_16__24_, r_n_16__23_, r_n_16__22_, r_n_16__21_, r_n_16__20_, r_n_16__19_, r_n_16__18_, r_n_16__17_, r_n_16__16_, r_n_16__15_, r_n_16__14_, r_n_16__13_, r_n_16__12_, r_n_16__11_, r_n_16__10_, r_n_16__9_, r_n_16__8_, r_n_16__7_, r_n_16__6_, r_n_16__5_, r_n_16__4_, r_n_16__3_, r_n_16__2_, r_n_16__1_, r_n_16__0_ } = (N32)? { r_17__63_, r_17__62_, r_17__61_, r_17__60_, r_17__59_, r_17__58_, r_17__57_, r_17__56_, r_17__55_, r_17__54_, r_17__53_, r_17__52_, r_17__51_, r_17__50_, r_17__49_, r_17__48_, r_17__47_, r_17__46_, r_17__45_, r_17__44_, r_17__43_, r_17__42_, r_17__41_, r_17__40_, r_17__39_, r_17__38_, r_17__37_, r_17__36_, r_17__35_, r_17__34_, r_17__33_, r_17__32_, r_17__31_, r_17__30_, r_17__29_, r_17__28_, r_17__27_, r_17__26_, r_17__25_, r_17__24_, r_17__23_, r_17__22_, r_17__21_, r_17__20_, r_17__19_, r_17__18_, r_17__17_, r_17__16_, r_17__15_, r_17__14_, r_17__13_, r_17__12_, r_17__11_, r_17__10_, r_17__9_, r_17__8_, r_17__7_, r_17__6_, r_17__5_, r_17__4_, r_17__3_, r_17__2_, r_17__1_, r_17__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N33)? data_i : 1'b0;
  assign N32 = sel_i[32];
  assign N33 = N1108;
  assign { r_n_17__63_, r_n_17__62_, r_n_17__61_, r_n_17__60_, r_n_17__59_, r_n_17__58_, r_n_17__57_, r_n_17__56_, r_n_17__55_, r_n_17__54_, r_n_17__53_, r_n_17__52_, r_n_17__51_, r_n_17__50_, r_n_17__49_, r_n_17__48_, r_n_17__47_, r_n_17__46_, r_n_17__45_, r_n_17__44_, r_n_17__43_, r_n_17__42_, r_n_17__41_, r_n_17__40_, r_n_17__39_, r_n_17__38_, r_n_17__37_, r_n_17__36_, r_n_17__35_, r_n_17__34_, r_n_17__33_, r_n_17__32_, r_n_17__31_, r_n_17__30_, r_n_17__29_, r_n_17__28_, r_n_17__27_, r_n_17__26_, r_n_17__25_, r_n_17__24_, r_n_17__23_, r_n_17__22_, r_n_17__21_, r_n_17__20_, r_n_17__19_, r_n_17__18_, r_n_17__17_, r_n_17__16_, r_n_17__15_, r_n_17__14_, r_n_17__13_, r_n_17__12_, r_n_17__11_, r_n_17__10_, r_n_17__9_, r_n_17__8_, r_n_17__7_, r_n_17__6_, r_n_17__5_, r_n_17__4_, r_n_17__3_, r_n_17__2_, r_n_17__1_, r_n_17__0_ } = (N34)? { r_18__63_, r_18__62_, r_18__61_, r_18__60_, r_18__59_, r_18__58_, r_18__57_, r_18__56_, r_18__55_, r_18__54_, r_18__53_, r_18__52_, r_18__51_, r_18__50_, r_18__49_, r_18__48_, r_18__47_, r_18__46_, r_18__45_, r_18__44_, r_18__43_, r_18__42_, r_18__41_, r_18__40_, r_18__39_, r_18__38_, r_18__37_, r_18__36_, r_18__35_, r_18__34_, r_18__33_, r_18__32_, r_18__31_, r_18__30_, r_18__29_, r_18__28_, r_18__27_, r_18__26_, r_18__25_, r_18__24_, r_18__23_, r_18__22_, r_18__21_, r_18__20_, r_18__19_, r_18__18_, r_18__17_, r_18__16_, r_18__15_, r_18__14_, r_18__13_, r_18__12_, r_18__11_, r_18__10_, r_18__9_, r_18__8_, r_18__7_, r_18__6_, r_18__5_, r_18__4_, r_18__3_, r_18__2_, r_18__1_, r_18__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N35)? data_i : 1'b0;
  assign N34 = sel_i[34];
  assign N35 = N1113;
  assign { r_n_18__63_, r_n_18__62_, r_n_18__61_, r_n_18__60_, r_n_18__59_, r_n_18__58_, r_n_18__57_, r_n_18__56_, r_n_18__55_, r_n_18__54_, r_n_18__53_, r_n_18__52_, r_n_18__51_, r_n_18__50_, r_n_18__49_, r_n_18__48_, r_n_18__47_, r_n_18__46_, r_n_18__45_, r_n_18__44_, r_n_18__43_, r_n_18__42_, r_n_18__41_, r_n_18__40_, r_n_18__39_, r_n_18__38_, r_n_18__37_, r_n_18__36_, r_n_18__35_, r_n_18__34_, r_n_18__33_, r_n_18__32_, r_n_18__31_, r_n_18__30_, r_n_18__29_, r_n_18__28_, r_n_18__27_, r_n_18__26_, r_n_18__25_, r_n_18__24_, r_n_18__23_, r_n_18__22_, r_n_18__21_, r_n_18__20_, r_n_18__19_, r_n_18__18_, r_n_18__17_, r_n_18__16_, r_n_18__15_, r_n_18__14_, r_n_18__13_, r_n_18__12_, r_n_18__11_, r_n_18__10_, r_n_18__9_, r_n_18__8_, r_n_18__7_, r_n_18__6_, r_n_18__5_, r_n_18__4_, r_n_18__3_, r_n_18__2_, r_n_18__1_, r_n_18__0_ } = (N36)? { r_19__63_, r_19__62_, r_19__61_, r_19__60_, r_19__59_, r_19__58_, r_19__57_, r_19__56_, r_19__55_, r_19__54_, r_19__53_, r_19__52_, r_19__51_, r_19__50_, r_19__49_, r_19__48_, r_19__47_, r_19__46_, r_19__45_, r_19__44_, r_19__43_, r_19__42_, r_19__41_, r_19__40_, r_19__39_, r_19__38_, r_19__37_, r_19__36_, r_19__35_, r_19__34_, r_19__33_, r_19__32_, r_19__31_, r_19__30_, r_19__29_, r_19__28_, r_19__27_, r_19__26_, r_19__25_, r_19__24_, r_19__23_, r_19__22_, r_19__21_, r_19__20_, r_19__19_, r_19__18_, r_19__17_, r_19__16_, r_19__15_, r_19__14_, r_19__13_, r_19__12_, r_19__11_, r_19__10_, r_19__9_, r_19__8_, r_19__7_, r_19__6_, r_19__5_, r_19__4_, r_19__3_, r_19__2_, r_19__1_, r_19__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N37)? data_i : 1'b0;
  assign N36 = sel_i[36];
  assign N37 = N1118;
  assign { r_n_19__63_, r_n_19__62_, r_n_19__61_, r_n_19__60_, r_n_19__59_, r_n_19__58_, r_n_19__57_, r_n_19__56_, r_n_19__55_, r_n_19__54_, r_n_19__53_, r_n_19__52_, r_n_19__51_, r_n_19__50_, r_n_19__49_, r_n_19__48_, r_n_19__47_, r_n_19__46_, r_n_19__45_, r_n_19__44_, r_n_19__43_, r_n_19__42_, r_n_19__41_, r_n_19__40_, r_n_19__39_, r_n_19__38_, r_n_19__37_, r_n_19__36_, r_n_19__35_, r_n_19__34_, r_n_19__33_, r_n_19__32_, r_n_19__31_, r_n_19__30_, r_n_19__29_, r_n_19__28_, r_n_19__27_, r_n_19__26_, r_n_19__25_, r_n_19__24_, r_n_19__23_, r_n_19__22_, r_n_19__21_, r_n_19__20_, r_n_19__19_, r_n_19__18_, r_n_19__17_, r_n_19__16_, r_n_19__15_, r_n_19__14_, r_n_19__13_, r_n_19__12_, r_n_19__11_, r_n_19__10_, r_n_19__9_, r_n_19__8_, r_n_19__7_, r_n_19__6_, r_n_19__5_, r_n_19__4_, r_n_19__3_, r_n_19__2_, r_n_19__1_, r_n_19__0_ } = (N38)? { r_20__63_, r_20__62_, r_20__61_, r_20__60_, r_20__59_, r_20__58_, r_20__57_, r_20__56_, r_20__55_, r_20__54_, r_20__53_, r_20__52_, r_20__51_, r_20__50_, r_20__49_, r_20__48_, r_20__47_, r_20__46_, r_20__45_, r_20__44_, r_20__43_, r_20__42_, r_20__41_, r_20__40_, r_20__39_, r_20__38_, r_20__37_, r_20__36_, r_20__35_, r_20__34_, r_20__33_, r_20__32_, r_20__31_, r_20__30_, r_20__29_, r_20__28_, r_20__27_, r_20__26_, r_20__25_, r_20__24_, r_20__23_, r_20__22_, r_20__21_, r_20__20_, r_20__19_, r_20__18_, r_20__17_, r_20__16_, r_20__15_, r_20__14_, r_20__13_, r_20__12_, r_20__11_, r_20__10_, r_20__9_, r_20__8_, r_20__7_, r_20__6_, r_20__5_, r_20__4_, r_20__3_, r_20__2_, r_20__1_, r_20__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N39)? data_i : 1'b0;
  assign N38 = sel_i[38];
  assign N39 = N1123;
  assign { r_n_20__63_, r_n_20__62_, r_n_20__61_, r_n_20__60_, r_n_20__59_, r_n_20__58_, r_n_20__57_, r_n_20__56_, r_n_20__55_, r_n_20__54_, r_n_20__53_, r_n_20__52_, r_n_20__51_, r_n_20__50_, r_n_20__49_, r_n_20__48_, r_n_20__47_, r_n_20__46_, r_n_20__45_, r_n_20__44_, r_n_20__43_, r_n_20__42_, r_n_20__41_, r_n_20__40_, r_n_20__39_, r_n_20__38_, r_n_20__37_, r_n_20__36_, r_n_20__35_, r_n_20__34_, r_n_20__33_, r_n_20__32_, r_n_20__31_, r_n_20__30_, r_n_20__29_, r_n_20__28_, r_n_20__27_, r_n_20__26_, r_n_20__25_, r_n_20__24_, r_n_20__23_, r_n_20__22_, r_n_20__21_, r_n_20__20_, r_n_20__19_, r_n_20__18_, r_n_20__17_, r_n_20__16_, r_n_20__15_, r_n_20__14_, r_n_20__13_, r_n_20__12_, r_n_20__11_, r_n_20__10_, r_n_20__9_, r_n_20__8_, r_n_20__7_, r_n_20__6_, r_n_20__5_, r_n_20__4_, r_n_20__3_, r_n_20__2_, r_n_20__1_, r_n_20__0_ } = (N40)? { r_21__63_, r_21__62_, r_21__61_, r_21__60_, r_21__59_, r_21__58_, r_21__57_, r_21__56_, r_21__55_, r_21__54_, r_21__53_, r_21__52_, r_21__51_, r_21__50_, r_21__49_, r_21__48_, r_21__47_, r_21__46_, r_21__45_, r_21__44_, r_21__43_, r_21__42_, r_21__41_, r_21__40_, r_21__39_, r_21__38_, r_21__37_, r_21__36_, r_21__35_, r_21__34_, r_21__33_, r_21__32_, r_21__31_, r_21__30_, r_21__29_, r_21__28_, r_21__27_, r_21__26_, r_21__25_, r_21__24_, r_21__23_, r_21__22_, r_21__21_, r_21__20_, r_21__19_, r_21__18_, r_21__17_, r_21__16_, r_21__15_, r_21__14_, r_21__13_, r_21__12_, r_21__11_, r_21__10_, r_21__9_, r_21__8_, r_21__7_, r_21__6_, r_21__5_, r_21__4_, r_21__3_, r_21__2_, r_21__1_, r_21__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N41)? data_i : 1'b0;
  assign N40 = sel_i[40];
  assign N41 = N1128;
  assign { r_n_21__63_, r_n_21__62_, r_n_21__61_, r_n_21__60_, r_n_21__59_, r_n_21__58_, r_n_21__57_, r_n_21__56_, r_n_21__55_, r_n_21__54_, r_n_21__53_, r_n_21__52_, r_n_21__51_, r_n_21__50_, r_n_21__49_, r_n_21__48_, r_n_21__47_, r_n_21__46_, r_n_21__45_, r_n_21__44_, r_n_21__43_, r_n_21__42_, r_n_21__41_, r_n_21__40_, r_n_21__39_, r_n_21__38_, r_n_21__37_, r_n_21__36_, r_n_21__35_, r_n_21__34_, r_n_21__33_, r_n_21__32_, r_n_21__31_, r_n_21__30_, r_n_21__29_, r_n_21__28_, r_n_21__27_, r_n_21__26_, r_n_21__25_, r_n_21__24_, r_n_21__23_, r_n_21__22_, r_n_21__21_, r_n_21__20_, r_n_21__19_, r_n_21__18_, r_n_21__17_, r_n_21__16_, r_n_21__15_, r_n_21__14_, r_n_21__13_, r_n_21__12_, r_n_21__11_, r_n_21__10_, r_n_21__9_, r_n_21__8_, r_n_21__7_, r_n_21__6_, r_n_21__5_, r_n_21__4_, r_n_21__3_, r_n_21__2_, r_n_21__1_, r_n_21__0_ } = (N42)? { r_22__63_, r_22__62_, r_22__61_, r_22__60_, r_22__59_, r_22__58_, r_22__57_, r_22__56_, r_22__55_, r_22__54_, r_22__53_, r_22__52_, r_22__51_, r_22__50_, r_22__49_, r_22__48_, r_22__47_, r_22__46_, r_22__45_, r_22__44_, r_22__43_, r_22__42_, r_22__41_, r_22__40_, r_22__39_, r_22__38_, r_22__37_, r_22__36_, r_22__35_, r_22__34_, r_22__33_, r_22__32_, r_22__31_, r_22__30_, r_22__29_, r_22__28_, r_22__27_, r_22__26_, r_22__25_, r_22__24_, r_22__23_, r_22__22_, r_22__21_, r_22__20_, r_22__19_, r_22__18_, r_22__17_, r_22__16_, r_22__15_, r_22__14_, r_22__13_, r_22__12_, r_22__11_, r_22__10_, r_22__9_, r_22__8_, r_22__7_, r_22__6_, r_22__5_, r_22__4_, r_22__3_, r_22__2_, r_22__1_, r_22__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N43)? data_i : 1'b0;
  assign N42 = sel_i[42];
  assign N43 = N1133;
  assign { r_n_22__63_, r_n_22__62_, r_n_22__61_, r_n_22__60_, r_n_22__59_, r_n_22__58_, r_n_22__57_, r_n_22__56_, r_n_22__55_, r_n_22__54_, r_n_22__53_, r_n_22__52_, r_n_22__51_, r_n_22__50_, r_n_22__49_, r_n_22__48_, r_n_22__47_, r_n_22__46_, r_n_22__45_, r_n_22__44_, r_n_22__43_, r_n_22__42_, r_n_22__41_, r_n_22__40_, r_n_22__39_, r_n_22__38_, r_n_22__37_, r_n_22__36_, r_n_22__35_, r_n_22__34_, r_n_22__33_, r_n_22__32_, r_n_22__31_, r_n_22__30_, r_n_22__29_, r_n_22__28_, r_n_22__27_, r_n_22__26_, r_n_22__25_, r_n_22__24_, r_n_22__23_, r_n_22__22_, r_n_22__21_, r_n_22__20_, r_n_22__19_, r_n_22__18_, r_n_22__17_, r_n_22__16_, r_n_22__15_, r_n_22__14_, r_n_22__13_, r_n_22__12_, r_n_22__11_, r_n_22__10_, r_n_22__9_, r_n_22__8_, r_n_22__7_, r_n_22__6_, r_n_22__5_, r_n_22__4_, r_n_22__3_, r_n_22__2_, r_n_22__1_, r_n_22__0_ } = (N44)? { r_23__63_, r_23__62_, r_23__61_, r_23__60_, r_23__59_, r_23__58_, r_23__57_, r_23__56_, r_23__55_, r_23__54_, r_23__53_, r_23__52_, r_23__51_, r_23__50_, r_23__49_, r_23__48_, r_23__47_, r_23__46_, r_23__45_, r_23__44_, r_23__43_, r_23__42_, r_23__41_, r_23__40_, r_23__39_, r_23__38_, r_23__37_, r_23__36_, r_23__35_, r_23__34_, r_23__33_, r_23__32_, r_23__31_, r_23__30_, r_23__29_, r_23__28_, r_23__27_, r_23__26_, r_23__25_, r_23__24_, r_23__23_, r_23__22_, r_23__21_, r_23__20_, r_23__19_, r_23__18_, r_23__17_, r_23__16_, r_23__15_, r_23__14_, r_23__13_, r_23__12_, r_23__11_, r_23__10_, r_23__9_, r_23__8_, r_23__7_, r_23__6_, r_23__5_, r_23__4_, r_23__3_, r_23__2_, r_23__1_, r_23__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N45)? data_i : 1'b0;
  assign N44 = sel_i[44];
  assign N45 = N1138;
  assign { r_n_23__63_, r_n_23__62_, r_n_23__61_, r_n_23__60_, r_n_23__59_, r_n_23__58_, r_n_23__57_, r_n_23__56_, r_n_23__55_, r_n_23__54_, r_n_23__53_, r_n_23__52_, r_n_23__51_, r_n_23__50_, r_n_23__49_, r_n_23__48_, r_n_23__47_, r_n_23__46_, r_n_23__45_, r_n_23__44_, r_n_23__43_, r_n_23__42_, r_n_23__41_, r_n_23__40_, r_n_23__39_, r_n_23__38_, r_n_23__37_, r_n_23__36_, r_n_23__35_, r_n_23__34_, r_n_23__33_, r_n_23__32_, r_n_23__31_, r_n_23__30_, r_n_23__29_, r_n_23__28_, r_n_23__27_, r_n_23__26_, r_n_23__25_, r_n_23__24_, r_n_23__23_, r_n_23__22_, r_n_23__21_, r_n_23__20_, r_n_23__19_, r_n_23__18_, r_n_23__17_, r_n_23__16_, r_n_23__15_, r_n_23__14_, r_n_23__13_, r_n_23__12_, r_n_23__11_, r_n_23__10_, r_n_23__9_, r_n_23__8_, r_n_23__7_, r_n_23__6_, r_n_23__5_, r_n_23__4_, r_n_23__3_, r_n_23__2_, r_n_23__1_, r_n_23__0_ } = (N46)? { r_24__63_, r_24__62_, r_24__61_, r_24__60_, r_24__59_, r_24__58_, r_24__57_, r_24__56_, r_24__55_, r_24__54_, r_24__53_, r_24__52_, r_24__51_, r_24__50_, r_24__49_, r_24__48_, r_24__47_, r_24__46_, r_24__45_, r_24__44_, r_24__43_, r_24__42_, r_24__41_, r_24__40_, r_24__39_, r_24__38_, r_24__37_, r_24__36_, r_24__35_, r_24__34_, r_24__33_, r_24__32_, r_24__31_, r_24__30_, r_24__29_, r_24__28_, r_24__27_, r_24__26_, r_24__25_, r_24__24_, r_24__23_, r_24__22_, r_24__21_, r_24__20_, r_24__19_, r_24__18_, r_24__17_, r_24__16_, r_24__15_, r_24__14_, r_24__13_, r_24__12_, r_24__11_, r_24__10_, r_24__9_, r_24__8_, r_24__7_, r_24__6_, r_24__5_, r_24__4_, r_24__3_, r_24__2_, r_24__1_, r_24__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N47)? data_i : 1'b0;
  assign N46 = sel_i[46];
  assign N47 = N1143;
  assign { r_n_24__63_, r_n_24__62_, r_n_24__61_, r_n_24__60_, r_n_24__59_, r_n_24__58_, r_n_24__57_, r_n_24__56_, r_n_24__55_, r_n_24__54_, r_n_24__53_, r_n_24__52_, r_n_24__51_, r_n_24__50_, r_n_24__49_, r_n_24__48_, r_n_24__47_, r_n_24__46_, r_n_24__45_, r_n_24__44_, r_n_24__43_, r_n_24__42_, r_n_24__41_, r_n_24__40_, r_n_24__39_, r_n_24__38_, r_n_24__37_, r_n_24__36_, r_n_24__35_, r_n_24__34_, r_n_24__33_, r_n_24__32_, r_n_24__31_, r_n_24__30_, r_n_24__29_, r_n_24__28_, r_n_24__27_, r_n_24__26_, r_n_24__25_, r_n_24__24_, r_n_24__23_, r_n_24__22_, r_n_24__21_, r_n_24__20_, r_n_24__19_, r_n_24__18_, r_n_24__17_, r_n_24__16_, r_n_24__15_, r_n_24__14_, r_n_24__13_, r_n_24__12_, r_n_24__11_, r_n_24__10_, r_n_24__9_, r_n_24__8_, r_n_24__7_, r_n_24__6_, r_n_24__5_, r_n_24__4_, r_n_24__3_, r_n_24__2_, r_n_24__1_, r_n_24__0_ } = (N48)? { r_25__63_, r_25__62_, r_25__61_, r_25__60_, r_25__59_, r_25__58_, r_25__57_, r_25__56_, r_25__55_, r_25__54_, r_25__53_, r_25__52_, r_25__51_, r_25__50_, r_25__49_, r_25__48_, r_25__47_, r_25__46_, r_25__45_, r_25__44_, r_25__43_, r_25__42_, r_25__41_, r_25__40_, r_25__39_, r_25__38_, r_25__37_, r_25__36_, r_25__35_, r_25__34_, r_25__33_, r_25__32_, r_25__31_, r_25__30_, r_25__29_, r_25__28_, r_25__27_, r_25__26_, r_25__25_, r_25__24_, r_25__23_, r_25__22_, r_25__21_, r_25__20_, r_25__19_, r_25__18_, r_25__17_, r_25__16_, r_25__15_, r_25__14_, r_25__13_, r_25__12_, r_25__11_, r_25__10_, r_25__9_, r_25__8_, r_25__7_, r_25__6_, r_25__5_, r_25__4_, r_25__3_, r_25__2_, r_25__1_, r_25__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N49)? data_i : 1'b0;
  assign N48 = sel_i[48];
  assign N49 = N1148;
  assign { r_n_25__63_, r_n_25__62_, r_n_25__61_, r_n_25__60_, r_n_25__59_, r_n_25__58_, r_n_25__57_, r_n_25__56_, r_n_25__55_, r_n_25__54_, r_n_25__53_, r_n_25__52_, r_n_25__51_, r_n_25__50_, r_n_25__49_, r_n_25__48_, r_n_25__47_, r_n_25__46_, r_n_25__45_, r_n_25__44_, r_n_25__43_, r_n_25__42_, r_n_25__41_, r_n_25__40_, r_n_25__39_, r_n_25__38_, r_n_25__37_, r_n_25__36_, r_n_25__35_, r_n_25__34_, r_n_25__33_, r_n_25__32_, r_n_25__31_, r_n_25__30_, r_n_25__29_, r_n_25__28_, r_n_25__27_, r_n_25__26_, r_n_25__25_, r_n_25__24_, r_n_25__23_, r_n_25__22_, r_n_25__21_, r_n_25__20_, r_n_25__19_, r_n_25__18_, r_n_25__17_, r_n_25__16_, r_n_25__15_, r_n_25__14_, r_n_25__13_, r_n_25__12_, r_n_25__11_, r_n_25__10_, r_n_25__9_, r_n_25__8_, r_n_25__7_, r_n_25__6_, r_n_25__5_, r_n_25__4_, r_n_25__3_, r_n_25__2_, r_n_25__1_, r_n_25__0_ } = (N50)? { r_26__63_, r_26__62_, r_26__61_, r_26__60_, r_26__59_, r_26__58_, r_26__57_, r_26__56_, r_26__55_, r_26__54_, r_26__53_, r_26__52_, r_26__51_, r_26__50_, r_26__49_, r_26__48_, r_26__47_, r_26__46_, r_26__45_, r_26__44_, r_26__43_, r_26__42_, r_26__41_, r_26__40_, r_26__39_, r_26__38_, r_26__37_, r_26__36_, r_26__35_, r_26__34_, r_26__33_, r_26__32_, r_26__31_, r_26__30_, r_26__29_, r_26__28_, r_26__27_, r_26__26_, r_26__25_, r_26__24_, r_26__23_, r_26__22_, r_26__21_, r_26__20_, r_26__19_, r_26__18_, r_26__17_, r_26__16_, r_26__15_, r_26__14_, r_26__13_, r_26__12_, r_26__11_, r_26__10_, r_26__9_, r_26__8_, r_26__7_, r_26__6_, r_26__5_, r_26__4_, r_26__3_, r_26__2_, r_26__1_, r_26__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N51)? data_i : 1'b0;
  assign N50 = sel_i[50];
  assign N51 = N1153;
  assign { r_n_26__63_, r_n_26__62_, r_n_26__61_, r_n_26__60_, r_n_26__59_, r_n_26__58_, r_n_26__57_, r_n_26__56_, r_n_26__55_, r_n_26__54_, r_n_26__53_, r_n_26__52_, r_n_26__51_, r_n_26__50_, r_n_26__49_, r_n_26__48_, r_n_26__47_, r_n_26__46_, r_n_26__45_, r_n_26__44_, r_n_26__43_, r_n_26__42_, r_n_26__41_, r_n_26__40_, r_n_26__39_, r_n_26__38_, r_n_26__37_, r_n_26__36_, r_n_26__35_, r_n_26__34_, r_n_26__33_, r_n_26__32_, r_n_26__31_, r_n_26__30_, r_n_26__29_, r_n_26__28_, r_n_26__27_, r_n_26__26_, r_n_26__25_, r_n_26__24_, r_n_26__23_, r_n_26__22_, r_n_26__21_, r_n_26__20_, r_n_26__19_, r_n_26__18_, r_n_26__17_, r_n_26__16_, r_n_26__15_, r_n_26__14_, r_n_26__13_, r_n_26__12_, r_n_26__11_, r_n_26__10_, r_n_26__9_, r_n_26__8_, r_n_26__7_, r_n_26__6_, r_n_26__5_, r_n_26__4_, r_n_26__3_, r_n_26__2_, r_n_26__1_, r_n_26__0_ } = (N52)? { r_27__63_, r_27__62_, r_27__61_, r_27__60_, r_27__59_, r_27__58_, r_27__57_, r_27__56_, r_27__55_, r_27__54_, r_27__53_, r_27__52_, r_27__51_, r_27__50_, r_27__49_, r_27__48_, r_27__47_, r_27__46_, r_27__45_, r_27__44_, r_27__43_, r_27__42_, r_27__41_, r_27__40_, r_27__39_, r_27__38_, r_27__37_, r_27__36_, r_27__35_, r_27__34_, r_27__33_, r_27__32_, r_27__31_, r_27__30_, r_27__29_, r_27__28_, r_27__27_, r_27__26_, r_27__25_, r_27__24_, r_27__23_, r_27__22_, r_27__21_, r_27__20_, r_27__19_, r_27__18_, r_27__17_, r_27__16_, r_27__15_, r_27__14_, r_27__13_, r_27__12_, r_27__11_, r_27__10_, r_27__9_, r_27__8_, r_27__7_, r_27__6_, r_27__5_, r_27__4_, r_27__3_, r_27__2_, r_27__1_, r_27__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N53)? data_i : 1'b0;
  assign N52 = sel_i[52];
  assign N53 = N1158;
  assign { r_n_27__63_, r_n_27__62_, r_n_27__61_, r_n_27__60_, r_n_27__59_, r_n_27__58_, r_n_27__57_, r_n_27__56_, r_n_27__55_, r_n_27__54_, r_n_27__53_, r_n_27__52_, r_n_27__51_, r_n_27__50_, r_n_27__49_, r_n_27__48_, r_n_27__47_, r_n_27__46_, r_n_27__45_, r_n_27__44_, r_n_27__43_, r_n_27__42_, r_n_27__41_, r_n_27__40_, r_n_27__39_, r_n_27__38_, r_n_27__37_, r_n_27__36_, r_n_27__35_, r_n_27__34_, r_n_27__33_, r_n_27__32_, r_n_27__31_, r_n_27__30_, r_n_27__29_, r_n_27__28_, r_n_27__27_, r_n_27__26_, r_n_27__25_, r_n_27__24_, r_n_27__23_, r_n_27__22_, r_n_27__21_, r_n_27__20_, r_n_27__19_, r_n_27__18_, r_n_27__17_, r_n_27__16_, r_n_27__15_, r_n_27__14_, r_n_27__13_, r_n_27__12_, r_n_27__11_, r_n_27__10_, r_n_27__9_, r_n_27__8_, r_n_27__7_, r_n_27__6_, r_n_27__5_, r_n_27__4_, r_n_27__3_, r_n_27__2_, r_n_27__1_, r_n_27__0_ } = (N54)? { r_28__63_, r_28__62_, r_28__61_, r_28__60_, r_28__59_, r_28__58_, r_28__57_, r_28__56_, r_28__55_, r_28__54_, r_28__53_, r_28__52_, r_28__51_, r_28__50_, r_28__49_, r_28__48_, r_28__47_, r_28__46_, r_28__45_, r_28__44_, r_28__43_, r_28__42_, r_28__41_, r_28__40_, r_28__39_, r_28__38_, r_28__37_, r_28__36_, r_28__35_, r_28__34_, r_28__33_, r_28__32_, r_28__31_, r_28__30_, r_28__29_, r_28__28_, r_28__27_, r_28__26_, r_28__25_, r_28__24_, r_28__23_, r_28__22_, r_28__21_, r_28__20_, r_28__19_, r_28__18_, r_28__17_, r_28__16_, r_28__15_, r_28__14_, r_28__13_, r_28__12_, r_28__11_, r_28__10_, r_28__9_, r_28__8_, r_28__7_, r_28__6_, r_28__5_, r_28__4_, r_28__3_, r_28__2_, r_28__1_, r_28__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N55)? data_i : 1'b0;
  assign N54 = sel_i[54];
  assign N55 = N1163;
  assign { r_n_28__63_, r_n_28__62_, r_n_28__61_, r_n_28__60_, r_n_28__59_, r_n_28__58_, r_n_28__57_, r_n_28__56_, r_n_28__55_, r_n_28__54_, r_n_28__53_, r_n_28__52_, r_n_28__51_, r_n_28__50_, r_n_28__49_, r_n_28__48_, r_n_28__47_, r_n_28__46_, r_n_28__45_, r_n_28__44_, r_n_28__43_, r_n_28__42_, r_n_28__41_, r_n_28__40_, r_n_28__39_, r_n_28__38_, r_n_28__37_, r_n_28__36_, r_n_28__35_, r_n_28__34_, r_n_28__33_, r_n_28__32_, r_n_28__31_, r_n_28__30_, r_n_28__29_, r_n_28__28_, r_n_28__27_, r_n_28__26_, r_n_28__25_, r_n_28__24_, r_n_28__23_, r_n_28__22_, r_n_28__21_, r_n_28__20_, r_n_28__19_, r_n_28__18_, r_n_28__17_, r_n_28__16_, r_n_28__15_, r_n_28__14_, r_n_28__13_, r_n_28__12_, r_n_28__11_, r_n_28__10_, r_n_28__9_, r_n_28__8_, r_n_28__7_, r_n_28__6_, r_n_28__5_, r_n_28__4_, r_n_28__3_, r_n_28__2_, r_n_28__1_, r_n_28__0_ } = (N56)? { r_29__63_, r_29__62_, r_29__61_, r_29__60_, r_29__59_, r_29__58_, r_29__57_, r_29__56_, r_29__55_, r_29__54_, r_29__53_, r_29__52_, r_29__51_, r_29__50_, r_29__49_, r_29__48_, r_29__47_, r_29__46_, r_29__45_, r_29__44_, r_29__43_, r_29__42_, r_29__41_, r_29__40_, r_29__39_, r_29__38_, r_29__37_, r_29__36_, r_29__35_, r_29__34_, r_29__33_, r_29__32_, r_29__31_, r_29__30_, r_29__29_, r_29__28_, r_29__27_, r_29__26_, r_29__25_, r_29__24_, r_29__23_, r_29__22_, r_29__21_, r_29__20_, r_29__19_, r_29__18_, r_29__17_, r_29__16_, r_29__15_, r_29__14_, r_29__13_, r_29__12_, r_29__11_, r_29__10_, r_29__9_, r_29__8_, r_29__7_, r_29__6_, r_29__5_, r_29__4_, r_29__3_, r_29__2_, r_29__1_, r_29__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N57)? data_i : 1'b0;
  assign N56 = sel_i[56];
  assign N57 = N1168;
  assign { r_n_29__63_, r_n_29__62_, r_n_29__61_, r_n_29__60_, r_n_29__59_, r_n_29__58_, r_n_29__57_, r_n_29__56_, r_n_29__55_, r_n_29__54_, r_n_29__53_, r_n_29__52_, r_n_29__51_, r_n_29__50_, r_n_29__49_, r_n_29__48_, r_n_29__47_, r_n_29__46_, r_n_29__45_, r_n_29__44_, r_n_29__43_, r_n_29__42_, r_n_29__41_, r_n_29__40_, r_n_29__39_, r_n_29__38_, r_n_29__37_, r_n_29__36_, r_n_29__35_, r_n_29__34_, r_n_29__33_, r_n_29__32_, r_n_29__31_, r_n_29__30_, r_n_29__29_, r_n_29__28_, r_n_29__27_, r_n_29__26_, r_n_29__25_, r_n_29__24_, r_n_29__23_, r_n_29__22_, r_n_29__21_, r_n_29__20_, r_n_29__19_, r_n_29__18_, r_n_29__17_, r_n_29__16_, r_n_29__15_, r_n_29__14_, r_n_29__13_, r_n_29__12_, r_n_29__11_, r_n_29__10_, r_n_29__9_, r_n_29__8_, r_n_29__7_, r_n_29__6_, r_n_29__5_, r_n_29__4_, r_n_29__3_, r_n_29__2_, r_n_29__1_, r_n_29__0_ } = (N58)? { r_30__63_, r_30__62_, r_30__61_, r_30__60_, r_30__59_, r_30__58_, r_30__57_, r_30__56_, r_30__55_, r_30__54_, r_30__53_, r_30__52_, r_30__51_, r_30__50_, r_30__49_, r_30__48_, r_30__47_, r_30__46_, r_30__45_, r_30__44_, r_30__43_, r_30__42_, r_30__41_, r_30__40_, r_30__39_, r_30__38_, r_30__37_, r_30__36_, r_30__35_, r_30__34_, r_30__33_, r_30__32_, r_30__31_, r_30__30_, r_30__29_, r_30__28_, r_30__27_, r_30__26_, r_30__25_, r_30__24_, r_30__23_, r_30__22_, r_30__21_, r_30__20_, r_30__19_, r_30__18_, r_30__17_, r_30__16_, r_30__15_, r_30__14_, r_30__13_, r_30__12_, r_30__11_, r_30__10_, r_30__9_, r_30__8_, r_30__7_, r_30__6_, r_30__5_, r_30__4_, r_30__3_, r_30__2_, r_30__1_, r_30__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N59)? data_i : 1'b0;
  assign N58 = sel_i[58];
  assign N59 = N1173;
  assign { r_n_30__63_, r_n_30__62_, r_n_30__61_, r_n_30__60_, r_n_30__59_, r_n_30__58_, r_n_30__57_, r_n_30__56_, r_n_30__55_, r_n_30__54_, r_n_30__53_, r_n_30__52_, r_n_30__51_, r_n_30__50_, r_n_30__49_, r_n_30__48_, r_n_30__47_, r_n_30__46_, r_n_30__45_, r_n_30__44_, r_n_30__43_, r_n_30__42_, r_n_30__41_, r_n_30__40_, r_n_30__39_, r_n_30__38_, r_n_30__37_, r_n_30__36_, r_n_30__35_, r_n_30__34_, r_n_30__33_, r_n_30__32_, r_n_30__31_, r_n_30__30_, r_n_30__29_, r_n_30__28_, r_n_30__27_, r_n_30__26_, r_n_30__25_, r_n_30__24_, r_n_30__23_, r_n_30__22_, r_n_30__21_, r_n_30__20_, r_n_30__19_, r_n_30__18_, r_n_30__17_, r_n_30__16_, r_n_30__15_, r_n_30__14_, r_n_30__13_, r_n_30__12_, r_n_30__11_, r_n_30__10_, r_n_30__9_, r_n_30__8_, r_n_30__7_, r_n_30__6_, r_n_30__5_, r_n_30__4_, r_n_30__3_, r_n_30__2_, r_n_30__1_, r_n_30__0_ } = (N60)? { r_31__63_, r_31__62_, r_31__61_, r_31__60_, r_31__59_, r_31__58_, r_31__57_, r_31__56_, r_31__55_, r_31__54_, r_31__53_, r_31__52_, r_31__51_, r_31__50_, r_31__49_, r_31__48_, r_31__47_, r_31__46_, r_31__45_, r_31__44_, r_31__43_, r_31__42_, r_31__41_, r_31__40_, r_31__39_, r_31__38_, r_31__37_, r_31__36_, r_31__35_, r_31__34_, r_31__33_, r_31__32_, r_31__31_, r_31__30_, r_31__29_, r_31__28_, r_31__27_, r_31__26_, r_31__25_, r_31__24_, r_31__23_, r_31__22_, r_31__21_, r_31__20_, r_31__19_, r_31__18_, r_31__17_, r_31__16_, r_31__15_, r_31__14_, r_31__13_, r_31__12_, r_31__11_, r_31__10_, r_31__9_, r_31__8_, r_31__7_, r_31__6_, r_31__5_, r_31__4_, r_31__3_, r_31__2_, r_31__1_, r_31__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N61)? data_i : 1'b0;
  assign N60 = sel_i[60];
  assign N61 = N1178;
  assign { r_n_31__63_, r_n_31__62_, r_n_31__61_, r_n_31__60_, r_n_31__59_, r_n_31__58_, r_n_31__57_, r_n_31__56_, r_n_31__55_, r_n_31__54_, r_n_31__53_, r_n_31__52_, r_n_31__51_, r_n_31__50_, r_n_31__49_, r_n_31__48_, r_n_31__47_, r_n_31__46_, r_n_31__45_, r_n_31__44_, r_n_31__43_, r_n_31__42_, r_n_31__41_, r_n_31__40_, r_n_31__39_, r_n_31__38_, r_n_31__37_, r_n_31__36_, r_n_31__35_, r_n_31__34_, r_n_31__33_, r_n_31__32_, r_n_31__31_, r_n_31__30_, r_n_31__29_, r_n_31__28_, r_n_31__27_, r_n_31__26_, r_n_31__25_, r_n_31__24_, r_n_31__23_, r_n_31__22_, r_n_31__21_, r_n_31__20_, r_n_31__19_, r_n_31__18_, r_n_31__17_, r_n_31__16_, r_n_31__15_, r_n_31__14_, r_n_31__13_, r_n_31__12_, r_n_31__11_, r_n_31__10_, r_n_31__9_, r_n_31__8_, r_n_31__7_, r_n_31__6_, r_n_31__5_, r_n_31__4_, r_n_31__3_, r_n_31__2_, r_n_31__1_, r_n_31__0_ } = (N62)? { r_32__63_, r_32__62_, r_32__61_, r_32__60_, r_32__59_, r_32__58_, r_32__57_, r_32__56_, r_32__55_, r_32__54_, r_32__53_, r_32__52_, r_32__51_, r_32__50_, r_32__49_, r_32__48_, r_32__47_, r_32__46_, r_32__45_, r_32__44_, r_32__43_, r_32__42_, r_32__41_, r_32__40_, r_32__39_, r_32__38_, r_32__37_, r_32__36_, r_32__35_, r_32__34_, r_32__33_, r_32__32_, r_32__31_, r_32__30_, r_32__29_, r_32__28_, r_32__27_, r_32__26_, r_32__25_, r_32__24_, r_32__23_, r_32__22_, r_32__21_, r_32__20_, r_32__19_, r_32__18_, r_32__17_, r_32__16_, r_32__15_, r_32__14_, r_32__13_, r_32__12_, r_32__11_, r_32__10_, r_32__9_, r_32__8_, r_32__7_, r_32__6_, r_32__5_, r_32__4_, r_32__3_, r_32__2_, r_32__1_, r_32__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N63)? data_i : 1'b0;
  assign N62 = sel_i[62];
  assign N63 = N1183;
  assign { r_n_32__63_, r_n_32__62_, r_n_32__61_, r_n_32__60_, r_n_32__59_, r_n_32__58_, r_n_32__57_, r_n_32__56_, r_n_32__55_, r_n_32__54_, r_n_32__53_, r_n_32__52_, r_n_32__51_, r_n_32__50_, r_n_32__49_, r_n_32__48_, r_n_32__47_, r_n_32__46_, r_n_32__45_, r_n_32__44_, r_n_32__43_, r_n_32__42_, r_n_32__41_, r_n_32__40_, r_n_32__39_, r_n_32__38_, r_n_32__37_, r_n_32__36_, r_n_32__35_, r_n_32__34_, r_n_32__33_, r_n_32__32_, r_n_32__31_, r_n_32__30_, r_n_32__29_, r_n_32__28_, r_n_32__27_, r_n_32__26_, r_n_32__25_, r_n_32__24_, r_n_32__23_, r_n_32__22_, r_n_32__21_, r_n_32__20_, r_n_32__19_, r_n_32__18_, r_n_32__17_, r_n_32__16_, r_n_32__15_, r_n_32__14_, r_n_32__13_, r_n_32__12_, r_n_32__11_, r_n_32__10_, r_n_32__9_, r_n_32__8_, r_n_32__7_, r_n_32__6_, r_n_32__5_, r_n_32__4_, r_n_32__3_, r_n_32__2_, r_n_32__1_, r_n_32__0_ } = (N64)? { r_33__63_, r_33__62_, r_33__61_, r_33__60_, r_33__59_, r_33__58_, r_33__57_, r_33__56_, r_33__55_, r_33__54_, r_33__53_, r_33__52_, r_33__51_, r_33__50_, r_33__49_, r_33__48_, r_33__47_, r_33__46_, r_33__45_, r_33__44_, r_33__43_, r_33__42_, r_33__41_, r_33__40_, r_33__39_, r_33__38_, r_33__37_, r_33__36_, r_33__35_, r_33__34_, r_33__33_, r_33__32_, r_33__31_, r_33__30_, r_33__29_, r_33__28_, r_33__27_, r_33__26_, r_33__25_, r_33__24_, r_33__23_, r_33__22_, r_33__21_, r_33__20_, r_33__19_, r_33__18_, r_33__17_, r_33__16_, r_33__15_, r_33__14_, r_33__13_, r_33__12_, r_33__11_, r_33__10_, r_33__9_, r_33__8_, r_33__7_, r_33__6_, r_33__5_, r_33__4_, r_33__3_, r_33__2_, r_33__1_, r_33__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N65)? data_i : 1'b0;
  assign N64 = sel_i[64];
  assign N65 = N1188;
  assign { r_n_33__63_, r_n_33__62_, r_n_33__61_, r_n_33__60_, r_n_33__59_, r_n_33__58_, r_n_33__57_, r_n_33__56_, r_n_33__55_, r_n_33__54_, r_n_33__53_, r_n_33__52_, r_n_33__51_, r_n_33__50_, r_n_33__49_, r_n_33__48_, r_n_33__47_, r_n_33__46_, r_n_33__45_, r_n_33__44_, r_n_33__43_, r_n_33__42_, r_n_33__41_, r_n_33__40_, r_n_33__39_, r_n_33__38_, r_n_33__37_, r_n_33__36_, r_n_33__35_, r_n_33__34_, r_n_33__33_, r_n_33__32_, r_n_33__31_, r_n_33__30_, r_n_33__29_, r_n_33__28_, r_n_33__27_, r_n_33__26_, r_n_33__25_, r_n_33__24_, r_n_33__23_, r_n_33__22_, r_n_33__21_, r_n_33__20_, r_n_33__19_, r_n_33__18_, r_n_33__17_, r_n_33__16_, r_n_33__15_, r_n_33__14_, r_n_33__13_, r_n_33__12_, r_n_33__11_, r_n_33__10_, r_n_33__9_, r_n_33__8_, r_n_33__7_, r_n_33__6_, r_n_33__5_, r_n_33__4_, r_n_33__3_, r_n_33__2_, r_n_33__1_, r_n_33__0_ } = (N66)? { r_34__63_, r_34__62_, r_34__61_, r_34__60_, r_34__59_, r_34__58_, r_34__57_, r_34__56_, r_34__55_, r_34__54_, r_34__53_, r_34__52_, r_34__51_, r_34__50_, r_34__49_, r_34__48_, r_34__47_, r_34__46_, r_34__45_, r_34__44_, r_34__43_, r_34__42_, r_34__41_, r_34__40_, r_34__39_, r_34__38_, r_34__37_, r_34__36_, r_34__35_, r_34__34_, r_34__33_, r_34__32_, r_34__31_, r_34__30_, r_34__29_, r_34__28_, r_34__27_, r_34__26_, r_34__25_, r_34__24_, r_34__23_, r_34__22_, r_34__21_, r_34__20_, r_34__19_, r_34__18_, r_34__17_, r_34__16_, r_34__15_, r_34__14_, r_34__13_, r_34__12_, r_34__11_, r_34__10_, r_34__9_, r_34__8_, r_34__7_, r_34__6_, r_34__5_, r_34__4_, r_34__3_, r_34__2_, r_34__1_, r_34__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N67)? data_i : 1'b0;
  assign N66 = sel_i[66];
  assign N67 = N1193;
  assign { r_n_34__63_, r_n_34__62_, r_n_34__61_, r_n_34__60_, r_n_34__59_, r_n_34__58_, r_n_34__57_, r_n_34__56_, r_n_34__55_, r_n_34__54_, r_n_34__53_, r_n_34__52_, r_n_34__51_, r_n_34__50_, r_n_34__49_, r_n_34__48_, r_n_34__47_, r_n_34__46_, r_n_34__45_, r_n_34__44_, r_n_34__43_, r_n_34__42_, r_n_34__41_, r_n_34__40_, r_n_34__39_, r_n_34__38_, r_n_34__37_, r_n_34__36_, r_n_34__35_, r_n_34__34_, r_n_34__33_, r_n_34__32_, r_n_34__31_, r_n_34__30_, r_n_34__29_, r_n_34__28_, r_n_34__27_, r_n_34__26_, r_n_34__25_, r_n_34__24_, r_n_34__23_, r_n_34__22_, r_n_34__21_, r_n_34__20_, r_n_34__19_, r_n_34__18_, r_n_34__17_, r_n_34__16_, r_n_34__15_, r_n_34__14_, r_n_34__13_, r_n_34__12_, r_n_34__11_, r_n_34__10_, r_n_34__9_, r_n_34__8_, r_n_34__7_, r_n_34__6_, r_n_34__5_, r_n_34__4_, r_n_34__3_, r_n_34__2_, r_n_34__1_, r_n_34__0_ } = (N68)? { r_35__63_, r_35__62_, r_35__61_, r_35__60_, r_35__59_, r_35__58_, r_35__57_, r_35__56_, r_35__55_, r_35__54_, r_35__53_, r_35__52_, r_35__51_, r_35__50_, r_35__49_, r_35__48_, r_35__47_, r_35__46_, r_35__45_, r_35__44_, r_35__43_, r_35__42_, r_35__41_, r_35__40_, r_35__39_, r_35__38_, r_35__37_, r_35__36_, r_35__35_, r_35__34_, r_35__33_, r_35__32_, r_35__31_, r_35__30_, r_35__29_, r_35__28_, r_35__27_, r_35__26_, r_35__25_, r_35__24_, r_35__23_, r_35__22_, r_35__21_, r_35__20_, r_35__19_, r_35__18_, r_35__17_, r_35__16_, r_35__15_, r_35__14_, r_35__13_, r_35__12_, r_35__11_, r_35__10_, r_35__9_, r_35__8_, r_35__7_, r_35__6_, r_35__5_, r_35__4_, r_35__3_, r_35__2_, r_35__1_, r_35__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N69)? data_i : 1'b0;
  assign N68 = sel_i[68];
  assign N69 = N1198;
  assign { r_n_35__63_, r_n_35__62_, r_n_35__61_, r_n_35__60_, r_n_35__59_, r_n_35__58_, r_n_35__57_, r_n_35__56_, r_n_35__55_, r_n_35__54_, r_n_35__53_, r_n_35__52_, r_n_35__51_, r_n_35__50_, r_n_35__49_, r_n_35__48_, r_n_35__47_, r_n_35__46_, r_n_35__45_, r_n_35__44_, r_n_35__43_, r_n_35__42_, r_n_35__41_, r_n_35__40_, r_n_35__39_, r_n_35__38_, r_n_35__37_, r_n_35__36_, r_n_35__35_, r_n_35__34_, r_n_35__33_, r_n_35__32_, r_n_35__31_, r_n_35__30_, r_n_35__29_, r_n_35__28_, r_n_35__27_, r_n_35__26_, r_n_35__25_, r_n_35__24_, r_n_35__23_, r_n_35__22_, r_n_35__21_, r_n_35__20_, r_n_35__19_, r_n_35__18_, r_n_35__17_, r_n_35__16_, r_n_35__15_, r_n_35__14_, r_n_35__13_, r_n_35__12_, r_n_35__11_, r_n_35__10_, r_n_35__9_, r_n_35__8_, r_n_35__7_, r_n_35__6_, r_n_35__5_, r_n_35__4_, r_n_35__3_, r_n_35__2_, r_n_35__1_, r_n_35__0_ } = (N70)? { r_36__63_, r_36__62_, r_36__61_, r_36__60_, r_36__59_, r_36__58_, r_36__57_, r_36__56_, r_36__55_, r_36__54_, r_36__53_, r_36__52_, r_36__51_, r_36__50_, r_36__49_, r_36__48_, r_36__47_, r_36__46_, r_36__45_, r_36__44_, r_36__43_, r_36__42_, r_36__41_, r_36__40_, r_36__39_, r_36__38_, r_36__37_, r_36__36_, r_36__35_, r_36__34_, r_36__33_, r_36__32_, r_36__31_, r_36__30_, r_36__29_, r_36__28_, r_36__27_, r_36__26_, r_36__25_, r_36__24_, r_36__23_, r_36__22_, r_36__21_, r_36__20_, r_36__19_, r_36__18_, r_36__17_, r_36__16_, r_36__15_, r_36__14_, r_36__13_, r_36__12_, r_36__11_, r_36__10_, r_36__9_, r_36__8_, r_36__7_, r_36__6_, r_36__5_, r_36__4_, r_36__3_, r_36__2_, r_36__1_, r_36__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N71)? data_i : 1'b0;
  assign N70 = sel_i[70];
  assign N71 = N1203;
  assign { r_n_36__63_, r_n_36__62_, r_n_36__61_, r_n_36__60_, r_n_36__59_, r_n_36__58_, r_n_36__57_, r_n_36__56_, r_n_36__55_, r_n_36__54_, r_n_36__53_, r_n_36__52_, r_n_36__51_, r_n_36__50_, r_n_36__49_, r_n_36__48_, r_n_36__47_, r_n_36__46_, r_n_36__45_, r_n_36__44_, r_n_36__43_, r_n_36__42_, r_n_36__41_, r_n_36__40_, r_n_36__39_, r_n_36__38_, r_n_36__37_, r_n_36__36_, r_n_36__35_, r_n_36__34_, r_n_36__33_, r_n_36__32_, r_n_36__31_, r_n_36__30_, r_n_36__29_, r_n_36__28_, r_n_36__27_, r_n_36__26_, r_n_36__25_, r_n_36__24_, r_n_36__23_, r_n_36__22_, r_n_36__21_, r_n_36__20_, r_n_36__19_, r_n_36__18_, r_n_36__17_, r_n_36__16_, r_n_36__15_, r_n_36__14_, r_n_36__13_, r_n_36__12_, r_n_36__11_, r_n_36__10_, r_n_36__9_, r_n_36__8_, r_n_36__7_, r_n_36__6_, r_n_36__5_, r_n_36__4_, r_n_36__3_, r_n_36__2_, r_n_36__1_, r_n_36__0_ } = (N72)? { r_37__63_, r_37__62_, r_37__61_, r_37__60_, r_37__59_, r_37__58_, r_37__57_, r_37__56_, r_37__55_, r_37__54_, r_37__53_, r_37__52_, r_37__51_, r_37__50_, r_37__49_, r_37__48_, r_37__47_, r_37__46_, r_37__45_, r_37__44_, r_37__43_, r_37__42_, r_37__41_, r_37__40_, r_37__39_, r_37__38_, r_37__37_, r_37__36_, r_37__35_, r_37__34_, r_37__33_, r_37__32_, r_37__31_, r_37__30_, r_37__29_, r_37__28_, r_37__27_, r_37__26_, r_37__25_, r_37__24_, r_37__23_, r_37__22_, r_37__21_, r_37__20_, r_37__19_, r_37__18_, r_37__17_, r_37__16_, r_37__15_, r_37__14_, r_37__13_, r_37__12_, r_37__11_, r_37__10_, r_37__9_, r_37__8_, r_37__7_, r_37__6_, r_37__5_, r_37__4_, r_37__3_, r_37__2_, r_37__1_, r_37__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N73)? data_i : 1'b0;
  assign N72 = sel_i[72];
  assign N73 = N1208;
  assign { r_n_37__63_, r_n_37__62_, r_n_37__61_, r_n_37__60_, r_n_37__59_, r_n_37__58_, r_n_37__57_, r_n_37__56_, r_n_37__55_, r_n_37__54_, r_n_37__53_, r_n_37__52_, r_n_37__51_, r_n_37__50_, r_n_37__49_, r_n_37__48_, r_n_37__47_, r_n_37__46_, r_n_37__45_, r_n_37__44_, r_n_37__43_, r_n_37__42_, r_n_37__41_, r_n_37__40_, r_n_37__39_, r_n_37__38_, r_n_37__37_, r_n_37__36_, r_n_37__35_, r_n_37__34_, r_n_37__33_, r_n_37__32_, r_n_37__31_, r_n_37__30_, r_n_37__29_, r_n_37__28_, r_n_37__27_, r_n_37__26_, r_n_37__25_, r_n_37__24_, r_n_37__23_, r_n_37__22_, r_n_37__21_, r_n_37__20_, r_n_37__19_, r_n_37__18_, r_n_37__17_, r_n_37__16_, r_n_37__15_, r_n_37__14_, r_n_37__13_, r_n_37__12_, r_n_37__11_, r_n_37__10_, r_n_37__9_, r_n_37__8_, r_n_37__7_, r_n_37__6_, r_n_37__5_, r_n_37__4_, r_n_37__3_, r_n_37__2_, r_n_37__1_, r_n_37__0_ } = (N74)? { r_38__63_, r_38__62_, r_38__61_, r_38__60_, r_38__59_, r_38__58_, r_38__57_, r_38__56_, r_38__55_, r_38__54_, r_38__53_, r_38__52_, r_38__51_, r_38__50_, r_38__49_, r_38__48_, r_38__47_, r_38__46_, r_38__45_, r_38__44_, r_38__43_, r_38__42_, r_38__41_, r_38__40_, r_38__39_, r_38__38_, r_38__37_, r_38__36_, r_38__35_, r_38__34_, r_38__33_, r_38__32_, r_38__31_, r_38__30_, r_38__29_, r_38__28_, r_38__27_, r_38__26_, r_38__25_, r_38__24_, r_38__23_, r_38__22_, r_38__21_, r_38__20_, r_38__19_, r_38__18_, r_38__17_, r_38__16_, r_38__15_, r_38__14_, r_38__13_, r_38__12_, r_38__11_, r_38__10_, r_38__9_, r_38__8_, r_38__7_, r_38__6_, r_38__5_, r_38__4_, r_38__3_, r_38__2_, r_38__1_, r_38__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N75)? data_i : 1'b0;
  assign N74 = sel_i[74];
  assign N75 = N1213;
  assign { r_n_38__63_, r_n_38__62_, r_n_38__61_, r_n_38__60_, r_n_38__59_, r_n_38__58_, r_n_38__57_, r_n_38__56_, r_n_38__55_, r_n_38__54_, r_n_38__53_, r_n_38__52_, r_n_38__51_, r_n_38__50_, r_n_38__49_, r_n_38__48_, r_n_38__47_, r_n_38__46_, r_n_38__45_, r_n_38__44_, r_n_38__43_, r_n_38__42_, r_n_38__41_, r_n_38__40_, r_n_38__39_, r_n_38__38_, r_n_38__37_, r_n_38__36_, r_n_38__35_, r_n_38__34_, r_n_38__33_, r_n_38__32_, r_n_38__31_, r_n_38__30_, r_n_38__29_, r_n_38__28_, r_n_38__27_, r_n_38__26_, r_n_38__25_, r_n_38__24_, r_n_38__23_, r_n_38__22_, r_n_38__21_, r_n_38__20_, r_n_38__19_, r_n_38__18_, r_n_38__17_, r_n_38__16_, r_n_38__15_, r_n_38__14_, r_n_38__13_, r_n_38__12_, r_n_38__11_, r_n_38__10_, r_n_38__9_, r_n_38__8_, r_n_38__7_, r_n_38__6_, r_n_38__5_, r_n_38__4_, r_n_38__3_, r_n_38__2_, r_n_38__1_, r_n_38__0_ } = (N76)? { r_39__63_, r_39__62_, r_39__61_, r_39__60_, r_39__59_, r_39__58_, r_39__57_, r_39__56_, r_39__55_, r_39__54_, r_39__53_, r_39__52_, r_39__51_, r_39__50_, r_39__49_, r_39__48_, r_39__47_, r_39__46_, r_39__45_, r_39__44_, r_39__43_, r_39__42_, r_39__41_, r_39__40_, r_39__39_, r_39__38_, r_39__37_, r_39__36_, r_39__35_, r_39__34_, r_39__33_, r_39__32_, r_39__31_, r_39__30_, r_39__29_, r_39__28_, r_39__27_, r_39__26_, r_39__25_, r_39__24_, r_39__23_, r_39__22_, r_39__21_, r_39__20_, r_39__19_, r_39__18_, r_39__17_, r_39__16_, r_39__15_, r_39__14_, r_39__13_, r_39__12_, r_39__11_, r_39__10_, r_39__9_, r_39__8_, r_39__7_, r_39__6_, r_39__5_, r_39__4_, r_39__3_, r_39__2_, r_39__1_, r_39__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N77)? data_i : 1'b0;
  assign N76 = sel_i[76];
  assign N77 = N1218;
  assign { r_n_39__63_, r_n_39__62_, r_n_39__61_, r_n_39__60_, r_n_39__59_, r_n_39__58_, r_n_39__57_, r_n_39__56_, r_n_39__55_, r_n_39__54_, r_n_39__53_, r_n_39__52_, r_n_39__51_, r_n_39__50_, r_n_39__49_, r_n_39__48_, r_n_39__47_, r_n_39__46_, r_n_39__45_, r_n_39__44_, r_n_39__43_, r_n_39__42_, r_n_39__41_, r_n_39__40_, r_n_39__39_, r_n_39__38_, r_n_39__37_, r_n_39__36_, r_n_39__35_, r_n_39__34_, r_n_39__33_, r_n_39__32_, r_n_39__31_, r_n_39__30_, r_n_39__29_, r_n_39__28_, r_n_39__27_, r_n_39__26_, r_n_39__25_, r_n_39__24_, r_n_39__23_, r_n_39__22_, r_n_39__21_, r_n_39__20_, r_n_39__19_, r_n_39__18_, r_n_39__17_, r_n_39__16_, r_n_39__15_, r_n_39__14_, r_n_39__13_, r_n_39__12_, r_n_39__11_, r_n_39__10_, r_n_39__9_, r_n_39__8_, r_n_39__7_, r_n_39__6_, r_n_39__5_, r_n_39__4_, r_n_39__3_, r_n_39__2_, r_n_39__1_, r_n_39__0_ } = (N78)? { r_40__63_, r_40__62_, r_40__61_, r_40__60_, r_40__59_, r_40__58_, r_40__57_, r_40__56_, r_40__55_, r_40__54_, r_40__53_, r_40__52_, r_40__51_, r_40__50_, r_40__49_, r_40__48_, r_40__47_, r_40__46_, r_40__45_, r_40__44_, r_40__43_, r_40__42_, r_40__41_, r_40__40_, r_40__39_, r_40__38_, r_40__37_, r_40__36_, r_40__35_, r_40__34_, r_40__33_, r_40__32_, r_40__31_, r_40__30_, r_40__29_, r_40__28_, r_40__27_, r_40__26_, r_40__25_, r_40__24_, r_40__23_, r_40__22_, r_40__21_, r_40__20_, r_40__19_, r_40__18_, r_40__17_, r_40__16_, r_40__15_, r_40__14_, r_40__13_, r_40__12_, r_40__11_, r_40__10_, r_40__9_, r_40__8_, r_40__7_, r_40__6_, r_40__5_, r_40__4_, r_40__3_, r_40__2_, r_40__1_, r_40__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N79)? data_i : 1'b0;
  assign N78 = sel_i[78];
  assign N79 = N1223;
  assign { r_n_40__63_, r_n_40__62_, r_n_40__61_, r_n_40__60_, r_n_40__59_, r_n_40__58_, r_n_40__57_, r_n_40__56_, r_n_40__55_, r_n_40__54_, r_n_40__53_, r_n_40__52_, r_n_40__51_, r_n_40__50_, r_n_40__49_, r_n_40__48_, r_n_40__47_, r_n_40__46_, r_n_40__45_, r_n_40__44_, r_n_40__43_, r_n_40__42_, r_n_40__41_, r_n_40__40_, r_n_40__39_, r_n_40__38_, r_n_40__37_, r_n_40__36_, r_n_40__35_, r_n_40__34_, r_n_40__33_, r_n_40__32_, r_n_40__31_, r_n_40__30_, r_n_40__29_, r_n_40__28_, r_n_40__27_, r_n_40__26_, r_n_40__25_, r_n_40__24_, r_n_40__23_, r_n_40__22_, r_n_40__21_, r_n_40__20_, r_n_40__19_, r_n_40__18_, r_n_40__17_, r_n_40__16_, r_n_40__15_, r_n_40__14_, r_n_40__13_, r_n_40__12_, r_n_40__11_, r_n_40__10_, r_n_40__9_, r_n_40__8_, r_n_40__7_, r_n_40__6_, r_n_40__5_, r_n_40__4_, r_n_40__3_, r_n_40__2_, r_n_40__1_, r_n_40__0_ } = (N80)? { r_41__63_, r_41__62_, r_41__61_, r_41__60_, r_41__59_, r_41__58_, r_41__57_, r_41__56_, r_41__55_, r_41__54_, r_41__53_, r_41__52_, r_41__51_, r_41__50_, r_41__49_, r_41__48_, r_41__47_, r_41__46_, r_41__45_, r_41__44_, r_41__43_, r_41__42_, r_41__41_, r_41__40_, r_41__39_, r_41__38_, r_41__37_, r_41__36_, r_41__35_, r_41__34_, r_41__33_, r_41__32_, r_41__31_, r_41__30_, r_41__29_, r_41__28_, r_41__27_, r_41__26_, r_41__25_, r_41__24_, r_41__23_, r_41__22_, r_41__21_, r_41__20_, r_41__19_, r_41__18_, r_41__17_, r_41__16_, r_41__15_, r_41__14_, r_41__13_, r_41__12_, r_41__11_, r_41__10_, r_41__9_, r_41__8_, r_41__7_, r_41__6_, r_41__5_, r_41__4_, r_41__3_, r_41__2_, r_41__1_, r_41__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N81)? data_i : 1'b0;
  assign N80 = sel_i[80];
  assign N81 = N1228;
  assign { r_n_41__63_, r_n_41__62_, r_n_41__61_, r_n_41__60_, r_n_41__59_, r_n_41__58_, r_n_41__57_, r_n_41__56_, r_n_41__55_, r_n_41__54_, r_n_41__53_, r_n_41__52_, r_n_41__51_, r_n_41__50_, r_n_41__49_, r_n_41__48_, r_n_41__47_, r_n_41__46_, r_n_41__45_, r_n_41__44_, r_n_41__43_, r_n_41__42_, r_n_41__41_, r_n_41__40_, r_n_41__39_, r_n_41__38_, r_n_41__37_, r_n_41__36_, r_n_41__35_, r_n_41__34_, r_n_41__33_, r_n_41__32_, r_n_41__31_, r_n_41__30_, r_n_41__29_, r_n_41__28_, r_n_41__27_, r_n_41__26_, r_n_41__25_, r_n_41__24_, r_n_41__23_, r_n_41__22_, r_n_41__21_, r_n_41__20_, r_n_41__19_, r_n_41__18_, r_n_41__17_, r_n_41__16_, r_n_41__15_, r_n_41__14_, r_n_41__13_, r_n_41__12_, r_n_41__11_, r_n_41__10_, r_n_41__9_, r_n_41__8_, r_n_41__7_, r_n_41__6_, r_n_41__5_, r_n_41__4_, r_n_41__3_, r_n_41__2_, r_n_41__1_, r_n_41__0_ } = (N82)? { r_42__63_, r_42__62_, r_42__61_, r_42__60_, r_42__59_, r_42__58_, r_42__57_, r_42__56_, r_42__55_, r_42__54_, r_42__53_, r_42__52_, r_42__51_, r_42__50_, r_42__49_, r_42__48_, r_42__47_, r_42__46_, r_42__45_, r_42__44_, r_42__43_, r_42__42_, r_42__41_, r_42__40_, r_42__39_, r_42__38_, r_42__37_, r_42__36_, r_42__35_, r_42__34_, r_42__33_, r_42__32_, r_42__31_, r_42__30_, r_42__29_, r_42__28_, r_42__27_, r_42__26_, r_42__25_, r_42__24_, r_42__23_, r_42__22_, r_42__21_, r_42__20_, r_42__19_, r_42__18_, r_42__17_, r_42__16_, r_42__15_, r_42__14_, r_42__13_, r_42__12_, r_42__11_, r_42__10_, r_42__9_, r_42__8_, r_42__7_, r_42__6_, r_42__5_, r_42__4_, r_42__3_, r_42__2_, r_42__1_, r_42__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N83)? data_i : 1'b0;
  assign N82 = sel_i[82];
  assign N83 = N1233;
  assign { r_n_42__63_, r_n_42__62_, r_n_42__61_, r_n_42__60_, r_n_42__59_, r_n_42__58_, r_n_42__57_, r_n_42__56_, r_n_42__55_, r_n_42__54_, r_n_42__53_, r_n_42__52_, r_n_42__51_, r_n_42__50_, r_n_42__49_, r_n_42__48_, r_n_42__47_, r_n_42__46_, r_n_42__45_, r_n_42__44_, r_n_42__43_, r_n_42__42_, r_n_42__41_, r_n_42__40_, r_n_42__39_, r_n_42__38_, r_n_42__37_, r_n_42__36_, r_n_42__35_, r_n_42__34_, r_n_42__33_, r_n_42__32_, r_n_42__31_, r_n_42__30_, r_n_42__29_, r_n_42__28_, r_n_42__27_, r_n_42__26_, r_n_42__25_, r_n_42__24_, r_n_42__23_, r_n_42__22_, r_n_42__21_, r_n_42__20_, r_n_42__19_, r_n_42__18_, r_n_42__17_, r_n_42__16_, r_n_42__15_, r_n_42__14_, r_n_42__13_, r_n_42__12_, r_n_42__11_, r_n_42__10_, r_n_42__9_, r_n_42__8_, r_n_42__7_, r_n_42__6_, r_n_42__5_, r_n_42__4_, r_n_42__3_, r_n_42__2_, r_n_42__1_, r_n_42__0_ } = (N84)? { r_43__63_, r_43__62_, r_43__61_, r_43__60_, r_43__59_, r_43__58_, r_43__57_, r_43__56_, r_43__55_, r_43__54_, r_43__53_, r_43__52_, r_43__51_, r_43__50_, r_43__49_, r_43__48_, r_43__47_, r_43__46_, r_43__45_, r_43__44_, r_43__43_, r_43__42_, r_43__41_, r_43__40_, r_43__39_, r_43__38_, r_43__37_, r_43__36_, r_43__35_, r_43__34_, r_43__33_, r_43__32_, r_43__31_, r_43__30_, r_43__29_, r_43__28_, r_43__27_, r_43__26_, r_43__25_, r_43__24_, r_43__23_, r_43__22_, r_43__21_, r_43__20_, r_43__19_, r_43__18_, r_43__17_, r_43__16_, r_43__15_, r_43__14_, r_43__13_, r_43__12_, r_43__11_, r_43__10_, r_43__9_, r_43__8_, r_43__7_, r_43__6_, r_43__5_, r_43__4_, r_43__3_, r_43__2_, r_43__1_, r_43__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N85)? data_i : 1'b0;
  assign N84 = sel_i[84];
  assign N85 = N1238;
  assign { r_n_43__63_, r_n_43__62_, r_n_43__61_, r_n_43__60_, r_n_43__59_, r_n_43__58_, r_n_43__57_, r_n_43__56_, r_n_43__55_, r_n_43__54_, r_n_43__53_, r_n_43__52_, r_n_43__51_, r_n_43__50_, r_n_43__49_, r_n_43__48_, r_n_43__47_, r_n_43__46_, r_n_43__45_, r_n_43__44_, r_n_43__43_, r_n_43__42_, r_n_43__41_, r_n_43__40_, r_n_43__39_, r_n_43__38_, r_n_43__37_, r_n_43__36_, r_n_43__35_, r_n_43__34_, r_n_43__33_, r_n_43__32_, r_n_43__31_, r_n_43__30_, r_n_43__29_, r_n_43__28_, r_n_43__27_, r_n_43__26_, r_n_43__25_, r_n_43__24_, r_n_43__23_, r_n_43__22_, r_n_43__21_, r_n_43__20_, r_n_43__19_, r_n_43__18_, r_n_43__17_, r_n_43__16_, r_n_43__15_, r_n_43__14_, r_n_43__13_, r_n_43__12_, r_n_43__11_, r_n_43__10_, r_n_43__9_, r_n_43__8_, r_n_43__7_, r_n_43__6_, r_n_43__5_, r_n_43__4_, r_n_43__3_, r_n_43__2_, r_n_43__1_, r_n_43__0_ } = (N86)? { r_44__63_, r_44__62_, r_44__61_, r_44__60_, r_44__59_, r_44__58_, r_44__57_, r_44__56_, r_44__55_, r_44__54_, r_44__53_, r_44__52_, r_44__51_, r_44__50_, r_44__49_, r_44__48_, r_44__47_, r_44__46_, r_44__45_, r_44__44_, r_44__43_, r_44__42_, r_44__41_, r_44__40_, r_44__39_, r_44__38_, r_44__37_, r_44__36_, r_44__35_, r_44__34_, r_44__33_, r_44__32_, r_44__31_, r_44__30_, r_44__29_, r_44__28_, r_44__27_, r_44__26_, r_44__25_, r_44__24_, r_44__23_, r_44__22_, r_44__21_, r_44__20_, r_44__19_, r_44__18_, r_44__17_, r_44__16_, r_44__15_, r_44__14_, r_44__13_, r_44__12_, r_44__11_, r_44__10_, r_44__9_, r_44__8_, r_44__7_, r_44__6_, r_44__5_, r_44__4_, r_44__3_, r_44__2_, r_44__1_, r_44__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N87)? data_i : 1'b0;
  assign N86 = sel_i[86];
  assign N87 = N1243;
  assign { r_n_44__63_, r_n_44__62_, r_n_44__61_, r_n_44__60_, r_n_44__59_, r_n_44__58_, r_n_44__57_, r_n_44__56_, r_n_44__55_, r_n_44__54_, r_n_44__53_, r_n_44__52_, r_n_44__51_, r_n_44__50_, r_n_44__49_, r_n_44__48_, r_n_44__47_, r_n_44__46_, r_n_44__45_, r_n_44__44_, r_n_44__43_, r_n_44__42_, r_n_44__41_, r_n_44__40_, r_n_44__39_, r_n_44__38_, r_n_44__37_, r_n_44__36_, r_n_44__35_, r_n_44__34_, r_n_44__33_, r_n_44__32_, r_n_44__31_, r_n_44__30_, r_n_44__29_, r_n_44__28_, r_n_44__27_, r_n_44__26_, r_n_44__25_, r_n_44__24_, r_n_44__23_, r_n_44__22_, r_n_44__21_, r_n_44__20_, r_n_44__19_, r_n_44__18_, r_n_44__17_, r_n_44__16_, r_n_44__15_, r_n_44__14_, r_n_44__13_, r_n_44__12_, r_n_44__11_, r_n_44__10_, r_n_44__9_, r_n_44__8_, r_n_44__7_, r_n_44__6_, r_n_44__5_, r_n_44__4_, r_n_44__3_, r_n_44__2_, r_n_44__1_, r_n_44__0_ } = (N88)? { r_45__63_, r_45__62_, r_45__61_, r_45__60_, r_45__59_, r_45__58_, r_45__57_, r_45__56_, r_45__55_, r_45__54_, r_45__53_, r_45__52_, r_45__51_, r_45__50_, r_45__49_, r_45__48_, r_45__47_, r_45__46_, r_45__45_, r_45__44_, r_45__43_, r_45__42_, r_45__41_, r_45__40_, r_45__39_, r_45__38_, r_45__37_, r_45__36_, r_45__35_, r_45__34_, r_45__33_, r_45__32_, r_45__31_, r_45__30_, r_45__29_, r_45__28_, r_45__27_, r_45__26_, r_45__25_, r_45__24_, r_45__23_, r_45__22_, r_45__21_, r_45__20_, r_45__19_, r_45__18_, r_45__17_, r_45__16_, r_45__15_, r_45__14_, r_45__13_, r_45__12_, r_45__11_, r_45__10_, r_45__9_, r_45__8_, r_45__7_, r_45__6_, r_45__5_, r_45__4_, r_45__3_, r_45__2_, r_45__1_, r_45__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N89)? data_i : 1'b0;
  assign N88 = sel_i[88];
  assign N89 = N1248;
  assign { r_n_45__63_, r_n_45__62_, r_n_45__61_, r_n_45__60_, r_n_45__59_, r_n_45__58_, r_n_45__57_, r_n_45__56_, r_n_45__55_, r_n_45__54_, r_n_45__53_, r_n_45__52_, r_n_45__51_, r_n_45__50_, r_n_45__49_, r_n_45__48_, r_n_45__47_, r_n_45__46_, r_n_45__45_, r_n_45__44_, r_n_45__43_, r_n_45__42_, r_n_45__41_, r_n_45__40_, r_n_45__39_, r_n_45__38_, r_n_45__37_, r_n_45__36_, r_n_45__35_, r_n_45__34_, r_n_45__33_, r_n_45__32_, r_n_45__31_, r_n_45__30_, r_n_45__29_, r_n_45__28_, r_n_45__27_, r_n_45__26_, r_n_45__25_, r_n_45__24_, r_n_45__23_, r_n_45__22_, r_n_45__21_, r_n_45__20_, r_n_45__19_, r_n_45__18_, r_n_45__17_, r_n_45__16_, r_n_45__15_, r_n_45__14_, r_n_45__13_, r_n_45__12_, r_n_45__11_, r_n_45__10_, r_n_45__9_, r_n_45__8_, r_n_45__7_, r_n_45__6_, r_n_45__5_, r_n_45__4_, r_n_45__3_, r_n_45__2_, r_n_45__1_, r_n_45__0_ } = (N90)? { r_46__63_, r_46__62_, r_46__61_, r_46__60_, r_46__59_, r_46__58_, r_46__57_, r_46__56_, r_46__55_, r_46__54_, r_46__53_, r_46__52_, r_46__51_, r_46__50_, r_46__49_, r_46__48_, r_46__47_, r_46__46_, r_46__45_, r_46__44_, r_46__43_, r_46__42_, r_46__41_, r_46__40_, r_46__39_, r_46__38_, r_46__37_, r_46__36_, r_46__35_, r_46__34_, r_46__33_, r_46__32_, r_46__31_, r_46__30_, r_46__29_, r_46__28_, r_46__27_, r_46__26_, r_46__25_, r_46__24_, r_46__23_, r_46__22_, r_46__21_, r_46__20_, r_46__19_, r_46__18_, r_46__17_, r_46__16_, r_46__15_, r_46__14_, r_46__13_, r_46__12_, r_46__11_, r_46__10_, r_46__9_, r_46__8_, r_46__7_, r_46__6_, r_46__5_, r_46__4_, r_46__3_, r_46__2_, r_46__1_, r_46__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N91)? data_i : 1'b0;
  assign N90 = sel_i[90];
  assign N91 = N1253;
  assign { r_n_46__63_, r_n_46__62_, r_n_46__61_, r_n_46__60_, r_n_46__59_, r_n_46__58_, r_n_46__57_, r_n_46__56_, r_n_46__55_, r_n_46__54_, r_n_46__53_, r_n_46__52_, r_n_46__51_, r_n_46__50_, r_n_46__49_, r_n_46__48_, r_n_46__47_, r_n_46__46_, r_n_46__45_, r_n_46__44_, r_n_46__43_, r_n_46__42_, r_n_46__41_, r_n_46__40_, r_n_46__39_, r_n_46__38_, r_n_46__37_, r_n_46__36_, r_n_46__35_, r_n_46__34_, r_n_46__33_, r_n_46__32_, r_n_46__31_, r_n_46__30_, r_n_46__29_, r_n_46__28_, r_n_46__27_, r_n_46__26_, r_n_46__25_, r_n_46__24_, r_n_46__23_, r_n_46__22_, r_n_46__21_, r_n_46__20_, r_n_46__19_, r_n_46__18_, r_n_46__17_, r_n_46__16_, r_n_46__15_, r_n_46__14_, r_n_46__13_, r_n_46__12_, r_n_46__11_, r_n_46__10_, r_n_46__9_, r_n_46__8_, r_n_46__7_, r_n_46__6_, r_n_46__5_, r_n_46__4_, r_n_46__3_, r_n_46__2_, r_n_46__1_, r_n_46__0_ } = (N92)? { r_47__63_, r_47__62_, r_47__61_, r_47__60_, r_47__59_, r_47__58_, r_47__57_, r_47__56_, r_47__55_, r_47__54_, r_47__53_, r_47__52_, r_47__51_, r_47__50_, r_47__49_, r_47__48_, r_47__47_, r_47__46_, r_47__45_, r_47__44_, r_47__43_, r_47__42_, r_47__41_, r_47__40_, r_47__39_, r_47__38_, r_47__37_, r_47__36_, r_47__35_, r_47__34_, r_47__33_, r_47__32_, r_47__31_, r_47__30_, r_47__29_, r_47__28_, r_47__27_, r_47__26_, r_47__25_, r_47__24_, r_47__23_, r_47__22_, r_47__21_, r_47__20_, r_47__19_, r_47__18_, r_47__17_, r_47__16_, r_47__15_, r_47__14_, r_47__13_, r_47__12_, r_47__11_, r_47__10_, r_47__9_, r_47__8_, r_47__7_, r_47__6_, r_47__5_, r_47__4_, r_47__3_, r_47__2_, r_47__1_, r_47__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N93)? data_i : 1'b0;
  assign N92 = sel_i[92];
  assign N93 = N1258;
  assign { r_n_47__63_, r_n_47__62_, r_n_47__61_, r_n_47__60_, r_n_47__59_, r_n_47__58_, r_n_47__57_, r_n_47__56_, r_n_47__55_, r_n_47__54_, r_n_47__53_, r_n_47__52_, r_n_47__51_, r_n_47__50_, r_n_47__49_, r_n_47__48_, r_n_47__47_, r_n_47__46_, r_n_47__45_, r_n_47__44_, r_n_47__43_, r_n_47__42_, r_n_47__41_, r_n_47__40_, r_n_47__39_, r_n_47__38_, r_n_47__37_, r_n_47__36_, r_n_47__35_, r_n_47__34_, r_n_47__33_, r_n_47__32_, r_n_47__31_, r_n_47__30_, r_n_47__29_, r_n_47__28_, r_n_47__27_, r_n_47__26_, r_n_47__25_, r_n_47__24_, r_n_47__23_, r_n_47__22_, r_n_47__21_, r_n_47__20_, r_n_47__19_, r_n_47__18_, r_n_47__17_, r_n_47__16_, r_n_47__15_, r_n_47__14_, r_n_47__13_, r_n_47__12_, r_n_47__11_, r_n_47__10_, r_n_47__9_, r_n_47__8_, r_n_47__7_, r_n_47__6_, r_n_47__5_, r_n_47__4_, r_n_47__3_, r_n_47__2_, r_n_47__1_, r_n_47__0_ } = (N94)? { r_48__63_, r_48__62_, r_48__61_, r_48__60_, r_48__59_, r_48__58_, r_48__57_, r_48__56_, r_48__55_, r_48__54_, r_48__53_, r_48__52_, r_48__51_, r_48__50_, r_48__49_, r_48__48_, r_48__47_, r_48__46_, r_48__45_, r_48__44_, r_48__43_, r_48__42_, r_48__41_, r_48__40_, r_48__39_, r_48__38_, r_48__37_, r_48__36_, r_48__35_, r_48__34_, r_48__33_, r_48__32_, r_48__31_, r_48__30_, r_48__29_, r_48__28_, r_48__27_, r_48__26_, r_48__25_, r_48__24_, r_48__23_, r_48__22_, r_48__21_, r_48__20_, r_48__19_, r_48__18_, r_48__17_, r_48__16_, r_48__15_, r_48__14_, r_48__13_, r_48__12_, r_48__11_, r_48__10_, r_48__9_, r_48__8_, r_48__7_, r_48__6_, r_48__5_, r_48__4_, r_48__3_, r_48__2_, r_48__1_, r_48__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N95)? data_i : 1'b0;
  assign N94 = sel_i[94];
  assign N95 = N1263;
  assign { r_n_48__63_, r_n_48__62_, r_n_48__61_, r_n_48__60_, r_n_48__59_, r_n_48__58_, r_n_48__57_, r_n_48__56_, r_n_48__55_, r_n_48__54_, r_n_48__53_, r_n_48__52_, r_n_48__51_, r_n_48__50_, r_n_48__49_, r_n_48__48_, r_n_48__47_, r_n_48__46_, r_n_48__45_, r_n_48__44_, r_n_48__43_, r_n_48__42_, r_n_48__41_, r_n_48__40_, r_n_48__39_, r_n_48__38_, r_n_48__37_, r_n_48__36_, r_n_48__35_, r_n_48__34_, r_n_48__33_, r_n_48__32_, r_n_48__31_, r_n_48__30_, r_n_48__29_, r_n_48__28_, r_n_48__27_, r_n_48__26_, r_n_48__25_, r_n_48__24_, r_n_48__23_, r_n_48__22_, r_n_48__21_, r_n_48__20_, r_n_48__19_, r_n_48__18_, r_n_48__17_, r_n_48__16_, r_n_48__15_, r_n_48__14_, r_n_48__13_, r_n_48__12_, r_n_48__11_, r_n_48__10_, r_n_48__9_, r_n_48__8_, r_n_48__7_, r_n_48__6_, r_n_48__5_, r_n_48__4_, r_n_48__3_, r_n_48__2_, r_n_48__1_, r_n_48__0_ } = (N96)? { r_49__63_, r_49__62_, r_49__61_, r_49__60_, r_49__59_, r_49__58_, r_49__57_, r_49__56_, r_49__55_, r_49__54_, r_49__53_, r_49__52_, r_49__51_, r_49__50_, r_49__49_, r_49__48_, r_49__47_, r_49__46_, r_49__45_, r_49__44_, r_49__43_, r_49__42_, r_49__41_, r_49__40_, r_49__39_, r_49__38_, r_49__37_, r_49__36_, r_49__35_, r_49__34_, r_49__33_, r_49__32_, r_49__31_, r_49__30_, r_49__29_, r_49__28_, r_49__27_, r_49__26_, r_49__25_, r_49__24_, r_49__23_, r_49__22_, r_49__21_, r_49__20_, r_49__19_, r_49__18_, r_49__17_, r_49__16_, r_49__15_, r_49__14_, r_49__13_, r_49__12_, r_49__11_, r_49__10_, r_49__9_, r_49__8_, r_49__7_, r_49__6_, r_49__5_, r_49__4_, r_49__3_, r_49__2_, r_49__1_, r_49__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N97)? data_i : 1'b0;
  assign N96 = sel_i[96];
  assign N97 = N1268;
  assign { r_n_49__63_, r_n_49__62_, r_n_49__61_, r_n_49__60_, r_n_49__59_, r_n_49__58_, r_n_49__57_, r_n_49__56_, r_n_49__55_, r_n_49__54_, r_n_49__53_, r_n_49__52_, r_n_49__51_, r_n_49__50_, r_n_49__49_, r_n_49__48_, r_n_49__47_, r_n_49__46_, r_n_49__45_, r_n_49__44_, r_n_49__43_, r_n_49__42_, r_n_49__41_, r_n_49__40_, r_n_49__39_, r_n_49__38_, r_n_49__37_, r_n_49__36_, r_n_49__35_, r_n_49__34_, r_n_49__33_, r_n_49__32_, r_n_49__31_, r_n_49__30_, r_n_49__29_, r_n_49__28_, r_n_49__27_, r_n_49__26_, r_n_49__25_, r_n_49__24_, r_n_49__23_, r_n_49__22_, r_n_49__21_, r_n_49__20_, r_n_49__19_, r_n_49__18_, r_n_49__17_, r_n_49__16_, r_n_49__15_, r_n_49__14_, r_n_49__13_, r_n_49__12_, r_n_49__11_, r_n_49__10_, r_n_49__9_, r_n_49__8_, r_n_49__7_, r_n_49__6_, r_n_49__5_, r_n_49__4_, r_n_49__3_, r_n_49__2_, r_n_49__1_, r_n_49__0_ } = (N98)? { r_50__63_, r_50__62_, r_50__61_, r_50__60_, r_50__59_, r_50__58_, r_50__57_, r_50__56_, r_50__55_, r_50__54_, r_50__53_, r_50__52_, r_50__51_, r_50__50_, r_50__49_, r_50__48_, r_50__47_, r_50__46_, r_50__45_, r_50__44_, r_50__43_, r_50__42_, r_50__41_, r_50__40_, r_50__39_, r_50__38_, r_50__37_, r_50__36_, r_50__35_, r_50__34_, r_50__33_, r_50__32_, r_50__31_, r_50__30_, r_50__29_, r_50__28_, r_50__27_, r_50__26_, r_50__25_, r_50__24_, r_50__23_, r_50__22_, r_50__21_, r_50__20_, r_50__19_, r_50__18_, r_50__17_, r_50__16_, r_50__15_, r_50__14_, r_50__13_, r_50__12_, r_50__11_, r_50__10_, r_50__9_, r_50__8_, r_50__7_, r_50__6_, r_50__5_, r_50__4_, r_50__3_, r_50__2_, r_50__1_, r_50__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N99)? data_i : 1'b0;
  assign N98 = sel_i[98];
  assign N99 = N1273;
  assign { r_n_50__63_, r_n_50__62_, r_n_50__61_, r_n_50__60_, r_n_50__59_, r_n_50__58_, r_n_50__57_, r_n_50__56_, r_n_50__55_, r_n_50__54_, r_n_50__53_, r_n_50__52_, r_n_50__51_, r_n_50__50_, r_n_50__49_, r_n_50__48_, r_n_50__47_, r_n_50__46_, r_n_50__45_, r_n_50__44_, r_n_50__43_, r_n_50__42_, r_n_50__41_, r_n_50__40_, r_n_50__39_, r_n_50__38_, r_n_50__37_, r_n_50__36_, r_n_50__35_, r_n_50__34_, r_n_50__33_, r_n_50__32_, r_n_50__31_, r_n_50__30_, r_n_50__29_, r_n_50__28_, r_n_50__27_, r_n_50__26_, r_n_50__25_, r_n_50__24_, r_n_50__23_, r_n_50__22_, r_n_50__21_, r_n_50__20_, r_n_50__19_, r_n_50__18_, r_n_50__17_, r_n_50__16_, r_n_50__15_, r_n_50__14_, r_n_50__13_, r_n_50__12_, r_n_50__11_, r_n_50__10_, r_n_50__9_, r_n_50__8_, r_n_50__7_, r_n_50__6_, r_n_50__5_, r_n_50__4_, r_n_50__3_, r_n_50__2_, r_n_50__1_, r_n_50__0_ } = (N100)? { r_51__63_, r_51__62_, r_51__61_, r_51__60_, r_51__59_, r_51__58_, r_51__57_, r_51__56_, r_51__55_, r_51__54_, r_51__53_, r_51__52_, r_51__51_, r_51__50_, r_51__49_, r_51__48_, r_51__47_, r_51__46_, r_51__45_, r_51__44_, r_51__43_, r_51__42_, r_51__41_, r_51__40_, r_51__39_, r_51__38_, r_51__37_, r_51__36_, r_51__35_, r_51__34_, r_51__33_, r_51__32_, r_51__31_, r_51__30_, r_51__29_, r_51__28_, r_51__27_, r_51__26_, r_51__25_, r_51__24_, r_51__23_, r_51__22_, r_51__21_, r_51__20_, r_51__19_, r_51__18_, r_51__17_, r_51__16_, r_51__15_, r_51__14_, r_51__13_, r_51__12_, r_51__11_, r_51__10_, r_51__9_, r_51__8_, r_51__7_, r_51__6_, r_51__5_, r_51__4_, r_51__3_, r_51__2_, r_51__1_, r_51__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N101)? data_i : 1'b0;
  assign N100 = sel_i[100];
  assign N101 = N1278;
  assign { r_n_51__63_, r_n_51__62_, r_n_51__61_, r_n_51__60_, r_n_51__59_, r_n_51__58_, r_n_51__57_, r_n_51__56_, r_n_51__55_, r_n_51__54_, r_n_51__53_, r_n_51__52_, r_n_51__51_, r_n_51__50_, r_n_51__49_, r_n_51__48_, r_n_51__47_, r_n_51__46_, r_n_51__45_, r_n_51__44_, r_n_51__43_, r_n_51__42_, r_n_51__41_, r_n_51__40_, r_n_51__39_, r_n_51__38_, r_n_51__37_, r_n_51__36_, r_n_51__35_, r_n_51__34_, r_n_51__33_, r_n_51__32_, r_n_51__31_, r_n_51__30_, r_n_51__29_, r_n_51__28_, r_n_51__27_, r_n_51__26_, r_n_51__25_, r_n_51__24_, r_n_51__23_, r_n_51__22_, r_n_51__21_, r_n_51__20_, r_n_51__19_, r_n_51__18_, r_n_51__17_, r_n_51__16_, r_n_51__15_, r_n_51__14_, r_n_51__13_, r_n_51__12_, r_n_51__11_, r_n_51__10_, r_n_51__9_, r_n_51__8_, r_n_51__7_, r_n_51__6_, r_n_51__5_, r_n_51__4_, r_n_51__3_, r_n_51__2_, r_n_51__1_, r_n_51__0_ } = (N102)? { r_52__63_, r_52__62_, r_52__61_, r_52__60_, r_52__59_, r_52__58_, r_52__57_, r_52__56_, r_52__55_, r_52__54_, r_52__53_, r_52__52_, r_52__51_, r_52__50_, r_52__49_, r_52__48_, r_52__47_, r_52__46_, r_52__45_, r_52__44_, r_52__43_, r_52__42_, r_52__41_, r_52__40_, r_52__39_, r_52__38_, r_52__37_, r_52__36_, r_52__35_, r_52__34_, r_52__33_, r_52__32_, r_52__31_, r_52__30_, r_52__29_, r_52__28_, r_52__27_, r_52__26_, r_52__25_, r_52__24_, r_52__23_, r_52__22_, r_52__21_, r_52__20_, r_52__19_, r_52__18_, r_52__17_, r_52__16_, r_52__15_, r_52__14_, r_52__13_, r_52__12_, r_52__11_, r_52__10_, r_52__9_, r_52__8_, r_52__7_, r_52__6_, r_52__5_, r_52__4_, r_52__3_, r_52__2_, r_52__1_, r_52__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N103)? data_i : 1'b0;
  assign N102 = sel_i[102];
  assign N103 = N1283;
  assign { r_n_52__63_, r_n_52__62_, r_n_52__61_, r_n_52__60_, r_n_52__59_, r_n_52__58_, r_n_52__57_, r_n_52__56_, r_n_52__55_, r_n_52__54_, r_n_52__53_, r_n_52__52_, r_n_52__51_, r_n_52__50_, r_n_52__49_, r_n_52__48_, r_n_52__47_, r_n_52__46_, r_n_52__45_, r_n_52__44_, r_n_52__43_, r_n_52__42_, r_n_52__41_, r_n_52__40_, r_n_52__39_, r_n_52__38_, r_n_52__37_, r_n_52__36_, r_n_52__35_, r_n_52__34_, r_n_52__33_, r_n_52__32_, r_n_52__31_, r_n_52__30_, r_n_52__29_, r_n_52__28_, r_n_52__27_, r_n_52__26_, r_n_52__25_, r_n_52__24_, r_n_52__23_, r_n_52__22_, r_n_52__21_, r_n_52__20_, r_n_52__19_, r_n_52__18_, r_n_52__17_, r_n_52__16_, r_n_52__15_, r_n_52__14_, r_n_52__13_, r_n_52__12_, r_n_52__11_, r_n_52__10_, r_n_52__9_, r_n_52__8_, r_n_52__7_, r_n_52__6_, r_n_52__5_, r_n_52__4_, r_n_52__3_, r_n_52__2_, r_n_52__1_, r_n_52__0_ } = (N104)? { r_53__63_, r_53__62_, r_53__61_, r_53__60_, r_53__59_, r_53__58_, r_53__57_, r_53__56_, r_53__55_, r_53__54_, r_53__53_, r_53__52_, r_53__51_, r_53__50_, r_53__49_, r_53__48_, r_53__47_, r_53__46_, r_53__45_, r_53__44_, r_53__43_, r_53__42_, r_53__41_, r_53__40_, r_53__39_, r_53__38_, r_53__37_, r_53__36_, r_53__35_, r_53__34_, r_53__33_, r_53__32_, r_53__31_, r_53__30_, r_53__29_, r_53__28_, r_53__27_, r_53__26_, r_53__25_, r_53__24_, r_53__23_, r_53__22_, r_53__21_, r_53__20_, r_53__19_, r_53__18_, r_53__17_, r_53__16_, r_53__15_, r_53__14_, r_53__13_, r_53__12_, r_53__11_, r_53__10_, r_53__9_, r_53__8_, r_53__7_, r_53__6_, r_53__5_, r_53__4_, r_53__3_, r_53__2_, r_53__1_, r_53__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N105)? data_i : 1'b0;
  assign N104 = sel_i[104];
  assign N105 = N1288;
  assign { r_n_53__63_, r_n_53__62_, r_n_53__61_, r_n_53__60_, r_n_53__59_, r_n_53__58_, r_n_53__57_, r_n_53__56_, r_n_53__55_, r_n_53__54_, r_n_53__53_, r_n_53__52_, r_n_53__51_, r_n_53__50_, r_n_53__49_, r_n_53__48_, r_n_53__47_, r_n_53__46_, r_n_53__45_, r_n_53__44_, r_n_53__43_, r_n_53__42_, r_n_53__41_, r_n_53__40_, r_n_53__39_, r_n_53__38_, r_n_53__37_, r_n_53__36_, r_n_53__35_, r_n_53__34_, r_n_53__33_, r_n_53__32_, r_n_53__31_, r_n_53__30_, r_n_53__29_, r_n_53__28_, r_n_53__27_, r_n_53__26_, r_n_53__25_, r_n_53__24_, r_n_53__23_, r_n_53__22_, r_n_53__21_, r_n_53__20_, r_n_53__19_, r_n_53__18_, r_n_53__17_, r_n_53__16_, r_n_53__15_, r_n_53__14_, r_n_53__13_, r_n_53__12_, r_n_53__11_, r_n_53__10_, r_n_53__9_, r_n_53__8_, r_n_53__7_, r_n_53__6_, r_n_53__5_, r_n_53__4_, r_n_53__3_, r_n_53__2_, r_n_53__1_, r_n_53__0_ } = (N106)? { r_54__63_, r_54__62_, r_54__61_, r_54__60_, r_54__59_, r_54__58_, r_54__57_, r_54__56_, r_54__55_, r_54__54_, r_54__53_, r_54__52_, r_54__51_, r_54__50_, r_54__49_, r_54__48_, r_54__47_, r_54__46_, r_54__45_, r_54__44_, r_54__43_, r_54__42_, r_54__41_, r_54__40_, r_54__39_, r_54__38_, r_54__37_, r_54__36_, r_54__35_, r_54__34_, r_54__33_, r_54__32_, r_54__31_, r_54__30_, r_54__29_, r_54__28_, r_54__27_, r_54__26_, r_54__25_, r_54__24_, r_54__23_, r_54__22_, r_54__21_, r_54__20_, r_54__19_, r_54__18_, r_54__17_, r_54__16_, r_54__15_, r_54__14_, r_54__13_, r_54__12_, r_54__11_, r_54__10_, r_54__9_, r_54__8_, r_54__7_, r_54__6_, r_54__5_, r_54__4_, r_54__3_, r_54__2_, r_54__1_, r_54__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N107)? data_i : 1'b0;
  assign N106 = sel_i[106];
  assign N107 = N1293;
  assign { r_n_54__63_, r_n_54__62_, r_n_54__61_, r_n_54__60_, r_n_54__59_, r_n_54__58_, r_n_54__57_, r_n_54__56_, r_n_54__55_, r_n_54__54_, r_n_54__53_, r_n_54__52_, r_n_54__51_, r_n_54__50_, r_n_54__49_, r_n_54__48_, r_n_54__47_, r_n_54__46_, r_n_54__45_, r_n_54__44_, r_n_54__43_, r_n_54__42_, r_n_54__41_, r_n_54__40_, r_n_54__39_, r_n_54__38_, r_n_54__37_, r_n_54__36_, r_n_54__35_, r_n_54__34_, r_n_54__33_, r_n_54__32_, r_n_54__31_, r_n_54__30_, r_n_54__29_, r_n_54__28_, r_n_54__27_, r_n_54__26_, r_n_54__25_, r_n_54__24_, r_n_54__23_, r_n_54__22_, r_n_54__21_, r_n_54__20_, r_n_54__19_, r_n_54__18_, r_n_54__17_, r_n_54__16_, r_n_54__15_, r_n_54__14_, r_n_54__13_, r_n_54__12_, r_n_54__11_, r_n_54__10_, r_n_54__9_, r_n_54__8_, r_n_54__7_, r_n_54__6_, r_n_54__5_, r_n_54__4_, r_n_54__3_, r_n_54__2_, r_n_54__1_, r_n_54__0_ } = (N108)? { r_55__63_, r_55__62_, r_55__61_, r_55__60_, r_55__59_, r_55__58_, r_55__57_, r_55__56_, r_55__55_, r_55__54_, r_55__53_, r_55__52_, r_55__51_, r_55__50_, r_55__49_, r_55__48_, r_55__47_, r_55__46_, r_55__45_, r_55__44_, r_55__43_, r_55__42_, r_55__41_, r_55__40_, r_55__39_, r_55__38_, r_55__37_, r_55__36_, r_55__35_, r_55__34_, r_55__33_, r_55__32_, r_55__31_, r_55__30_, r_55__29_, r_55__28_, r_55__27_, r_55__26_, r_55__25_, r_55__24_, r_55__23_, r_55__22_, r_55__21_, r_55__20_, r_55__19_, r_55__18_, r_55__17_, r_55__16_, r_55__15_, r_55__14_, r_55__13_, r_55__12_, r_55__11_, r_55__10_, r_55__9_, r_55__8_, r_55__7_, r_55__6_, r_55__5_, r_55__4_, r_55__3_, r_55__2_, r_55__1_, r_55__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N109)? data_i : 1'b0;
  assign N108 = sel_i[108];
  assign N109 = N1298;
  assign { r_n_55__63_, r_n_55__62_, r_n_55__61_, r_n_55__60_, r_n_55__59_, r_n_55__58_, r_n_55__57_, r_n_55__56_, r_n_55__55_, r_n_55__54_, r_n_55__53_, r_n_55__52_, r_n_55__51_, r_n_55__50_, r_n_55__49_, r_n_55__48_, r_n_55__47_, r_n_55__46_, r_n_55__45_, r_n_55__44_, r_n_55__43_, r_n_55__42_, r_n_55__41_, r_n_55__40_, r_n_55__39_, r_n_55__38_, r_n_55__37_, r_n_55__36_, r_n_55__35_, r_n_55__34_, r_n_55__33_, r_n_55__32_, r_n_55__31_, r_n_55__30_, r_n_55__29_, r_n_55__28_, r_n_55__27_, r_n_55__26_, r_n_55__25_, r_n_55__24_, r_n_55__23_, r_n_55__22_, r_n_55__21_, r_n_55__20_, r_n_55__19_, r_n_55__18_, r_n_55__17_, r_n_55__16_, r_n_55__15_, r_n_55__14_, r_n_55__13_, r_n_55__12_, r_n_55__11_, r_n_55__10_, r_n_55__9_, r_n_55__8_, r_n_55__7_, r_n_55__6_, r_n_55__5_, r_n_55__4_, r_n_55__3_, r_n_55__2_, r_n_55__1_, r_n_55__0_ } = (N110)? { r_56__63_, r_56__62_, r_56__61_, r_56__60_, r_56__59_, r_56__58_, r_56__57_, r_56__56_, r_56__55_, r_56__54_, r_56__53_, r_56__52_, r_56__51_, r_56__50_, r_56__49_, r_56__48_, r_56__47_, r_56__46_, r_56__45_, r_56__44_, r_56__43_, r_56__42_, r_56__41_, r_56__40_, r_56__39_, r_56__38_, r_56__37_, r_56__36_, r_56__35_, r_56__34_, r_56__33_, r_56__32_, r_56__31_, r_56__30_, r_56__29_, r_56__28_, r_56__27_, r_56__26_, r_56__25_, r_56__24_, r_56__23_, r_56__22_, r_56__21_, r_56__20_, r_56__19_, r_56__18_, r_56__17_, r_56__16_, r_56__15_, r_56__14_, r_56__13_, r_56__12_, r_56__11_, r_56__10_, r_56__9_, r_56__8_, r_56__7_, r_56__6_, r_56__5_, r_56__4_, r_56__3_, r_56__2_, r_56__1_, r_56__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N111)? data_i : 1'b0;
  assign N110 = sel_i[110];
  assign N111 = N1303;
  assign { r_n_56__63_, r_n_56__62_, r_n_56__61_, r_n_56__60_, r_n_56__59_, r_n_56__58_, r_n_56__57_, r_n_56__56_, r_n_56__55_, r_n_56__54_, r_n_56__53_, r_n_56__52_, r_n_56__51_, r_n_56__50_, r_n_56__49_, r_n_56__48_, r_n_56__47_, r_n_56__46_, r_n_56__45_, r_n_56__44_, r_n_56__43_, r_n_56__42_, r_n_56__41_, r_n_56__40_, r_n_56__39_, r_n_56__38_, r_n_56__37_, r_n_56__36_, r_n_56__35_, r_n_56__34_, r_n_56__33_, r_n_56__32_, r_n_56__31_, r_n_56__30_, r_n_56__29_, r_n_56__28_, r_n_56__27_, r_n_56__26_, r_n_56__25_, r_n_56__24_, r_n_56__23_, r_n_56__22_, r_n_56__21_, r_n_56__20_, r_n_56__19_, r_n_56__18_, r_n_56__17_, r_n_56__16_, r_n_56__15_, r_n_56__14_, r_n_56__13_, r_n_56__12_, r_n_56__11_, r_n_56__10_, r_n_56__9_, r_n_56__8_, r_n_56__7_, r_n_56__6_, r_n_56__5_, r_n_56__4_, r_n_56__3_, r_n_56__2_, r_n_56__1_, r_n_56__0_ } = (N112)? { r_57__63_, r_57__62_, r_57__61_, r_57__60_, r_57__59_, r_57__58_, r_57__57_, r_57__56_, r_57__55_, r_57__54_, r_57__53_, r_57__52_, r_57__51_, r_57__50_, r_57__49_, r_57__48_, r_57__47_, r_57__46_, r_57__45_, r_57__44_, r_57__43_, r_57__42_, r_57__41_, r_57__40_, r_57__39_, r_57__38_, r_57__37_, r_57__36_, r_57__35_, r_57__34_, r_57__33_, r_57__32_, r_57__31_, r_57__30_, r_57__29_, r_57__28_, r_57__27_, r_57__26_, r_57__25_, r_57__24_, r_57__23_, r_57__22_, r_57__21_, r_57__20_, r_57__19_, r_57__18_, r_57__17_, r_57__16_, r_57__15_, r_57__14_, r_57__13_, r_57__12_, r_57__11_, r_57__10_, r_57__9_, r_57__8_, r_57__7_, r_57__6_, r_57__5_, r_57__4_, r_57__3_, r_57__2_, r_57__1_, r_57__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N113)? data_i : 1'b0;
  assign N112 = sel_i[112];
  assign N113 = N1308;
  assign { r_n_57__63_, r_n_57__62_, r_n_57__61_, r_n_57__60_, r_n_57__59_, r_n_57__58_, r_n_57__57_, r_n_57__56_, r_n_57__55_, r_n_57__54_, r_n_57__53_, r_n_57__52_, r_n_57__51_, r_n_57__50_, r_n_57__49_, r_n_57__48_, r_n_57__47_, r_n_57__46_, r_n_57__45_, r_n_57__44_, r_n_57__43_, r_n_57__42_, r_n_57__41_, r_n_57__40_, r_n_57__39_, r_n_57__38_, r_n_57__37_, r_n_57__36_, r_n_57__35_, r_n_57__34_, r_n_57__33_, r_n_57__32_, r_n_57__31_, r_n_57__30_, r_n_57__29_, r_n_57__28_, r_n_57__27_, r_n_57__26_, r_n_57__25_, r_n_57__24_, r_n_57__23_, r_n_57__22_, r_n_57__21_, r_n_57__20_, r_n_57__19_, r_n_57__18_, r_n_57__17_, r_n_57__16_, r_n_57__15_, r_n_57__14_, r_n_57__13_, r_n_57__12_, r_n_57__11_, r_n_57__10_, r_n_57__9_, r_n_57__8_, r_n_57__7_, r_n_57__6_, r_n_57__5_, r_n_57__4_, r_n_57__3_, r_n_57__2_, r_n_57__1_, r_n_57__0_ } = (N114)? { r_58__63_, r_58__62_, r_58__61_, r_58__60_, r_58__59_, r_58__58_, r_58__57_, r_58__56_, r_58__55_, r_58__54_, r_58__53_, r_58__52_, r_58__51_, r_58__50_, r_58__49_, r_58__48_, r_58__47_, r_58__46_, r_58__45_, r_58__44_, r_58__43_, r_58__42_, r_58__41_, r_58__40_, r_58__39_, r_58__38_, r_58__37_, r_58__36_, r_58__35_, r_58__34_, r_58__33_, r_58__32_, r_58__31_, r_58__30_, r_58__29_, r_58__28_, r_58__27_, r_58__26_, r_58__25_, r_58__24_, r_58__23_, r_58__22_, r_58__21_, r_58__20_, r_58__19_, r_58__18_, r_58__17_, r_58__16_, r_58__15_, r_58__14_, r_58__13_, r_58__12_, r_58__11_, r_58__10_, r_58__9_, r_58__8_, r_58__7_, r_58__6_, r_58__5_, r_58__4_, r_58__3_, r_58__2_, r_58__1_, r_58__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N115)? data_i : 1'b0;
  assign N114 = sel_i[114];
  assign N115 = N1313;
  assign { r_n_58__63_, r_n_58__62_, r_n_58__61_, r_n_58__60_, r_n_58__59_, r_n_58__58_, r_n_58__57_, r_n_58__56_, r_n_58__55_, r_n_58__54_, r_n_58__53_, r_n_58__52_, r_n_58__51_, r_n_58__50_, r_n_58__49_, r_n_58__48_, r_n_58__47_, r_n_58__46_, r_n_58__45_, r_n_58__44_, r_n_58__43_, r_n_58__42_, r_n_58__41_, r_n_58__40_, r_n_58__39_, r_n_58__38_, r_n_58__37_, r_n_58__36_, r_n_58__35_, r_n_58__34_, r_n_58__33_, r_n_58__32_, r_n_58__31_, r_n_58__30_, r_n_58__29_, r_n_58__28_, r_n_58__27_, r_n_58__26_, r_n_58__25_, r_n_58__24_, r_n_58__23_, r_n_58__22_, r_n_58__21_, r_n_58__20_, r_n_58__19_, r_n_58__18_, r_n_58__17_, r_n_58__16_, r_n_58__15_, r_n_58__14_, r_n_58__13_, r_n_58__12_, r_n_58__11_, r_n_58__10_, r_n_58__9_, r_n_58__8_, r_n_58__7_, r_n_58__6_, r_n_58__5_, r_n_58__4_, r_n_58__3_, r_n_58__2_, r_n_58__1_, r_n_58__0_ } = (N116)? { r_59__63_, r_59__62_, r_59__61_, r_59__60_, r_59__59_, r_59__58_, r_59__57_, r_59__56_, r_59__55_, r_59__54_, r_59__53_, r_59__52_, r_59__51_, r_59__50_, r_59__49_, r_59__48_, r_59__47_, r_59__46_, r_59__45_, r_59__44_, r_59__43_, r_59__42_, r_59__41_, r_59__40_, r_59__39_, r_59__38_, r_59__37_, r_59__36_, r_59__35_, r_59__34_, r_59__33_, r_59__32_, r_59__31_, r_59__30_, r_59__29_, r_59__28_, r_59__27_, r_59__26_, r_59__25_, r_59__24_, r_59__23_, r_59__22_, r_59__21_, r_59__20_, r_59__19_, r_59__18_, r_59__17_, r_59__16_, r_59__15_, r_59__14_, r_59__13_, r_59__12_, r_59__11_, r_59__10_, r_59__9_, r_59__8_, r_59__7_, r_59__6_, r_59__5_, r_59__4_, r_59__3_, r_59__2_, r_59__1_, r_59__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N117)? data_i : 1'b0;
  assign N116 = sel_i[116];
  assign N117 = N1318;
  assign { r_n_59__63_, r_n_59__62_, r_n_59__61_, r_n_59__60_, r_n_59__59_, r_n_59__58_, r_n_59__57_, r_n_59__56_, r_n_59__55_, r_n_59__54_, r_n_59__53_, r_n_59__52_, r_n_59__51_, r_n_59__50_, r_n_59__49_, r_n_59__48_, r_n_59__47_, r_n_59__46_, r_n_59__45_, r_n_59__44_, r_n_59__43_, r_n_59__42_, r_n_59__41_, r_n_59__40_, r_n_59__39_, r_n_59__38_, r_n_59__37_, r_n_59__36_, r_n_59__35_, r_n_59__34_, r_n_59__33_, r_n_59__32_, r_n_59__31_, r_n_59__30_, r_n_59__29_, r_n_59__28_, r_n_59__27_, r_n_59__26_, r_n_59__25_, r_n_59__24_, r_n_59__23_, r_n_59__22_, r_n_59__21_, r_n_59__20_, r_n_59__19_, r_n_59__18_, r_n_59__17_, r_n_59__16_, r_n_59__15_, r_n_59__14_, r_n_59__13_, r_n_59__12_, r_n_59__11_, r_n_59__10_, r_n_59__9_, r_n_59__8_, r_n_59__7_, r_n_59__6_, r_n_59__5_, r_n_59__4_, r_n_59__3_, r_n_59__2_, r_n_59__1_, r_n_59__0_ } = (N118)? { r_60__63_, r_60__62_, r_60__61_, r_60__60_, r_60__59_, r_60__58_, r_60__57_, r_60__56_, r_60__55_, r_60__54_, r_60__53_, r_60__52_, r_60__51_, r_60__50_, r_60__49_, r_60__48_, r_60__47_, r_60__46_, r_60__45_, r_60__44_, r_60__43_, r_60__42_, r_60__41_, r_60__40_, r_60__39_, r_60__38_, r_60__37_, r_60__36_, r_60__35_, r_60__34_, r_60__33_, r_60__32_, r_60__31_, r_60__30_, r_60__29_, r_60__28_, r_60__27_, r_60__26_, r_60__25_, r_60__24_, r_60__23_, r_60__22_, r_60__21_, r_60__20_, r_60__19_, r_60__18_, r_60__17_, r_60__16_, r_60__15_, r_60__14_, r_60__13_, r_60__12_, r_60__11_, r_60__10_, r_60__9_, r_60__8_, r_60__7_, r_60__6_, r_60__5_, r_60__4_, r_60__3_, r_60__2_, r_60__1_, r_60__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N119)? data_i : 1'b0;
  assign N118 = sel_i[118];
  assign N119 = N1323;
  assign { r_n_60__63_, r_n_60__62_, r_n_60__61_, r_n_60__60_, r_n_60__59_, r_n_60__58_, r_n_60__57_, r_n_60__56_, r_n_60__55_, r_n_60__54_, r_n_60__53_, r_n_60__52_, r_n_60__51_, r_n_60__50_, r_n_60__49_, r_n_60__48_, r_n_60__47_, r_n_60__46_, r_n_60__45_, r_n_60__44_, r_n_60__43_, r_n_60__42_, r_n_60__41_, r_n_60__40_, r_n_60__39_, r_n_60__38_, r_n_60__37_, r_n_60__36_, r_n_60__35_, r_n_60__34_, r_n_60__33_, r_n_60__32_, r_n_60__31_, r_n_60__30_, r_n_60__29_, r_n_60__28_, r_n_60__27_, r_n_60__26_, r_n_60__25_, r_n_60__24_, r_n_60__23_, r_n_60__22_, r_n_60__21_, r_n_60__20_, r_n_60__19_, r_n_60__18_, r_n_60__17_, r_n_60__16_, r_n_60__15_, r_n_60__14_, r_n_60__13_, r_n_60__12_, r_n_60__11_, r_n_60__10_, r_n_60__9_, r_n_60__8_, r_n_60__7_, r_n_60__6_, r_n_60__5_, r_n_60__4_, r_n_60__3_, r_n_60__2_, r_n_60__1_, r_n_60__0_ } = (N120)? { r_61__63_, r_61__62_, r_61__61_, r_61__60_, r_61__59_, r_61__58_, r_61__57_, r_61__56_, r_61__55_, r_61__54_, r_61__53_, r_61__52_, r_61__51_, r_61__50_, r_61__49_, r_61__48_, r_61__47_, r_61__46_, r_61__45_, r_61__44_, r_61__43_, r_61__42_, r_61__41_, r_61__40_, r_61__39_, r_61__38_, r_61__37_, r_61__36_, r_61__35_, r_61__34_, r_61__33_, r_61__32_, r_61__31_, r_61__30_, r_61__29_, r_61__28_, r_61__27_, r_61__26_, r_61__25_, r_61__24_, r_61__23_, r_61__22_, r_61__21_, r_61__20_, r_61__19_, r_61__18_, r_61__17_, r_61__16_, r_61__15_, r_61__14_, r_61__13_, r_61__12_, r_61__11_, r_61__10_, r_61__9_, r_61__8_, r_61__7_, r_61__6_, r_61__5_, r_61__4_, r_61__3_, r_61__2_, r_61__1_, r_61__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N121)? data_i : 1'b0;
  assign N120 = sel_i[120];
  assign N121 = N1328;
  assign { r_n_61__63_, r_n_61__62_, r_n_61__61_, r_n_61__60_, r_n_61__59_, r_n_61__58_, r_n_61__57_, r_n_61__56_, r_n_61__55_, r_n_61__54_, r_n_61__53_, r_n_61__52_, r_n_61__51_, r_n_61__50_, r_n_61__49_, r_n_61__48_, r_n_61__47_, r_n_61__46_, r_n_61__45_, r_n_61__44_, r_n_61__43_, r_n_61__42_, r_n_61__41_, r_n_61__40_, r_n_61__39_, r_n_61__38_, r_n_61__37_, r_n_61__36_, r_n_61__35_, r_n_61__34_, r_n_61__33_, r_n_61__32_, r_n_61__31_, r_n_61__30_, r_n_61__29_, r_n_61__28_, r_n_61__27_, r_n_61__26_, r_n_61__25_, r_n_61__24_, r_n_61__23_, r_n_61__22_, r_n_61__21_, r_n_61__20_, r_n_61__19_, r_n_61__18_, r_n_61__17_, r_n_61__16_, r_n_61__15_, r_n_61__14_, r_n_61__13_, r_n_61__12_, r_n_61__11_, r_n_61__10_, r_n_61__9_, r_n_61__8_, r_n_61__7_, r_n_61__6_, r_n_61__5_, r_n_61__4_, r_n_61__3_, r_n_61__2_, r_n_61__1_, r_n_61__0_ } = (N122)? { r_62__63_, r_62__62_, r_62__61_, r_62__60_, r_62__59_, r_62__58_, r_62__57_, r_62__56_, r_62__55_, r_62__54_, r_62__53_, r_62__52_, r_62__51_, r_62__50_, r_62__49_, r_62__48_, r_62__47_, r_62__46_, r_62__45_, r_62__44_, r_62__43_, r_62__42_, r_62__41_, r_62__40_, r_62__39_, r_62__38_, r_62__37_, r_62__36_, r_62__35_, r_62__34_, r_62__33_, r_62__32_, r_62__31_, r_62__30_, r_62__29_, r_62__28_, r_62__27_, r_62__26_, r_62__25_, r_62__24_, r_62__23_, r_62__22_, r_62__21_, r_62__20_, r_62__19_, r_62__18_, r_62__17_, r_62__16_, r_62__15_, r_62__14_, r_62__13_, r_62__12_, r_62__11_, r_62__10_, r_62__9_, r_62__8_, r_62__7_, r_62__6_, r_62__5_, r_62__4_, r_62__3_, r_62__2_, r_62__1_, r_62__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N123)? data_i : 1'b0;
  assign N122 = sel_i[122];
  assign N123 = N1333;
  assign { r_n_62__63_, r_n_62__62_, r_n_62__61_, r_n_62__60_, r_n_62__59_, r_n_62__58_, r_n_62__57_, r_n_62__56_, r_n_62__55_, r_n_62__54_, r_n_62__53_, r_n_62__52_, r_n_62__51_, r_n_62__50_, r_n_62__49_, r_n_62__48_, r_n_62__47_, r_n_62__46_, r_n_62__45_, r_n_62__44_, r_n_62__43_, r_n_62__42_, r_n_62__41_, r_n_62__40_, r_n_62__39_, r_n_62__38_, r_n_62__37_, r_n_62__36_, r_n_62__35_, r_n_62__34_, r_n_62__33_, r_n_62__32_, r_n_62__31_, r_n_62__30_, r_n_62__29_, r_n_62__28_, r_n_62__27_, r_n_62__26_, r_n_62__25_, r_n_62__24_, r_n_62__23_, r_n_62__22_, r_n_62__21_, r_n_62__20_, r_n_62__19_, r_n_62__18_, r_n_62__17_, r_n_62__16_, r_n_62__15_, r_n_62__14_, r_n_62__13_, r_n_62__12_, r_n_62__11_, r_n_62__10_, r_n_62__9_, r_n_62__8_, r_n_62__7_, r_n_62__6_, r_n_62__5_, r_n_62__4_, r_n_62__3_, r_n_62__2_, r_n_62__1_, r_n_62__0_ } = (N124)? { r_63__63_, r_63__62_, r_63__61_, r_63__60_, r_63__59_, r_63__58_, r_63__57_, r_63__56_, r_63__55_, r_63__54_, r_63__53_, r_63__52_, r_63__51_, r_63__50_, r_63__49_, r_63__48_, r_63__47_, r_63__46_, r_63__45_, r_63__44_, r_63__43_, r_63__42_, r_63__41_, r_63__40_, r_63__39_, r_63__38_, r_63__37_, r_63__36_, r_63__35_, r_63__34_, r_63__33_, r_63__32_, r_63__31_, r_63__30_, r_63__29_, r_63__28_, r_63__27_, r_63__26_, r_63__25_, r_63__24_, r_63__23_, r_63__22_, r_63__21_, r_63__20_, r_63__19_, r_63__18_, r_63__17_, r_63__16_, r_63__15_, r_63__14_, r_63__13_, r_63__12_, r_63__11_, r_63__10_, r_63__9_, r_63__8_, r_63__7_, r_63__6_, r_63__5_, r_63__4_, r_63__3_, r_63__2_, r_63__1_, r_63__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N125)? data_i : 1'b0;
  assign N124 = sel_i[124];
  assign N125 = N1338;
  assign { r_n_63__63_, r_n_63__62_, r_n_63__61_, r_n_63__60_, r_n_63__59_, r_n_63__58_, r_n_63__57_, r_n_63__56_, r_n_63__55_, r_n_63__54_, r_n_63__53_, r_n_63__52_, r_n_63__51_, r_n_63__50_, r_n_63__49_, r_n_63__48_, r_n_63__47_, r_n_63__46_, r_n_63__45_, r_n_63__44_, r_n_63__43_, r_n_63__42_, r_n_63__41_, r_n_63__40_, r_n_63__39_, r_n_63__38_, r_n_63__37_, r_n_63__36_, r_n_63__35_, r_n_63__34_, r_n_63__33_, r_n_63__32_, r_n_63__31_, r_n_63__30_, r_n_63__29_, r_n_63__28_, r_n_63__27_, r_n_63__26_, r_n_63__25_, r_n_63__24_, r_n_63__23_, r_n_63__22_, r_n_63__21_, r_n_63__20_, r_n_63__19_, r_n_63__18_, r_n_63__17_, r_n_63__16_, r_n_63__15_, r_n_63__14_, r_n_63__13_, r_n_63__12_, r_n_63__11_, r_n_63__10_, r_n_63__9_, r_n_63__8_, r_n_63__7_, r_n_63__6_, r_n_63__5_, r_n_63__4_, r_n_63__3_, r_n_63__2_, r_n_63__1_, r_n_63__0_ } = (N126)? { r_64__63_, r_64__62_, r_64__61_, r_64__60_, r_64__59_, r_64__58_, r_64__57_, r_64__56_, r_64__55_, r_64__54_, r_64__53_, r_64__52_, r_64__51_, r_64__50_, r_64__49_, r_64__48_, r_64__47_, r_64__46_, r_64__45_, r_64__44_, r_64__43_, r_64__42_, r_64__41_, r_64__40_, r_64__39_, r_64__38_, r_64__37_, r_64__36_, r_64__35_, r_64__34_, r_64__33_, r_64__32_, r_64__31_, r_64__30_, r_64__29_, r_64__28_, r_64__27_, r_64__26_, r_64__25_, r_64__24_, r_64__23_, r_64__22_, r_64__21_, r_64__20_, r_64__19_, r_64__18_, r_64__17_, r_64__16_, r_64__15_, r_64__14_, r_64__13_, r_64__12_, r_64__11_, r_64__10_, r_64__9_, r_64__8_, r_64__7_, r_64__6_, r_64__5_, r_64__4_, r_64__3_, r_64__2_, r_64__1_, r_64__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N127)? data_i : 1'b0;
  assign N126 = sel_i[126];
  assign N127 = N1343;
  assign { r_n_64__63_, r_n_64__62_, r_n_64__61_, r_n_64__60_, r_n_64__59_, r_n_64__58_, r_n_64__57_, r_n_64__56_, r_n_64__55_, r_n_64__54_, r_n_64__53_, r_n_64__52_, r_n_64__51_, r_n_64__50_, r_n_64__49_, r_n_64__48_, r_n_64__47_, r_n_64__46_, r_n_64__45_, r_n_64__44_, r_n_64__43_, r_n_64__42_, r_n_64__41_, r_n_64__40_, r_n_64__39_, r_n_64__38_, r_n_64__37_, r_n_64__36_, r_n_64__35_, r_n_64__34_, r_n_64__33_, r_n_64__32_, r_n_64__31_, r_n_64__30_, r_n_64__29_, r_n_64__28_, r_n_64__27_, r_n_64__26_, r_n_64__25_, r_n_64__24_, r_n_64__23_, r_n_64__22_, r_n_64__21_, r_n_64__20_, r_n_64__19_, r_n_64__18_, r_n_64__17_, r_n_64__16_, r_n_64__15_, r_n_64__14_, r_n_64__13_, r_n_64__12_, r_n_64__11_, r_n_64__10_, r_n_64__9_, r_n_64__8_, r_n_64__7_, r_n_64__6_, r_n_64__5_, r_n_64__4_, r_n_64__3_, r_n_64__2_, r_n_64__1_, r_n_64__0_ } = (N128)? { r_65__63_, r_65__62_, r_65__61_, r_65__60_, r_65__59_, r_65__58_, r_65__57_, r_65__56_, r_65__55_, r_65__54_, r_65__53_, r_65__52_, r_65__51_, r_65__50_, r_65__49_, r_65__48_, r_65__47_, r_65__46_, r_65__45_, r_65__44_, r_65__43_, r_65__42_, r_65__41_, r_65__40_, r_65__39_, r_65__38_, r_65__37_, r_65__36_, r_65__35_, r_65__34_, r_65__33_, r_65__32_, r_65__31_, r_65__30_, r_65__29_, r_65__28_, r_65__27_, r_65__26_, r_65__25_, r_65__24_, r_65__23_, r_65__22_, r_65__21_, r_65__20_, r_65__19_, r_65__18_, r_65__17_, r_65__16_, r_65__15_, r_65__14_, r_65__13_, r_65__12_, r_65__11_, r_65__10_, r_65__9_, r_65__8_, r_65__7_, r_65__6_, r_65__5_, r_65__4_, r_65__3_, r_65__2_, r_65__1_, r_65__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N129)? data_i : 1'b0;
  assign N128 = sel_i[128];
  assign N129 = N1348;
  assign { r_n_65__63_, r_n_65__62_, r_n_65__61_, r_n_65__60_, r_n_65__59_, r_n_65__58_, r_n_65__57_, r_n_65__56_, r_n_65__55_, r_n_65__54_, r_n_65__53_, r_n_65__52_, r_n_65__51_, r_n_65__50_, r_n_65__49_, r_n_65__48_, r_n_65__47_, r_n_65__46_, r_n_65__45_, r_n_65__44_, r_n_65__43_, r_n_65__42_, r_n_65__41_, r_n_65__40_, r_n_65__39_, r_n_65__38_, r_n_65__37_, r_n_65__36_, r_n_65__35_, r_n_65__34_, r_n_65__33_, r_n_65__32_, r_n_65__31_, r_n_65__30_, r_n_65__29_, r_n_65__28_, r_n_65__27_, r_n_65__26_, r_n_65__25_, r_n_65__24_, r_n_65__23_, r_n_65__22_, r_n_65__21_, r_n_65__20_, r_n_65__19_, r_n_65__18_, r_n_65__17_, r_n_65__16_, r_n_65__15_, r_n_65__14_, r_n_65__13_, r_n_65__12_, r_n_65__11_, r_n_65__10_, r_n_65__9_, r_n_65__8_, r_n_65__7_, r_n_65__6_, r_n_65__5_, r_n_65__4_, r_n_65__3_, r_n_65__2_, r_n_65__1_, r_n_65__0_ } = (N130)? { r_66__63_, r_66__62_, r_66__61_, r_66__60_, r_66__59_, r_66__58_, r_66__57_, r_66__56_, r_66__55_, r_66__54_, r_66__53_, r_66__52_, r_66__51_, r_66__50_, r_66__49_, r_66__48_, r_66__47_, r_66__46_, r_66__45_, r_66__44_, r_66__43_, r_66__42_, r_66__41_, r_66__40_, r_66__39_, r_66__38_, r_66__37_, r_66__36_, r_66__35_, r_66__34_, r_66__33_, r_66__32_, r_66__31_, r_66__30_, r_66__29_, r_66__28_, r_66__27_, r_66__26_, r_66__25_, r_66__24_, r_66__23_, r_66__22_, r_66__21_, r_66__20_, r_66__19_, r_66__18_, r_66__17_, r_66__16_, r_66__15_, r_66__14_, r_66__13_, r_66__12_, r_66__11_, r_66__10_, r_66__9_, r_66__8_, r_66__7_, r_66__6_, r_66__5_, r_66__4_, r_66__3_, r_66__2_, r_66__1_, r_66__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N131)? data_i : 1'b0;
  assign N130 = sel_i[130];
  assign N131 = N1353;
  assign { r_n_66__63_, r_n_66__62_, r_n_66__61_, r_n_66__60_, r_n_66__59_, r_n_66__58_, r_n_66__57_, r_n_66__56_, r_n_66__55_, r_n_66__54_, r_n_66__53_, r_n_66__52_, r_n_66__51_, r_n_66__50_, r_n_66__49_, r_n_66__48_, r_n_66__47_, r_n_66__46_, r_n_66__45_, r_n_66__44_, r_n_66__43_, r_n_66__42_, r_n_66__41_, r_n_66__40_, r_n_66__39_, r_n_66__38_, r_n_66__37_, r_n_66__36_, r_n_66__35_, r_n_66__34_, r_n_66__33_, r_n_66__32_, r_n_66__31_, r_n_66__30_, r_n_66__29_, r_n_66__28_, r_n_66__27_, r_n_66__26_, r_n_66__25_, r_n_66__24_, r_n_66__23_, r_n_66__22_, r_n_66__21_, r_n_66__20_, r_n_66__19_, r_n_66__18_, r_n_66__17_, r_n_66__16_, r_n_66__15_, r_n_66__14_, r_n_66__13_, r_n_66__12_, r_n_66__11_, r_n_66__10_, r_n_66__9_, r_n_66__8_, r_n_66__7_, r_n_66__6_, r_n_66__5_, r_n_66__4_, r_n_66__3_, r_n_66__2_, r_n_66__1_, r_n_66__0_ } = (N132)? { r_67__63_, r_67__62_, r_67__61_, r_67__60_, r_67__59_, r_67__58_, r_67__57_, r_67__56_, r_67__55_, r_67__54_, r_67__53_, r_67__52_, r_67__51_, r_67__50_, r_67__49_, r_67__48_, r_67__47_, r_67__46_, r_67__45_, r_67__44_, r_67__43_, r_67__42_, r_67__41_, r_67__40_, r_67__39_, r_67__38_, r_67__37_, r_67__36_, r_67__35_, r_67__34_, r_67__33_, r_67__32_, r_67__31_, r_67__30_, r_67__29_, r_67__28_, r_67__27_, r_67__26_, r_67__25_, r_67__24_, r_67__23_, r_67__22_, r_67__21_, r_67__20_, r_67__19_, r_67__18_, r_67__17_, r_67__16_, r_67__15_, r_67__14_, r_67__13_, r_67__12_, r_67__11_, r_67__10_, r_67__9_, r_67__8_, r_67__7_, r_67__6_, r_67__5_, r_67__4_, r_67__3_, r_67__2_, r_67__1_, r_67__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N133)? data_i : 1'b0;
  assign N132 = sel_i[132];
  assign N133 = N1358;
  assign { r_n_67__63_, r_n_67__62_, r_n_67__61_, r_n_67__60_, r_n_67__59_, r_n_67__58_, r_n_67__57_, r_n_67__56_, r_n_67__55_, r_n_67__54_, r_n_67__53_, r_n_67__52_, r_n_67__51_, r_n_67__50_, r_n_67__49_, r_n_67__48_, r_n_67__47_, r_n_67__46_, r_n_67__45_, r_n_67__44_, r_n_67__43_, r_n_67__42_, r_n_67__41_, r_n_67__40_, r_n_67__39_, r_n_67__38_, r_n_67__37_, r_n_67__36_, r_n_67__35_, r_n_67__34_, r_n_67__33_, r_n_67__32_, r_n_67__31_, r_n_67__30_, r_n_67__29_, r_n_67__28_, r_n_67__27_, r_n_67__26_, r_n_67__25_, r_n_67__24_, r_n_67__23_, r_n_67__22_, r_n_67__21_, r_n_67__20_, r_n_67__19_, r_n_67__18_, r_n_67__17_, r_n_67__16_, r_n_67__15_, r_n_67__14_, r_n_67__13_, r_n_67__12_, r_n_67__11_, r_n_67__10_, r_n_67__9_, r_n_67__8_, r_n_67__7_, r_n_67__6_, r_n_67__5_, r_n_67__4_, r_n_67__3_, r_n_67__2_, r_n_67__1_, r_n_67__0_ } = (N134)? { r_68__63_, r_68__62_, r_68__61_, r_68__60_, r_68__59_, r_68__58_, r_68__57_, r_68__56_, r_68__55_, r_68__54_, r_68__53_, r_68__52_, r_68__51_, r_68__50_, r_68__49_, r_68__48_, r_68__47_, r_68__46_, r_68__45_, r_68__44_, r_68__43_, r_68__42_, r_68__41_, r_68__40_, r_68__39_, r_68__38_, r_68__37_, r_68__36_, r_68__35_, r_68__34_, r_68__33_, r_68__32_, r_68__31_, r_68__30_, r_68__29_, r_68__28_, r_68__27_, r_68__26_, r_68__25_, r_68__24_, r_68__23_, r_68__22_, r_68__21_, r_68__20_, r_68__19_, r_68__18_, r_68__17_, r_68__16_, r_68__15_, r_68__14_, r_68__13_, r_68__12_, r_68__11_, r_68__10_, r_68__9_, r_68__8_, r_68__7_, r_68__6_, r_68__5_, r_68__4_, r_68__3_, r_68__2_, r_68__1_, r_68__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N135)? data_i : 1'b0;
  assign N134 = sel_i[134];
  assign N135 = N1363;
  assign { r_n_68__63_, r_n_68__62_, r_n_68__61_, r_n_68__60_, r_n_68__59_, r_n_68__58_, r_n_68__57_, r_n_68__56_, r_n_68__55_, r_n_68__54_, r_n_68__53_, r_n_68__52_, r_n_68__51_, r_n_68__50_, r_n_68__49_, r_n_68__48_, r_n_68__47_, r_n_68__46_, r_n_68__45_, r_n_68__44_, r_n_68__43_, r_n_68__42_, r_n_68__41_, r_n_68__40_, r_n_68__39_, r_n_68__38_, r_n_68__37_, r_n_68__36_, r_n_68__35_, r_n_68__34_, r_n_68__33_, r_n_68__32_, r_n_68__31_, r_n_68__30_, r_n_68__29_, r_n_68__28_, r_n_68__27_, r_n_68__26_, r_n_68__25_, r_n_68__24_, r_n_68__23_, r_n_68__22_, r_n_68__21_, r_n_68__20_, r_n_68__19_, r_n_68__18_, r_n_68__17_, r_n_68__16_, r_n_68__15_, r_n_68__14_, r_n_68__13_, r_n_68__12_, r_n_68__11_, r_n_68__10_, r_n_68__9_, r_n_68__8_, r_n_68__7_, r_n_68__6_, r_n_68__5_, r_n_68__4_, r_n_68__3_, r_n_68__2_, r_n_68__1_, r_n_68__0_ } = (N136)? { r_69__63_, r_69__62_, r_69__61_, r_69__60_, r_69__59_, r_69__58_, r_69__57_, r_69__56_, r_69__55_, r_69__54_, r_69__53_, r_69__52_, r_69__51_, r_69__50_, r_69__49_, r_69__48_, r_69__47_, r_69__46_, r_69__45_, r_69__44_, r_69__43_, r_69__42_, r_69__41_, r_69__40_, r_69__39_, r_69__38_, r_69__37_, r_69__36_, r_69__35_, r_69__34_, r_69__33_, r_69__32_, r_69__31_, r_69__30_, r_69__29_, r_69__28_, r_69__27_, r_69__26_, r_69__25_, r_69__24_, r_69__23_, r_69__22_, r_69__21_, r_69__20_, r_69__19_, r_69__18_, r_69__17_, r_69__16_, r_69__15_, r_69__14_, r_69__13_, r_69__12_, r_69__11_, r_69__10_, r_69__9_, r_69__8_, r_69__7_, r_69__6_, r_69__5_, r_69__4_, r_69__3_, r_69__2_, r_69__1_, r_69__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N137)? data_i : 1'b0;
  assign N136 = sel_i[136];
  assign N137 = N1368;
  assign { r_n_69__63_, r_n_69__62_, r_n_69__61_, r_n_69__60_, r_n_69__59_, r_n_69__58_, r_n_69__57_, r_n_69__56_, r_n_69__55_, r_n_69__54_, r_n_69__53_, r_n_69__52_, r_n_69__51_, r_n_69__50_, r_n_69__49_, r_n_69__48_, r_n_69__47_, r_n_69__46_, r_n_69__45_, r_n_69__44_, r_n_69__43_, r_n_69__42_, r_n_69__41_, r_n_69__40_, r_n_69__39_, r_n_69__38_, r_n_69__37_, r_n_69__36_, r_n_69__35_, r_n_69__34_, r_n_69__33_, r_n_69__32_, r_n_69__31_, r_n_69__30_, r_n_69__29_, r_n_69__28_, r_n_69__27_, r_n_69__26_, r_n_69__25_, r_n_69__24_, r_n_69__23_, r_n_69__22_, r_n_69__21_, r_n_69__20_, r_n_69__19_, r_n_69__18_, r_n_69__17_, r_n_69__16_, r_n_69__15_, r_n_69__14_, r_n_69__13_, r_n_69__12_, r_n_69__11_, r_n_69__10_, r_n_69__9_, r_n_69__8_, r_n_69__7_, r_n_69__6_, r_n_69__5_, r_n_69__4_, r_n_69__3_, r_n_69__2_, r_n_69__1_, r_n_69__0_ } = (N138)? { r_70__63_, r_70__62_, r_70__61_, r_70__60_, r_70__59_, r_70__58_, r_70__57_, r_70__56_, r_70__55_, r_70__54_, r_70__53_, r_70__52_, r_70__51_, r_70__50_, r_70__49_, r_70__48_, r_70__47_, r_70__46_, r_70__45_, r_70__44_, r_70__43_, r_70__42_, r_70__41_, r_70__40_, r_70__39_, r_70__38_, r_70__37_, r_70__36_, r_70__35_, r_70__34_, r_70__33_, r_70__32_, r_70__31_, r_70__30_, r_70__29_, r_70__28_, r_70__27_, r_70__26_, r_70__25_, r_70__24_, r_70__23_, r_70__22_, r_70__21_, r_70__20_, r_70__19_, r_70__18_, r_70__17_, r_70__16_, r_70__15_, r_70__14_, r_70__13_, r_70__12_, r_70__11_, r_70__10_, r_70__9_, r_70__8_, r_70__7_, r_70__6_, r_70__5_, r_70__4_, r_70__3_, r_70__2_, r_70__1_, r_70__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N139)? data_i : 1'b0;
  assign N138 = sel_i[138];
  assign N139 = N1373;
  assign { r_n_70__63_, r_n_70__62_, r_n_70__61_, r_n_70__60_, r_n_70__59_, r_n_70__58_, r_n_70__57_, r_n_70__56_, r_n_70__55_, r_n_70__54_, r_n_70__53_, r_n_70__52_, r_n_70__51_, r_n_70__50_, r_n_70__49_, r_n_70__48_, r_n_70__47_, r_n_70__46_, r_n_70__45_, r_n_70__44_, r_n_70__43_, r_n_70__42_, r_n_70__41_, r_n_70__40_, r_n_70__39_, r_n_70__38_, r_n_70__37_, r_n_70__36_, r_n_70__35_, r_n_70__34_, r_n_70__33_, r_n_70__32_, r_n_70__31_, r_n_70__30_, r_n_70__29_, r_n_70__28_, r_n_70__27_, r_n_70__26_, r_n_70__25_, r_n_70__24_, r_n_70__23_, r_n_70__22_, r_n_70__21_, r_n_70__20_, r_n_70__19_, r_n_70__18_, r_n_70__17_, r_n_70__16_, r_n_70__15_, r_n_70__14_, r_n_70__13_, r_n_70__12_, r_n_70__11_, r_n_70__10_, r_n_70__9_, r_n_70__8_, r_n_70__7_, r_n_70__6_, r_n_70__5_, r_n_70__4_, r_n_70__3_, r_n_70__2_, r_n_70__1_, r_n_70__0_ } = (N140)? { r_71__63_, r_71__62_, r_71__61_, r_71__60_, r_71__59_, r_71__58_, r_71__57_, r_71__56_, r_71__55_, r_71__54_, r_71__53_, r_71__52_, r_71__51_, r_71__50_, r_71__49_, r_71__48_, r_71__47_, r_71__46_, r_71__45_, r_71__44_, r_71__43_, r_71__42_, r_71__41_, r_71__40_, r_71__39_, r_71__38_, r_71__37_, r_71__36_, r_71__35_, r_71__34_, r_71__33_, r_71__32_, r_71__31_, r_71__30_, r_71__29_, r_71__28_, r_71__27_, r_71__26_, r_71__25_, r_71__24_, r_71__23_, r_71__22_, r_71__21_, r_71__20_, r_71__19_, r_71__18_, r_71__17_, r_71__16_, r_71__15_, r_71__14_, r_71__13_, r_71__12_, r_71__11_, r_71__10_, r_71__9_, r_71__8_, r_71__7_, r_71__6_, r_71__5_, r_71__4_, r_71__3_, r_71__2_, r_71__1_, r_71__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N141)? data_i : 1'b0;
  assign N140 = sel_i[140];
  assign N141 = N1378;
  assign { r_n_71__63_, r_n_71__62_, r_n_71__61_, r_n_71__60_, r_n_71__59_, r_n_71__58_, r_n_71__57_, r_n_71__56_, r_n_71__55_, r_n_71__54_, r_n_71__53_, r_n_71__52_, r_n_71__51_, r_n_71__50_, r_n_71__49_, r_n_71__48_, r_n_71__47_, r_n_71__46_, r_n_71__45_, r_n_71__44_, r_n_71__43_, r_n_71__42_, r_n_71__41_, r_n_71__40_, r_n_71__39_, r_n_71__38_, r_n_71__37_, r_n_71__36_, r_n_71__35_, r_n_71__34_, r_n_71__33_, r_n_71__32_, r_n_71__31_, r_n_71__30_, r_n_71__29_, r_n_71__28_, r_n_71__27_, r_n_71__26_, r_n_71__25_, r_n_71__24_, r_n_71__23_, r_n_71__22_, r_n_71__21_, r_n_71__20_, r_n_71__19_, r_n_71__18_, r_n_71__17_, r_n_71__16_, r_n_71__15_, r_n_71__14_, r_n_71__13_, r_n_71__12_, r_n_71__11_, r_n_71__10_, r_n_71__9_, r_n_71__8_, r_n_71__7_, r_n_71__6_, r_n_71__5_, r_n_71__4_, r_n_71__3_, r_n_71__2_, r_n_71__1_, r_n_71__0_ } = (N142)? { r_72__63_, r_72__62_, r_72__61_, r_72__60_, r_72__59_, r_72__58_, r_72__57_, r_72__56_, r_72__55_, r_72__54_, r_72__53_, r_72__52_, r_72__51_, r_72__50_, r_72__49_, r_72__48_, r_72__47_, r_72__46_, r_72__45_, r_72__44_, r_72__43_, r_72__42_, r_72__41_, r_72__40_, r_72__39_, r_72__38_, r_72__37_, r_72__36_, r_72__35_, r_72__34_, r_72__33_, r_72__32_, r_72__31_, r_72__30_, r_72__29_, r_72__28_, r_72__27_, r_72__26_, r_72__25_, r_72__24_, r_72__23_, r_72__22_, r_72__21_, r_72__20_, r_72__19_, r_72__18_, r_72__17_, r_72__16_, r_72__15_, r_72__14_, r_72__13_, r_72__12_, r_72__11_, r_72__10_, r_72__9_, r_72__8_, r_72__7_, r_72__6_, r_72__5_, r_72__4_, r_72__3_, r_72__2_, r_72__1_, r_72__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N143)? data_i : 1'b0;
  assign N142 = sel_i[142];
  assign N143 = N1383;
  assign { r_n_72__63_, r_n_72__62_, r_n_72__61_, r_n_72__60_, r_n_72__59_, r_n_72__58_, r_n_72__57_, r_n_72__56_, r_n_72__55_, r_n_72__54_, r_n_72__53_, r_n_72__52_, r_n_72__51_, r_n_72__50_, r_n_72__49_, r_n_72__48_, r_n_72__47_, r_n_72__46_, r_n_72__45_, r_n_72__44_, r_n_72__43_, r_n_72__42_, r_n_72__41_, r_n_72__40_, r_n_72__39_, r_n_72__38_, r_n_72__37_, r_n_72__36_, r_n_72__35_, r_n_72__34_, r_n_72__33_, r_n_72__32_, r_n_72__31_, r_n_72__30_, r_n_72__29_, r_n_72__28_, r_n_72__27_, r_n_72__26_, r_n_72__25_, r_n_72__24_, r_n_72__23_, r_n_72__22_, r_n_72__21_, r_n_72__20_, r_n_72__19_, r_n_72__18_, r_n_72__17_, r_n_72__16_, r_n_72__15_, r_n_72__14_, r_n_72__13_, r_n_72__12_, r_n_72__11_, r_n_72__10_, r_n_72__9_, r_n_72__8_, r_n_72__7_, r_n_72__6_, r_n_72__5_, r_n_72__4_, r_n_72__3_, r_n_72__2_, r_n_72__1_, r_n_72__0_ } = (N144)? { r_73__63_, r_73__62_, r_73__61_, r_73__60_, r_73__59_, r_73__58_, r_73__57_, r_73__56_, r_73__55_, r_73__54_, r_73__53_, r_73__52_, r_73__51_, r_73__50_, r_73__49_, r_73__48_, r_73__47_, r_73__46_, r_73__45_, r_73__44_, r_73__43_, r_73__42_, r_73__41_, r_73__40_, r_73__39_, r_73__38_, r_73__37_, r_73__36_, r_73__35_, r_73__34_, r_73__33_, r_73__32_, r_73__31_, r_73__30_, r_73__29_, r_73__28_, r_73__27_, r_73__26_, r_73__25_, r_73__24_, r_73__23_, r_73__22_, r_73__21_, r_73__20_, r_73__19_, r_73__18_, r_73__17_, r_73__16_, r_73__15_, r_73__14_, r_73__13_, r_73__12_, r_73__11_, r_73__10_, r_73__9_, r_73__8_, r_73__7_, r_73__6_, r_73__5_, r_73__4_, r_73__3_, r_73__2_, r_73__1_, r_73__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N145)? data_i : 1'b0;
  assign N144 = sel_i[144];
  assign N145 = N1388;
  assign { r_n_73__63_, r_n_73__62_, r_n_73__61_, r_n_73__60_, r_n_73__59_, r_n_73__58_, r_n_73__57_, r_n_73__56_, r_n_73__55_, r_n_73__54_, r_n_73__53_, r_n_73__52_, r_n_73__51_, r_n_73__50_, r_n_73__49_, r_n_73__48_, r_n_73__47_, r_n_73__46_, r_n_73__45_, r_n_73__44_, r_n_73__43_, r_n_73__42_, r_n_73__41_, r_n_73__40_, r_n_73__39_, r_n_73__38_, r_n_73__37_, r_n_73__36_, r_n_73__35_, r_n_73__34_, r_n_73__33_, r_n_73__32_, r_n_73__31_, r_n_73__30_, r_n_73__29_, r_n_73__28_, r_n_73__27_, r_n_73__26_, r_n_73__25_, r_n_73__24_, r_n_73__23_, r_n_73__22_, r_n_73__21_, r_n_73__20_, r_n_73__19_, r_n_73__18_, r_n_73__17_, r_n_73__16_, r_n_73__15_, r_n_73__14_, r_n_73__13_, r_n_73__12_, r_n_73__11_, r_n_73__10_, r_n_73__9_, r_n_73__8_, r_n_73__7_, r_n_73__6_, r_n_73__5_, r_n_73__4_, r_n_73__3_, r_n_73__2_, r_n_73__1_, r_n_73__0_ } = (N146)? { r_74__63_, r_74__62_, r_74__61_, r_74__60_, r_74__59_, r_74__58_, r_74__57_, r_74__56_, r_74__55_, r_74__54_, r_74__53_, r_74__52_, r_74__51_, r_74__50_, r_74__49_, r_74__48_, r_74__47_, r_74__46_, r_74__45_, r_74__44_, r_74__43_, r_74__42_, r_74__41_, r_74__40_, r_74__39_, r_74__38_, r_74__37_, r_74__36_, r_74__35_, r_74__34_, r_74__33_, r_74__32_, r_74__31_, r_74__30_, r_74__29_, r_74__28_, r_74__27_, r_74__26_, r_74__25_, r_74__24_, r_74__23_, r_74__22_, r_74__21_, r_74__20_, r_74__19_, r_74__18_, r_74__17_, r_74__16_, r_74__15_, r_74__14_, r_74__13_, r_74__12_, r_74__11_, r_74__10_, r_74__9_, r_74__8_, r_74__7_, r_74__6_, r_74__5_, r_74__4_, r_74__3_, r_74__2_, r_74__1_, r_74__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N147)? data_i : 1'b0;
  assign N146 = sel_i[146];
  assign N147 = N1393;
  assign { r_n_74__63_, r_n_74__62_, r_n_74__61_, r_n_74__60_, r_n_74__59_, r_n_74__58_, r_n_74__57_, r_n_74__56_, r_n_74__55_, r_n_74__54_, r_n_74__53_, r_n_74__52_, r_n_74__51_, r_n_74__50_, r_n_74__49_, r_n_74__48_, r_n_74__47_, r_n_74__46_, r_n_74__45_, r_n_74__44_, r_n_74__43_, r_n_74__42_, r_n_74__41_, r_n_74__40_, r_n_74__39_, r_n_74__38_, r_n_74__37_, r_n_74__36_, r_n_74__35_, r_n_74__34_, r_n_74__33_, r_n_74__32_, r_n_74__31_, r_n_74__30_, r_n_74__29_, r_n_74__28_, r_n_74__27_, r_n_74__26_, r_n_74__25_, r_n_74__24_, r_n_74__23_, r_n_74__22_, r_n_74__21_, r_n_74__20_, r_n_74__19_, r_n_74__18_, r_n_74__17_, r_n_74__16_, r_n_74__15_, r_n_74__14_, r_n_74__13_, r_n_74__12_, r_n_74__11_, r_n_74__10_, r_n_74__9_, r_n_74__8_, r_n_74__7_, r_n_74__6_, r_n_74__5_, r_n_74__4_, r_n_74__3_, r_n_74__2_, r_n_74__1_, r_n_74__0_ } = (N148)? { r_75__63_, r_75__62_, r_75__61_, r_75__60_, r_75__59_, r_75__58_, r_75__57_, r_75__56_, r_75__55_, r_75__54_, r_75__53_, r_75__52_, r_75__51_, r_75__50_, r_75__49_, r_75__48_, r_75__47_, r_75__46_, r_75__45_, r_75__44_, r_75__43_, r_75__42_, r_75__41_, r_75__40_, r_75__39_, r_75__38_, r_75__37_, r_75__36_, r_75__35_, r_75__34_, r_75__33_, r_75__32_, r_75__31_, r_75__30_, r_75__29_, r_75__28_, r_75__27_, r_75__26_, r_75__25_, r_75__24_, r_75__23_, r_75__22_, r_75__21_, r_75__20_, r_75__19_, r_75__18_, r_75__17_, r_75__16_, r_75__15_, r_75__14_, r_75__13_, r_75__12_, r_75__11_, r_75__10_, r_75__9_, r_75__8_, r_75__7_, r_75__6_, r_75__5_, r_75__4_, r_75__3_, r_75__2_, r_75__1_, r_75__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N149)? data_i : 1'b0;
  assign N148 = sel_i[148];
  assign N149 = N1398;
  assign { r_n_75__63_, r_n_75__62_, r_n_75__61_, r_n_75__60_, r_n_75__59_, r_n_75__58_, r_n_75__57_, r_n_75__56_, r_n_75__55_, r_n_75__54_, r_n_75__53_, r_n_75__52_, r_n_75__51_, r_n_75__50_, r_n_75__49_, r_n_75__48_, r_n_75__47_, r_n_75__46_, r_n_75__45_, r_n_75__44_, r_n_75__43_, r_n_75__42_, r_n_75__41_, r_n_75__40_, r_n_75__39_, r_n_75__38_, r_n_75__37_, r_n_75__36_, r_n_75__35_, r_n_75__34_, r_n_75__33_, r_n_75__32_, r_n_75__31_, r_n_75__30_, r_n_75__29_, r_n_75__28_, r_n_75__27_, r_n_75__26_, r_n_75__25_, r_n_75__24_, r_n_75__23_, r_n_75__22_, r_n_75__21_, r_n_75__20_, r_n_75__19_, r_n_75__18_, r_n_75__17_, r_n_75__16_, r_n_75__15_, r_n_75__14_, r_n_75__13_, r_n_75__12_, r_n_75__11_, r_n_75__10_, r_n_75__9_, r_n_75__8_, r_n_75__7_, r_n_75__6_, r_n_75__5_, r_n_75__4_, r_n_75__3_, r_n_75__2_, r_n_75__1_, r_n_75__0_ } = (N150)? { r_76__63_, r_76__62_, r_76__61_, r_76__60_, r_76__59_, r_76__58_, r_76__57_, r_76__56_, r_76__55_, r_76__54_, r_76__53_, r_76__52_, r_76__51_, r_76__50_, r_76__49_, r_76__48_, r_76__47_, r_76__46_, r_76__45_, r_76__44_, r_76__43_, r_76__42_, r_76__41_, r_76__40_, r_76__39_, r_76__38_, r_76__37_, r_76__36_, r_76__35_, r_76__34_, r_76__33_, r_76__32_, r_76__31_, r_76__30_, r_76__29_, r_76__28_, r_76__27_, r_76__26_, r_76__25_, r_76__24_, r_76__23_, r_76__22_, r_76__21_, r_76__20_, r_76__19_, r_76__18_, r_76__17_, r_76__16_, r_76__15_, r_76__14_, r_76__13_, r_76__12_, r_76__11_, r_76__10_, r_76__9_, r_76__8_, r_76__7_, r_76__6_, r_76__5_, r_76__4_, r_76__3_, r_76__2_, r_76__1_, r_76__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N151)? data_i : 1'b0;
  assign N150 = sel_i[150];
  assign N151 = N1403;
  assign { r_n_76__63_, r_n_76__62_, r_n_76__61_, r_n_76__60_, r_n_76__59_, r_n_76__58_, r_n_76__57_, r_n_76__56_, r_n_76__55_, r_n_76__54_, r_n_76__53_, r_n_76__52_, r_n_76__51_, r_n_76__50_, r_n_76__49_, r_n_76__48_, r_n_76__47_, r_n_76__46_, r_n_76__45_, r_n_76__44_, r_n_76__43_, r_n_76__42_, r_n_76__41_, r_n_76__40_, r_n_76__39_, r_n_76__38_, r_n_76__37_, r_n_76__36_, r_n_76__35_, r_n_76__34_, r_n_76__33_, r_n_76__32_, r_n_76__31_, r_n_76__30_, r_n_76__29_, r_n_76__28_, r_n_76__27_, r_n_76__26_, r_n_76__25_, r_n_76__24_, r_n_76__23_, r_n_76__22_, r_n_76__21_, r_n_76__20_, r_n_76__19_, r_n_76__18_, r_n_76__17_, r_n_76__16_, r_n_76__15_, r_n_76__14_, r_n_76__13_, r_n_76__12_, r_n_76__11_, r_n_76__10_, r_n_76__9_, r_n_76__8_, r_n_76__7_, r_n_76__6_, r_n_76__5_, r_n_76__4_, r_n_76__3_, r_n_76__2_, r_n_76__1_, r_n_76__0_ } = (N152)? { r_77__63_, r_77__62_, r_77__61_, r_77__60_, r_77__59_, r_77__58_, r_77__57_, r_77__56_, r_77__55_, r_77__54_, r_77__53_, r_77__52_, r_77__51_, r_77__50_, r_77__49_, r_77__48_, r_77__47_, r_77__46_, r_77__45_, r_77__44_, r_77__43_, r_77__42_, r_77__41_, r_77__40_, r_77__39_, r_77__38_, r_77__37_, r_77__36_, r_77__35_, r_77__34_, r_77__33_, r_77__32_, r_77__31_, r_77__30_, r_77__29_, r_77__28_, r_77__27_, r_77__26_, r_77__25_, r_77__24_, r_77__23_, r_77__22_, r_77__21_, r_77__20_, r_77__19_, r_77__18_, r_77__17_, r_77__16_, r_77__15_, r_77__14_, r_77__13_, r_77__12_, r_77__11_, r_77__10_, r_77__9_, r_77__8_, r_77__7_, r_77__6_, r_77__5_, r_77__4_, r_77__3_, r_77__2_, r_77__1_, r_77__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N153)? data_i : 1'b0;
  assign N152 = sel_i[152];
  assign N153 = N1408;
  assign { r_n_77__63_, r_n_77__62_, r_n_77__61_, r_n_77__60_, r_n_77__59_, r_n_77__58_, r_n_77__57_, r_n_77__56_, r_n_77__55_, r_n_77__54_, r_n_77__53_, r_n_77__52_, r_n_77__51_, r_n_77__50_, r_n_77__49_, r_n_77__48_, r_n_77__47_, r_n_77__46_, r_n_77__45_, r_n_77__44_, r_n_77__43_, r_n_77__42_, r_n_77__41_, r_n_77__40_, r_n_77__39_, r_n_77__38_, r_n_77__37_, r_n_77__36_, r_n_77__35_, r_n_77__34_, r_n_77__33_, r_n_77__32_, r_n_77__31_, r_n_77__30_, r_n_77__29_, r_n_77__28_, r_n_77__27_, r_n_77__26_, r_n_77__25_, r_n_77__24_, r_n_77__23_, r_n_77__22_, r_n_77__21_, r_n_77__20_, r_n_77__19_, r_n_77__18_, r_n_77__17_, r_n_77__16_, r_n_77__15_, r_n_77__14_, r_n_77__13_, r_n_77__12_, r_n_77__11_, r_n_77__10_, r_n_77__9_, r_n_77__8_, r_n_77__7_, r_n_77__6_, r_n_77__5_, r_n_77__4_, r_n_77__3_, r_n_77__2_, r_n_77__1_, r_n_77__0_ } = (N154)? { r_78__63_, r_78__62_, r_78__61_, r_78__60_, r_78__59_, r_78__58_, r_78__57_, r_78__56_, r_78__55_, r_78__54_, r_78__53_, r_78__52_, r_78__51_, r_78__50_, r_78__49_, r_78__48_, r_78__47_, r_78__46_, r_78__45_, r_78__44_, r_78__43_, r_78__42_, r_78__41_, r_78__40_, r_78__39_, r_78__38_, r_78__37_, r_78__36_, r_78__35_, r_78__34_, r_78__33_, r_78__32_, r_78__31_, r_78__30_, r_78__29_, r_78__28_, r_78__27_, r_78__26_, r_78__25_, r_78__24_, r_78__23_, r_78__22_, r_78__21_, r_78__20_, r_78__19_, r_78__18_, r_78__17_, r_78__16_, r_78__15_, r_78__14_, r_78__13_, r_78__12_, r_78__11_, r_78__10_, r_78__9_, r_78__8_, r_78__7_, r_78__6_, r_78__5_, r_78__4_, r_78__3_, r_78__2_, r_78__1_, r_78__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N155)? data_i : 1'b0;
  assign N154 = sel_i[154];
  assign N155 = N1413;
  assign { r_n_78__63_, r_n_78__62_, r_n_78__61_, r_n_78__60_, r_n_78__59_, r_n_78__58_, r_n_78__57_, r_n_78__56_, r_n_78__55_, r_n_78__54_, r_n_78__53_, r_n_78__52_, r_n_78__51_, r_n_78__50_, r_n_78__49_, r_n_78__48_, r_n_78__47_, r_n_78__46_, r_n_78__45_, r_n_78__44_, r_n_78__43_, r_n_78__42_, r_n_78__41_, r_n_78__40_, r_n_78__39_, r_n_78__38_, r_n_78__37_, r_n_78__36_, r_n_78__35_, r_n_78__34_, r_n_78__33_, r_n_78__32_, r_n_78__31_, r_n_78__30_, r_n_78__29_, r_n_78__28_, r_n_78__27_, r_n_78__26_, r_n_78__25_, r_n_78__24_, r_n_78__23_, r_n_78__22_, r_n_78__21_, r_n_78__20_, r_n_78__19_, r_n_78__18_, r_n_78__17_, r_n_78__16_, r_n_78__15_, r_n_78__14_, r_n_78__13_, r_n_78__12_, r_n_78__11_, r_n_78__10_, r_n_78__9_, r_n_78__8_, r_n_78__7_, r_n_78__6_, r_n_78__5_, r_n_78__4_, r_n_78__3_, r_n_78__2_, r_n_78__1_, r_n_78__0_ } = (N156)? { r_79__63_, r_79__62_, r_79__61_, r_79__60_, r_79__59_, r_79__58_, r_79__57_, r_79__56_, r_79__55_, r_79__54_, r_79__53_, r_79__52_, r_79__51_, r_79__50_, r_79__49_, r_79__48_, r_79__47_, r_79__46_, r_79__45_, r_79__44_, r_79__43_, r_79__42_, r_79__41_, r_79__40_, r_79__39_, r_79__38_, r_79__37_, r_79__36_, r_79__35_, r_79__34_, r_79__33_, r_79__32_, r_79__31_, r_79__30_, r_79__29_, r_79__28_, r_79__27_, r_79__26_, r_79__25_, r_79__24_, r_79__23_, r_79__22_, r_79__21_, r_79__20_, r_79__19_, r_79__18_, r_79__17_, r_79__16_, r_79__15_, r_79__14_, r_79__13_, r_79__12_, r_79__11_, r_79__10_, r_79__9_, r_79__8_, r_79__7_, r_79__6_, r_79__5_, r_79__4_, r_79__3_, r_79__2_, r_79__1_, r_79__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N157)? data_i : 1'b0;
  assign N156 = sel_i[156];
  assign N157 = N1418;
  assign { r_n_79__63_, r_n_79__62_, r_n_79__61_, r_n_79__60_, r_n_79__59_, r_n_79__58_, r_n_79__57_, r_n_79__56_, r_n_79__55_, r_n_79__54_, r_n_79__53_, r_n_79__52_, r_n_79__51_, r_n_79__50_, r_n_79__49_, r_n_79__48_, r_n_79__47_, r_n_79__46_, r_n_79__45_, r_n_79__44_, r_n_79__43_, r_n_79__42_, r_n_79__41_, r_n_79__40_, r_n_79__39_, r_n_79__38_, r_n_79__37_, r_n_79__36_, r_n_79__35_, r_n_79__34_, r_n_79__33_, r_n_79__32_, r_n_79__31_, r_n_79__30_, r_n_79__29_, r_n_79__28_, r_n_79__27_, r_n_79__26_, r_n_79__25_, r_n_79__24_, r_n_79__23_, r_n_79__22_, r_n_79__21_, r_n_79__20_, r_n_79__19_, r_n_79__18_, r_n_79__17_, r_n_79__16_, r_n_79__15_, r_n_79__14_, r_n_79__13_, r_n_79__12_, r_n_79__11_, r_n_79__10_, r_n_79__9_, r_n_79__8_, r_n_79__7_, r_n_79__6_, r_n_79__5_, r_n_79__4_, r_n_79__3_, r_n_79__2_, r_n_79__1_, r_n_79__0_ } = (N158)? { r_80__63_, r_80__62_, r_80__61_, r_80__60_, r_80__59_, r_80__58_, r_80__57_, r_80__56_, r_80__55_, r_80__54_, r_80__53_, r_80__52_, r_80__51_, r_80__50_, r_80__49_, r_80__48_, r_80__47_, r_80__46_, r_80__45_, r_80__44_, r_80__43_, r_80__42_, r_80__41_, r_80__40_, r_80__39_, r_80__38_, r_80__37_, r_80__36_, r_80__35_, r_80__34_, r_80__33_, r_80__32_, r_80__31_, r_80__30_, r_80__29_, r_80__28_, r_80__27_, r_80__26_, r_80__25_, r_80__24_, r_80__23_, r_80__22_, r_80__21_, r_80__20_, r_80__19_, r_80__18_, r_80__17_, r_80__16_, r_80__15_, r_80__14_, r_80__13_, r_80__12_, r_80__11_, r_80__10_, r_80__9_, r_80__8_, r_80__7_, r_80__6_, r_80__5_, r_80__4_, r_80__3_, r_80__2_, r_80__1_, r_80__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N159)? data_i : 1'b0;
  assign N158 = sel_i[158];
  assign N159 = N1423;
  assign { r_n_80__63_, r_n_80__62_, r_n_80__61_, r_n_80__60_, r_n_80__59_, r_n_80__58_, r_n_80__57_, r_n_80__56_, r_n_80__55_, r_n_80__54_, r_n_80__53_, r_n_80__52_, r_n_80__51_, r_n_80__50_, r_n_80__49_, r_n_80__48_, r_n_80__47_, r_n_80__46_, r_n_80__45_, r_n_80__44_, r_n_80__43_, r_n_80__42_, r_n_80__41_, r_n_80__40_, r_n_80__39_, r_n_80__38_, r_n_80__37_, r_n_80__36_, r_n_80__35_, r_n_80__34_, r_n_80__33_, r_n_80__32_, r_n_80__31_, r_n_80__30_, r_n_80__29_, r_n_80__28_, r_n_80__27_, r_n_80__26_, r_n_80__25_, r_n_80__24_, r_n_80__23_, r_n_80__22_, r_n_80__21_, r_n_80__20_, r_n_80__19_, r_n_80__18_, r_n_80__17_, r_n_80__16_, r_n_80__15_, r_n_80__14_, r_n_80__13_, r_n_80__12_, r_n_80__11_, r_n_80__10_, r_n_80__9_, r_n_80__8_, r_n_80__7_, r_n_80__6_, r_n_80__5_, r_n_80__4_, r_n_80__3_, r_n_80__2_, r_n_80__1_, r_n_80__0_ } = (N160)? { r_81__63_, r_81__62_, r_81__61_, r_81__60_, r_81__59_, r_81__58_, r_81__57_, r_81__56_, r_81__55_, r_81__54_, r_81__53_, r_81__52_, r_81__51_, r_81__50_, r_81__49_, r_81__48_, r_81__47_, r_81__46_, r_81__45_, r_81__44_, r_81__43_, r_81__42_, r_81__41_, r_81__40_, r_81__39_, r_81__38_, r_81__37_, r_81__36_, r_81__35_, r_81__34_, r_81__33_, r_81__32_, r_81__31_, r_81__30_, r_81__29_, r_81__28_, r_81__27_, r_81__26_, r_81__25_, r_81__24_, r_81__23_, r_81__22_, r_81__21_, r_81__20_, r_81__19_, r_81__18_, r_81__17_, r_81__16_, r_81__15_, r_81__14_, r_81__13_, r_81__12_, r_81__11_, r_81__10_, r_81__9_, r_81__8_, r_81__7_, r_81__6_, r_81__5_, r_81__4_, r_81__3_, r_81__2_, r_81__1_, r_81__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N161)? data_i : 1'b0;
  assign N160 = sel_i[160];
  assign N161 = N1428;
  assign { r_n_81__63_, r_n_81__62_, r_n_81__61_, r_n_81__60_, r_n_81__59_, r_n_81__58_, r_n_81__57_, r_n_81__56_, r_n_81__55_, r_n_81__54_, r_n_81__53_, r_n_81__52_, r_n_81__51_, r_n_81__50_, r_n_81__49_, r_n_81__48_, r_n_81__47_, r_n_81__46_, r_n_81__45_, r_n_81__44_, r_n_81__43_, r_n_81__42_, r_n_81__41_, r_n_81__40_, r_n_81__39_, r_n_81__38_, r_n_81__37_, r_n_81__36_, r_n_81__35_, r_n_81__34_, r_n_81__33_, r_n_81__32_, r_n_81__31_, r_n_81__30_, r_n_81__29_, r_n_81__28_, r_n_81__27_, r_n_81__26_, r_n_81__25_, r_n_81__24_, r_n_81__23_, r_n_81__22_, r_n_81__21_, r_n_81__20_, r_n_81__19_, r_n_81__18_, r_n_81__17_, r_n_81__16_, r_n_81__15_, r_n_81__14_, r_n_81__13_, r_n_81__12_, r_n_81__11_, r_n_81__10_, r_n_81__9_, r_n_81__8_, r_n_81__7_, r_n_81__6_, r_n_81__5_, r_n_81__4_, r_n_81__3_, r_n_81__2_, r_n_81__1_, r_n_81__0_ } = (N162)? { r_82__63_, r_82__62_, r_82__61_, r_82__60_, r_82__59_, r_82__58_, r_82__57_, r_82__56_, r_82__55_, r_82__54_, r_82__53_, r_82__52_, r_82__51_, r_82__50_, r_82__49_, r_82__48_, r_82__47_, r_82__46_, r_82__45_, r_82__44_, r_82__43_, r_82__42_, r_82__41_, r_82__40_, r_82__39_, r_82__38_, r_82__37_, r_82__36_, r_82__35_, r_82__34_, r_82__33_, r_82__32_, r_82__31_, r_82__30_, r_82__29_, r_82__28_, r_82__27_, r_82__26_, r_82__25_, r_82__24_, r_82__23_, r_82__22_, r_82__21_, r_82__20_, r_82__19_, r_82__18_, r_82__17_, r_82__16_, r_82__15_, r_82__14_, r_82__13_, r_82__12_, r_82__11_, r_82__10_, r_82__9_, r_82__8_, r_82__7_, r_82__6_, r_82__5_, r_82__4_, r_82__3_, r_82__2_, r_82__1_, r_82__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N163)? data_i : 1'b0;
  assign N162 = sel_i[162];
  assign N163 = N1433;
  assign { r_n_82__63_, r_n_82__62_, r_n_82__61_, r_n_82__60_, r_n_82__59_, r_n_82__58_, r_n_82__57_, r_n_82__56_, r_n_82__55_, r_n_82__54_, r_n_82__53_, r_n_82__52_, r_n_82__51_, r_n_82__50_, r_n_82__49_, r_n_82__48_, r_n_82__47_, r_n_82__46_, r_n_82__45_, r_n_82__44_, r_n_82__43_, r_n_82__42_, r_n_82__41_, r_n_82__40_, r_n_82__39_, r_n_82__38_, r_n_82__37_, r_n_82__36_, r_n_82__35_, r_n_82__34_, r_n_82__33_, r_n_82__32_, r_n_82__31_, r_n_82__30_, r_n_82__29_, r_n_82__28_, r_n_82__27_, r_n_82__26_, r_n_82__25_, r_n_82__24_, r_n_82__23_, r_n_82__22_, r_n_82__21_, r_n_82__20_, r_n_82__19_, r_n_82__18_, r_n_82__17_, r_n_82__16_, r_n_82__15_, r_n_82__14_, r_n_82__13_, r_n_82__12_, r_n_82__11_, r_n_82__10_, r_n_82__9_, r_n_82__8_, r_n_82__7_, r_n_82__6_, r_n_82__5_, r_n_82__4_, r_n_82__3_, r_n_82__2_, r_n_82__1_, r_n_82__0_ } = (N164)? { r_83__63_, r_83__62_, r_83__61_, r_83__60_, r_83__59_, r_83__58_, r_83__57_, r_83__56_, r_83__55_, r_83__54_, r_83__53_, r_83__52_, r_83__51_, r_83__50_, r_83__49_, r_83__48_, r_83__47_, r_83__46_, r_83__45_, r_83__44_, r_83__43_, r_83__42_, r_83__41_, r_83__40_, r_83__39_, r_83__38_, r_83__37_, r_83__36_, r_83__35_, r_83__34_, r_83__33_, r_83__32_, r_83__31_, r_83__30_, r_83__29_, r_83__28_, r_83__27_, r_83__26_, r_83__25_, r_83__24_, r_83__23_, r_83__22_, r_83__21_, r_83__20_, r_83__19_, r_83__18_, r_83__17_, r_83__16_, r_83__15_, r_83__14_, r_83__13_, r_83__12_, r_83__11_, r_83__10_, r_83__9_, r_83__8_, r_83__7_, r_83__6_, r_83__5_, r_83__4_, r_83__3_, r_83__2_, r_83__1_, r_83__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N165)? data_i : 1'b0;
  assign N164 = sel_i[164];
  assign N165 = N1438;
  assign { r_n_83__63_, r_n_83__62_, r_n_83__61_, r_n_83__60_, r_n_83__59_, r_n_83__58_, r_n_83__57_, r_n_83__56_, r_n_83__55_, r_n_83__54_, r_n_83__53_, r_n_83__52_, r_n_83__51_, r_n_83__50_, r_n_83__49_, r_n_83__48_, r_n_83__47_, r_n_83__46_, r_n_83__45_, r_n_83__44_, r_n_83__43_, r_n_83__42_, r_n_83__41_, r_n_83__40_, r_n_83__39_, r_n_83__38_, r_n_83__37_, r_n_83__36_, r_n_83__35_, r_n_83__34_, r_n_83__33_, r_n_83__32_, r_n_83__31_, r_n_83__30_, r_n_83__29_, r_n_83__28_, r_n_83__27_, r_n_83__26_, r_n_83__25_, r_n_83__24_, r_n_83__23_, r_n_83__22_, r_n_83__21_, r_n_83__20_, r_n_83__19_, r_n_83__18_, r_n_83__17_, r_n_83__16_, r_n_83__15_, r_n_83__14_, r_n_83__13_, r_n_83__12_, r_n_83__11_, r_n_83__10_, r_n_83__9_, r_n_83__8_, r_n_83__7_, r_n_83__6_, r_n_83__5_, r_n_83__4_, r_n_83__3_, r_n_83__2_, r_n_83__1_, r_n_83__0_ } = (N166)? { r_84__63_, r_84__62_, r_84__61_, r_84__60_, r_84__59_, r_84__58_, r_84__57_, r_84__56_, r_84__55_, r_84__54_, r_84__53_, r_84__52_, r_84__51_, r_84__50_, r_84__49_, r_84__48_, r_84__47_, r_84__46_, r_84__45_, r_84__44_, r_84__43_, r_84__42_, r_84__41_, r_84__40_, r_84__39_, r_84__38_, r_84__37_, r_84__36_, r_84__35_, r_84__34_, r_84__33_, r_84__32_, r_84__31_, r_84__30_, r_84__29_, r_84__28_, r_84__27_, r_84__26_, r_84__25_, r_84__24_, r_84__23_, r_84__22_, r_84__21_, r_84__20_, r_84__19_, r_84__18_, r_84__17_, r_84__16_, r_84__15_, r_84__14_, r_84__13_, r_84__12_, r_84__11_, r_84__10_, r_84__9_, r_84__8_, r_84__7_, r_84__6_, r_84__5_, r_84__4_, r_84__3_, r_84__2_, r_84__1_, r_84__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N167)? data_i : 1'b0;
  assign N166 = sel_i[166];
  assign N167 = N1443;
  assign { r_n_84__63_, r_n_84__62_, r_n_84__61_, r_n_84__60_, r_n_84__59_, r_n_84__58_, r_n_84__57_, r_n_84__56_, r_n_84__55_, r_n_84__54_, r_n_84__53_, r_n_84__52_, r_n_84__51_, r_n_84__50_, r_n_84__49_, r_n_84__48_, r_n_84__47_, r_n_84__46_, r_n_84__45_, r_n_84__44_, r_n_84__43_, r_n_84__42_, r_n_84__41_, r_n_84__40_, r_n_84__39_, r_n_84__38_, r_n_84__37_, r_n_84__36_, r_n_84__35_, r_n_84__34_, r_n_84__33_, r_n_84__32_, r_n_84__31_, r_n_84__30_, r_n_84__29_, r_n_84__28_, r_n_84__27_, r_n_84__26_, r_n_84__25_, r_n_84__24_, r_n_84__23_, r_n_84__22_, r_n_84__21_, r_n_84__20_, r_n_84__19_, r_n_84__18_, r_n_84__17_, r_n_84__16_, r_n_84__15_, r_n_84__14_, r_n_84__13_, r_n_84__12_, r_n_84__11_, r_n_84__10_, r_n_84__9_, r_n_84__8_, r_n_84__7_, r_n_84__6_, r_n_84__5_, r_n_84__4_, r_n_84__3_, r_n_84__2_, r_n_84__1_, r_n_84__0_ } = (N168)? { r_85__63_, r_85__62_, r_85__61_, r_85__60_, r_85__59_, r_85__58_, r_85__57_, r_85__56_, r_85__55_, r_85__54_, r_85__53_, r_85__52_, r_85__51_, r_85__50_, r_85__49_, r_85__48_, r_85__47_, r_85__46_, r_85__45_, r_85__44_, r_85__43_, r_85__42_, r_85__41_, r_85__40_, r_85__39_, r_85__38_, r_85__37_, r_85__36_, r_85__35_, r_85__34_, r_85__33_, r_85__32_, r_85__31_, r_85__30_, r_85__29_, r_85__28_, r_85__27_, r_85__26_, r_85__25_, r_85__24_, r_85__23_, r_85__22_, r_85__21_, r_85__20_, r_85__19_, r_85__18_, r_85__17_, r_85__16_, r_85__15_, r_85__14_, r_85__13_, r_85__12_, r_85__11_, r_85__10_, r_85__9_, r_85__8_, r_85__7_, r_85__6_, r_85__5_, r_85__4_, r_85__3_, r_85__2_, r_85__1_, r_85__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N169)? data_i : 1'b0;
  assign N168 = sel_i[168];
  assign N169 = N1448;
  assign { r_n_85__63_, r_n_85__62_, r_n_85__61_, r_n_85__60_, r_n_85__59_, r_n_85__58_, r_n_85__57_, r_n_85__56_, r_n_85__55_, r_n_85__54_, r_n_85__53_, r_n_85__52_, r_n_85__51_, r_n_85__50_, r_n_85__49_, r_n_85__48_, r_n_85__47_, r_n_85__46_, r_n_85__45_, r_n_85__44_, r_n_85__43_, r_n_85__42_, r_n_85__41_, r_n_85__40_, r_n_85__39_, r_n_85__38_, r_n_85__37_, r_n_85__36_, r_n_85__35_, r_n_85__34_, r_n_85__33_, r_n_85__32_, r_n_85__31_, r_n_85__30_, r_n_85__29_, r_n_85__28_, r_n_85__27_, r_n_85__26_, r_n_85__25_, r_n_85__24_, r_n_85__23_, r_n_85__22_, r_n_85__21_, r_n_85__20_, r_n_85__19_, r_n_85__18_, r_n_85__17_, r_n_85__16_, r_n_85__15_, r_n_85__14_, r_n_85__13_, r_n_85__12_, r_n_85__11_, r_n_85__10_, r_n_85__9_, r_n_85__8_, r_n_85__7_, r_n_85__6_, r_n_85__5_, r_n_85__4_, r_n_85__3_, r_n_85__2_, r_n_85__1_, r_n_85__0_ } = (N170)? { r_86__63_, r_86__62_, r_86__61_, r_86__60_, r_86__59_, r_86__58_, r_86__57_, r_86__56_, r_86__55_, r_86__54_, r_86__53_, r_86__52_, r_86__51_, r_86__50_, r_86__49_, r_86__48_, r_86__47_, r_86__46_, r_86__45_, r_86__44_, r_86__43_, r_86__42_, r_86__41_, r_86__40_, r_86__39_, r_86__38_, r_86__37_, r_86__36_, r_86__35_, r_86__34_, r_86__33_, r_86__32_, r_86__31_, r_86__30_, r_86__29_, r_86__28_, r_86__27_, r_86__26_, r_86__25_, r_86__24_, r_86__23_, r_86__22_, r_86__21_, r_86__20_, r_86__19_, r_86__18_, r_86__17_, r_86__16_, r_86__15_, r_86__14_, r_86__13_, r_86__12_, r_86__11_, r_86__10_, r_86__9_, r_86__8_, r_86__7_, r_86__6_, r_86__5_, r_86__4_, r_86__3_, r_86__2_, r_86__1_, r_86__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N171)? data_i : 1'b0;
  assign N170 = sel_i[170];
  assign N171 = N1453;
  assign { r_n_86__63_, r_n_86__62_, r_n_86__61_, r_n_86__60_, r_n_86__59_, r_n_86__58_, r_n_86__57_, r_n_86__56_, r_n_86__55_, r_n_86__54_, r_n_86__53_, r_n_86__52_, r_n_86__51_, r_n_86__50_, r_n_86__49_, r_n_86__48_, r_n_86__47_, r_n_86__46_, r_n_86__45_, r_n_86__44_, r_n_86__43_, r_n_86__42_, r_n_86__41_, r_n_86__40_, r_n_86__39_, r_n_86__38_, r_n_86__37_, r_n_86__36_, r_n_86__35_, r_n_86__34_, r_n_86__33_, r_n_86__32_, r_n_86__31_, r_n_86__30_, r_n_86__29_, r_n_86__28_, r_n_86__27_, r_n_86__26_, r_n_86__25_, r_n_86__24_, r_n_86__23_, r_n_86__22_, r_n_86__21_, r_n_86__20_, r_n_86__19_, r_n_86__18_, r_n_86__17_, r_n_86__16_, r_n_86__15_, r_n_86__14_, r_n_86__13_, r_n_86__12_, r_n_86__11_, r_n_86__10_, r_n_86__9_, r_n_86__8_, r_n_86__7_, r_n_86__6_, r_n_86__5_, r_n_86__4_, r_n_86__3_, r_n_86__2_, r_n_86__1_, r_n_86__0_ } = (N172)? { r_87__63_, r_87__62_, r_87__61_, r_87__60_, r_87__59_, r_87__58_, r_87__57_, r_87__56_, r_87__55_, r_87__54_, r_87__53_, r_87__52_, r_87__51_, r_87__50_, r_87__49_, r_87__48_, r_87__47_, r_87__46_, r_87__45_, r_87__44_, r_87__43_, r_87__42_, r_87__41_, r_87__40_, r_87__39_, r_87__38_, r_87__37_, r_87__36_, r_87__35_, r_87__34_, r_87__33_, r_87__32_, r_87__31_, r_87__30_, r_87__29_, r_87__28_, r_87__27_, r_87__26_, r_87__25_, r_87__24_, r_87__23_, r_87__22_, r_87__21_, r_87__20_, r_87__19_, r_87__18_, r_87__17_, r_87__16_, r_87__15_, r_87__14_, r_87__13_, r_87__12_, r_87__11_, r_87__10_, r_87__9_, r_87__8_, r_87__7_, r_87__6_, r_87__5_, r_87__4_, r_87__3_, r_87__2_, r_87__1_, r_87__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N173)? data_i : 1'b0;
  assign N172 = sel_i[172];
  assign N173 = N1458;
  assign { r_n_87__63_, r_n_87__62_, r_n_87__61_, r_n_87__60_, r_n_87__59_, r_n_87__58_, r_n_87__57_, r_n_87__56_, r_n_87__55_, r_n_87__54_, r_n_87__53_, r_n_87__52_, r_n_87__51_, r_n_87__50_, r_n_87__49_, r_n_87__48_, r_n_87__47_, r_n_87__46_, r_n_87__45_, r_n_87__44_, r_n_87__43_, r_n_87__42_, r_n_87__41_, r_n_87__40_, r_n_87__39_, r_n_87__38_, r_n_87__37_, r_n_87__36_, r_n_87__35_, r_n_87__34_, r_n_87__33_, r_n_87__32_, r_n_87__31_, r_n_87__30_, r_n_87__29_, r_n_87__28_, r_n_87__27_, r_n_87__26_, r_n_87__25_, r_n_87__24_, r_n_87__23_, r_n_87__22_, r_n_87__21_, r_n_87__20_, r_n_87__19_, r_n_87__18_, r_n_87__17_, r_n_87__16_, r_n_87__15_, r_n_87__14_, r_n_87__13_, r_n_87__12_, r_n_87__11_, r_n_87__10_, r_n_87__9_, r_n_87__8_, r_n_87__7_, r_n_87__6_, r_n_87__5_, r_n_87__4_, r_n_87__3_, r_n_87__2_, r_n_87__1_, r_n_87__0_ } = (N174)? { r_88__63_, r_88__62_, r_88__61_, r_88__60_, r_88__59_, r_88__58_, r_88__57_, r_88__56_, r_88__55_, r_88__54_, r_88__53_, r_88__52_, r_88__51_, r_88__50_, r_88__49_, r_88__48_, r_88__47_, r_88__46_, r_88__45_, r_88__44_, r_88__43_, r_88__42_, r_88__41_, r_88__40_, r_88__39_, r_88__38_, r_88__37_, r_88__36_, r_88__35_, r_88__34_, r_88__33_, r_88__32_, r_88__31_, r_88__30_, r_88__29_, r_88__28_, r_88__27_, r_88__26_, r_88__25_, r_88__24_, r_88__23_, r_88__22_, r_88__21_, r_88__20_, r_88__19_, r_88__18_, r_88__17_, r_88__16_, r_88__15_, r_88__14_, r_88__13_, r_88__12_, r_88__11_, r_88__10_, r_88__9_, r_88__8_, r_88__7_, r_88__6_, r_88__5_, r_88__4_, r_88__3_, r_88__2_, r_88__1_, r_88__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N175)? data_i : 1'b0;
  assign N174 = sel_i[174];
  assign N175 = N1463;
  assign { r_n_88__63_, r_n_88__62_, r_n_88__61_, r_n_88__60_, r_n_88__59_, r_n_88__58_, r_n_88__57_, r_n_88__56_, r_n_88__55_, r_n_88__54_, r_n_88__53_, r_n_88__52_, r_n_88__51_, r_n_88__50_, r_n_88__49_, r_n_88__48_, r_n_88__47_, r_n_88__46_, r_n_88__45_, r_n_88__44_, r_n_88__43_, r_n_88__42_, r_n_88__41_, r_n_88__40_, r_n_88__39_, r_n_88__38_, r_n_88__37_, r_n_88__36_, r_n_88__35_, r_n_88__34_, r_n_88__33_, r_n_88__32_, r_n_88__31_, r_n_88__30_, r_n_88__29_, r_n_88__28_, r_n_88__27_, r_n_88__26_, r_n_88__25_, r_n_88__24_, r_n_88__23_, r_n_88__22_, r_n_88__21_, r_n_88__20_, r_n_88__19_, r_n_88__18_, r_n_88__17_, r_n_88__16_, r_n_88__15_, r_n_88__14_, r_n_88__13_, r_n_88__12_, r_n_88__11_, r_n_88__10_, r_n_88__9_, r_n_88__8_, r_n_88__7_, r_n_88__6_, r_n_88__5_, r_n_88__4_, r_n_88__3_, r_n_88__2_, r_n_88__1_, r_n_88__0_ } = (N176)? { r_89__63_, r_89__62_, r_89__61_, r_89__60_, r_89__59_, r_89__58_, r_89__57_, r_89__56_, r_89__55_, r_89__54_, r_89__53_, r_89__52_, r_89__51_, r_89__50_, r_89__49_, r_89__48_, r_89__47_, r_89__46_, r_89__45_, r_89__44_, r_89__43_, r_89__42_, r_89__41_, r_89__40_, r_89__39_, r_89__38_, r_89__37_, r_89__36_, r_89__35_, r_89__34_, r_89__33_, r_89__32_, r_89__31_, r_89__30_, r_89__29_, r_89__28_, r_89__27_, r_89__26_, r_89__25_, r_89__24_, r_89__23_, r_89__22_, r_89__21_, r_89__20_, r_89__19_, r_89__18_, r_89__17_, r_89__16_, r_89__15_, r_89__14_, r_89__13_, r_89__12_, r_89__11_, r_89__10_, r_89__9_, r_89__8_, r_89__7_, r_89__6_, r_89__5_, r_89__4_, r_89__3_, r_89__2_, r_89__1_, r_89__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N177)? data_i : 1'b0;
  assign N176 = sel_i[176];
  assign N177 = N1468;
  assign { r_n_89__63_, r_n_89__62_, r_n_89__61_, r_n_89__60_, r_n_89__59_, r_n_89__58_, r_n_89__57_, r_n_89__56_, r_n_89__55_, r_n_89__54_, r_n_89__53_, r_n_89__52_, r_n_89__51_, r_n_89__50_, r_n_89__49_, r_n_89__48_, r_n_89__47_, r_n_89__46_, r_n_89__45_, r_n_89__44_, r_n_89__43_, r_n_89__42_, r_n_89__41_, r_n_89__40_, r_n_89__39_, r_n_89__38_, r_n_89__37_, r_n_89__36_, r_n_89__35_, r_n_89__34_, r_n_89__33_, r_n_89__32_, r_n_89__31_, r_n_89__30_, r_n_89__29_, r_n_89__28_, r_n_89__27_, r_n_89__26_, r_n_89__25_, r_n_89__24_, r_n_89__23_, r_n_89__22_, r_n_89__21_, r_n_89__20_, r_n_89__19_, r_n_89__18_, r_n_89__17_, r_n_89__16_, r_n_89__15_, r_n_89__14_, r_n_89__13_, r_n_89__12_, r_n_89__11_, r_n_89__10_, r_n_89__9_, r_n_89__8_, r_n_89__7_, r_n_89__6_, r_n_89__5_, r_n_89__4_, r_n_89__3_, r_n_89__2_, r_n_89__1_, r_n_89__0_ } = (N178)? { r_90__63_, r_90__62_, r_90__61_, r_90__60_, r_90__59_, r_90__58_, r_90__57_, r_90__56_, r_90__55_, r_90__54_, r_90__53_, r_90__52_, r_90__51_, r_90__50_, r_90__49_, r_90__48_, r_90__47_, r_90__46_, r_90__45_, r_90__44_, r_90__43_, r_90__42_, r_90__41_, r_90__40_, r_90__39_, r_90__38_, r_90__37_, r_90__36_, r_90__35_, r_90__34_, r_90__33_, r_90__32_, r_90__31_, r_90__30_, r_90__29_, r_90__28_, r_90__27_, r_90__26_, r_90__25_, r_90__24_, r_90__23_, r_90__22_, r_90__21_, r_90__20_, r_90__19_, r_90__18_, r_90__17_, r_90__16_, r_90__15_, r_90__14_, r_90__13_, r_90__12_, r_90__11_, r_90__10_, r_90__9_, r_90__8_, r_90__7_, r_90__6_, r_90__5_, r_90__4_, r_90__3_, r_90__2_, r_90__1_, r_90__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N179)? data_i : 1'b0;
  assign N178 = sel_i[178];
  assign N179 = N1473;
  assign { r_n_90__63_, r_n_90__62_, r_n_90__61_, r_n_90__60_, r_n_90__59_, r_n_90__58_, r_n_90__57_, r_n_90__56_, r_n_90__55_, r_n_90__54_, r_n_90__53_, r_n_90__52_, r_n_90__51_, r_n_90__50_, r_n_90__49_, r_n_90__48_, r_n_90__47_, r_n_90__46_, r_n_90__45_, r_n_90__44_, r_n_90__43_, r_n_90__42_, r_n_90__41_, r_n_90__40_, r_n_90__39_, r_n_90__38_, r_n_90__37_, r_n_90__36_, r_n_90__35_, r_n_90__34_, r_n_90__33_, r_n_90__32_, r_n_90__31_, r_n_90__30_, r_n_90__29_, r_n_90__28_, r_n_90__27_, r_n_90__26_, r_n_90__25_, r_n_90__24_, r_n_90__23_, r_n_90__22_, r_n_90__21_, r_n_90__20_, r_n_90__19_, r_n_90__18_, r_n_90__17_, r_n_90__16_, r_n_90__15_, r_n_90__14_, r_n_90__13_, r_n_90__12_, r_n_90__11_, r_n_90__10_, r_n_90__9_, r_n_90__8_, r_n_90__7_, r_n_90__6_, r_n_90__5_, r_n_90__4_, r_n_90__3_, r_n_90__2_, r_n_90__1_, r_n_90__0_ } = (N180)? { r_91__63_, r_91__62_, r_91__61_, r_91__60_, r_91__59_, r_91__58_, r_91__57_, r_91__56_, r_91__55_, r_91__54_, r_91__53_, r_91__52_, r_91__51_, r_91__50_, r_91__49_, r_91__48_, r_91__47_, r_91__46_, r_91__45_, r_91__44_, r_91__43_, r_91__42_, r_91__41_, r_91__40_, r_91__39_, r_91__38_, r_91__37_, r_91__36_, r_91__35_, r_91__34_, r_91__33_, r_91__32_, r_91__31_, r_91__30_, r_91__29_, r_91__28_, r_91__27_, r_91__26_, r_91__25_, r_91__24_, r_91__23_, r_91__22_, r_91__21_, r_91__20_, r_91__19_, r_91__18_, r_91__17_, r_91__16_, r_91__15_, r_91__14_, r_91__13_, r_91__12_, r_91__11_, r_91__10_, r_91__9_, r_91__8_, r_91__7_, r_91__6_, r_91__5_, r_91__4_, r_91__3_, r_91__2_, r_91__1_, r_91__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N181)? data_i : 1'b0;
  assign N180 = sel_i[180];
  assign N181 = N1478;
  assign { r_n_91__63_, r_n_91__62_, r_n_91__61_, r_n_91__60_, r_n_91__59_, r_n_91__58_, r_n_91__57_, r_n_91__56_, r_n_91__55_, r_n_91__54_, r_n_91__53_, r_n_91__52_, r_n_91__51_, r_n_91__50_, r_n_91__49_, r_n_91__48_, r_n_91__47_, r_n_91__46_, r_n_91__45_, r_n_91__44_, r_n_91__43_, r_n_91__42_, r_n_91__41_, r_n_91__40_, r_n_91__39_, r_n_91__38_, r_n_91__37_, r_n_91__36_, r_n_91__35_, r_n_91__34_, r_n_91__33_, r_n_91__32_, r_n_91__31_, r_n_91__30_, r_n_91__29_, r_n_91__28_, r_n_91__27_, r_n_91__26_, r_n_91__25_, r_n_91__24_, r_n_91__23_, r_n_91__22_, r_n_91__21_, r_n_91__20_, r_n_91__19_, r_n_91__18_, r_n_91__17_, r_n_91__16_, r_n_91__15_, r_n_91__14_, r_n_91__13_, r_n_91__12_, r_n_91__11_, r_n_91__10_, r_n_91__9_, r_n_91__8_, r_n_91__7_, r_n_91__6_, r_n_91__5_, r_n_91__4_, r_n_91__3_, r_n_91__2_, r_n_91__1_, r_n_91__0_ } = (N182)? { r_92__63_, r_92__62_, r_92__61_, r_92__60_, r_92__59_, r_92__58_, r_92__57_, r_92__56_, r_92__55_, r_92__54_, r_92__53_, r_92__52_, r_92__51_, r_92__50_, r_92__49_, r_92__48_, r_92__47_, r_92__46_, r_92__45_, r_92__44_, r_92__43_, r_92__42_, r_92__41_, r_92__40_, r_92__39_, r_92__38_, r_92__37_, r_92__36_, r_92__35_, r_92__34_, r_92__33_, r_92__32_, r_92__31_, r_92__30_, r_92__29_, r_92__28_, r_92__27_, r_92__26_, r_92__25_, r_92__24_, r_92__23_, r_92__22_, r_92__21_, r_92__20_, r_92__19_, r_92__18_, r_92__17_, r_92__16_, r_92__15_, r_92__14_, r_92__13_, r_92__12_, r_92__11_, r_92__10_, r_92__9_, r_92__8_, r_92__7_, r_92__6_, r_92__5_, r_92__4_, r_92__3_, r_92__2_, r_92__1_, r_92__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N183)? data_i : 1'b0;
  assign N182 = sel_i[182];
  assign N183 = N1483;
  assign { r_n_92__63_, r_n_92__62_, r_n_92__61_, r_n_92__60_, r_n_92__59_, r_n_92__58_, r_n_92__57_, r_n_92__56_, r_n_92__55_, r_n_92__54_, r_n_92__53_, r_n_92__52_, r_n_92__51_, r_n_92__50_, r_n_92__49_, r_n_92__48_, r_n_92__47_, r_n_92__46_, r_n_92__45_, r_n_92__44_, r_n_92__43_, r_n_92__42_, r_n_92__41_, r_n_92__40_, r_n_92__39_, r_n_92__38_, r_n_92__37_, r_n_92__36_, r_n_92__35_, r_n_92__34_, r_n_92__33_, r_n_92__32_, r_n_92__31_, r_n_92__30_, r_n_92__29_, r_n_92__28_, r_n_92__27_, r_n_92__26_, r_n_92__25_, r_n_92__24_, r_n_92__23_, r_n_92__22_, r_n_92__21_, r_n_92__20_, r_n_92__19_, r_n_92__18_, r_n_92__17_, r_n_92__16_, r_n_92__15_, r_n_92__14_, r_n_92__13_, r_n_92__12_, r_n_92__11_, r_n_92__10_, r_n_92__9_, r_n_92__8_, r_n_92__7_, r_n_92__6_, r_n_92__5_, r_n_92__4_, r_n_92__3_, r_n_92__2_, r_n_92__1_, r_n_92__0_ } = (N184)? { r_93__63_, r_93__62_, r_93__61_, r_93__60_, r_93__59_, r_93__58_, r_93__57_, r_93__56_, r_93__55_, r_93__54_, r_93__53_, r_93__52_, r_93__51_, r_93__50_, r_93__49_, r_93__48_, r_93__47_, r_93__46_, r_93__45_, r_93__44_, r_93__43_, r_93__42_, r_93__41_, r_93__40_, r_93__39_, r_93__38_, r_93__37_, r_93__36_, r_93__35_, r_93__34_, r_93__33_, r_93__32_, r_93__31_, r_93__30_, r_93__29_, r_93__28_, r_93__27_, r_93__26_, r_93__25_, r_93__24_, r_93__23_, r_93__22_, r_93__21_, r_93__20_, r_93__19_, r_93__18_, r_93__17_, r_93__16_, r_93__15_, r_93__14_, r_93__13_, r_93__12_, r_93__11_, r_93__10_, r_93__9_, r_93__8_, r_93__7_, r_93__6_, r_93__5_, r_93__4_, r_93__3_, r_93__2_, r_93__1_, r_93__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N185)? data_i : 1'b0;
  assign N184 = sel_i[184];
  assign N185 = N1488;
  assign { r_n_93__63_, r_n_93__62_, r_n_93__61_, r_n_93__60_, r_n_93__59_, r_n_93__58_, r_n_93__57_, r_n_93__56_, r_n_93__55_, r_n_93__54_, r_n_93__53_, r_n_93__52_, r_n_93__51_, r_n_93__50_, r_n_93__49_, r_n_93__48_, r_n_93__47_, r_n_93__46_, r_n_93__45_, r_n_93__44_, r_n_93__43_, r_n_93__42_, r_n_93__41_, r_n_93__40_, r_n_93__39_, r_n_93__38_, r_n_93__37_, r_n_93__36_, r_n_93__35_, r_n_93__34_, r_n_93__33_, r_n_93__32_, r_n_93__31_, r_n_93__30_, r_n_93__29_, r_n_93__28_, r_n_93__27_, r_n_93__26_, r_n_93__25_, r_n_93__24_, r_n_93__23_, r_n_93__22_, r_n_93__21_, r_n_93__20_, r_n_93__19_, r_n_93__18_, r_n_93__17_, r_n_93__16_, r_n_93__15_, r_n_93__14_, r_n_93__13_, r_n_93__12_, r_n_93__11_, r_n_93__10_, r_n_93__9_, r_n_93__8_, r_n_93__7_, r_n_93__6_, r_n_93__5_, r_n_93__4_, r_n_93__3_, r_n_93__2_, r_n_93__1_, r_n_93__0_ } = (N186)? { r_94__63_, r_94__62_, r_94__61_, r_94__60_, r_94__59_, r_94__58_, r_94__57_, r_94__56_, r_94__55_, r_94__54_, r_94__53_, r_94__52_, r_94__51_, r_94__50_, r_94__49_, r_94__48_, r_94__47_, r_94__46_, r_94__45_, r_94__44_, r_94__43_, r_94__42_, r_94__41_, r_94__40_, r_94__39_, r_94__38_, r_94__37_, r_94__36_, r_94__35_, r_94__34_, r_94__33_, r_94__32_, r_94__31_, r_94__30_, r_94__29_, r_94__28_, r_94__27_, r_94__26_, r_94__25_, r_94__24_, r_94__23_, r_94__22_, r_94__21_, r_94__20_, r_94__19_, r_94__18_, r_94__17_, r_94__16_, r_94__15_, r_94__14_, r_94__13_, r_94__12_, r_94__11_, r_94__10_, r_94__9_, r_94__8_, r_94__7_, r_94__6_, r_94__5_, r_94__4_, r_94__3_, r_94__2_, r_94__1_, r_94__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N187)? data_i : 1'b0;
  assign N186 = sel_i[186];
  assign N187 = N1493;
  assign { r_n_94__63_, r_n_94__62_, r_n_94__61_, r_n_94__60_, r_n_94__59_, r_n_94__58_, r_n_94__57_, r_n_94__56_, r_n_94__55_, r_n_94__54_, r_n_94__53_, r_n_94__52_, r_n_94__51_, r_n_94__50_, r_n_94__49_, r_n_94__48_, r_n_94__47_, r_n_94__46_, r_n_94__45_, r_n_94__44_, r_n_94__43_, r_n_94__42_, r_n_94__41_, r_n_94__40_, r_n_94__39_, r_n_94__38_, r_n_94__37_, r_n_94__36_, r_n_94__35_, r_n_94__34_, r_n_94__33_, r_n_94__32_, r_n_94__31_, r_n_94__30_, r_n_94__29_, r_n_94__28_, r_n_94__27_, r_n_94__26_, r_n_94__25_, r_n_94__24_, r_n_94__23_, r_n_94__22_, r_n_94__21_, r_n_94__20_, r_n_94__19_, r_n_94__18_, r_n_94__17_, r_n_94__16_, r_n_94__15_, r_n_94__14_, r_n_94__13_, r_n_94__12_, r_n_94__11_, r_n_94__10_, r_n_94__9_, r_n_94__8_, r_n_94__7_, r_n_94__6_, r_n_94__5_, r_n_94__4_, r_n_94__3_, r_n_94__2_, r_n_94__1_, r_n_94__0_ } = (N188)? { r_95__63_, r_95__62_, r_95__61_, r_95__60_, r_95__59_, r_95__58_, r_95__57_, r_95__56_, r_95__55_, r_95__54_, r_95__53_, r_95__52_, r_95__51_, r_95__50_, r_95__49_, r_95__48_, r_95__47_, r_95__46_, r_95__45_, r_95__44_, r_95__43_, r_95__42_, r_95__41_, r_95__40_, r_95__39_, r_95__38_, r_95__37_, r_95__36_, r_95__35_, r_95__34_, r_95__33_, r_95__32_, r_95__31_, r_95__30_, r_95__29_, r_95__28_, r_95__27_, r_95__26_, r_95__25_, r_95__24_, r_95__23_, r_95__22_, r_95__21_, r_95__20_, r_95__19_, r_95__18_, r_95__17_, r_95__16_, r_95__15_, r_95__14_, r_95__13_, r_95__12_, r_95__11_, r_95__10_, r_95__9_, r_95__8_, r_95__7_, r_95__6_, r_95__5_, r_95__4_, r_95__3_, r_95__2_, r_95__1_, r_95__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N189)? data_i : 1'b0;
  assign N188 = sel_i[188];
  assign N189 = N1498;
  assign { r_n_95__63_, r_n_95__62_, r_n_95__61_, r_n_95__60_, r_n_95__59_, r_n_95__58_, r_n_95__57_, r_n_95__56_, r_n_95__55_, r_n_95__54_, r_n_95__53_, r_n_95__52_, r_n_95__51_, r_n_95__50_, r_n_95__49_, r_n_95__48_, r_n_95__47_, r_n_95__46_, r_n_95__45_, r_n_95__44_, r_n_95__43_, r_n_95__42_, r_n_95__41_, r_n_95__40_, r_n_95__39_, r_n_95__38_, r_n_95__37_, r_n_95__36_, r_n_95__35_, r_n_95__34_, r_n_95__33_, r_n_95__32_, r_n_95__31_, r_n_95__30_, r_n_95__29_, r_n_95__28_, r_n_95__27_, r_n_95__26_, r_n_95__25_, r_n_95__24_, r_n_95__23_, r_n_95__22_, r_n_95__21_, r_n_95__20_, r_n_95__19_, r_n_95__18_, r_n_95__17_, r_n_95__16_, r_n_95__15_, r_n_95__14_, r_n_95__13_, r_n_95__12_, r_n_95__11_, r_n_95__10_, r_n_95__9_, r_n_95__8_, r_n_95__7_, r_n_95__6_, r_n_95__5_, r_n_95__4_, r_n_95__3_, r_n_95__2_, r_n_95__1_, r_n_95__0_ } = (N190)? { r_96__63_, r_96__62_, r_96__61_, r_96__60_, r_96__59_, r_96__58_, r_96__57_, r_96__56_, r_96__55_, r_96__54_, r_96__53_, r_96__52_, r_96__51_, r_96__50_, r_96__49_, r_96__48_, r_96__47_, r_96__46_, r_96__45_, r_96__44_, r_96__43_, r_96__42_, r_96__41_, r_96__40_, r_96__39_, r_96__38_, r_96__37_, r_96__36_, r_96__35_, r_96__34_, r_96__33_, r_96__32_, r_96__31_, r_96__30_, r_96__29_, r_96__28_, r_96__27_, r_96__26_, r_96__25_, r_96__24_, r_96__23_, r_96__22_, r_96__21_, r_96__20_, r_96__19_, r_96__18_, r_96__17_, r_96__16_, r_96__15_, r_96__14_, r_96__13_, r_96__12_, r_96__11_, r_96__10_, r_96__9_, r_96__8_, r_96__7_, r_96__6_, r_96__5_, r_96__4_, r_96__3_, r_96__2_, r_96__1_, r_96__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N191)? data_i : 1'b0;
  assign N190 = sel_i[190];
  assign N191 = N1503;
  assign { r_n_96__63_, r_n_96__62_, r_n_96__61_, r_n_96__60_, r_n_96__59_, r_n_96__58_, r_n_96__57_, r_n_96__56_, r_n_96__55_, r_n_96__54_, r_n_96__53_, r_n_96__52_, r_n_96__51_, r_n_96__50_, r_n_96__49_, r_n_96__48_, r_n_96__47_, r_n_96__46_, r_n_96__45_, r_n_96__44_, r_n_96__43_, r_n_96__42_, r_n_96__41_, r_n_96__40_, r_n_96__39_, r_n_96__38_, r_n_96__37_, r_n_96__36_, r_n_96__35_, r_n_96__34_, r_n_96__33_, r_n_96__32_, r_n_96__31_, r_n_96__30_, r_n_96__29_, r_n_96__28_, r_n_96__27_, r_n_96__26_, r_n_96__25_, r_n_96__24_, r_n_96__23_, r_n_96__22_, r_n_96__21_, r_n_96__20_, r_n_96__19_, r_n_96__18_, r_n_96__17_, r_n_96__16_, r_n_96__15_, r_n_96__14_, r_n_96__13_, r_n_96__12_, r_n_96__11_, r_n_96__10_, r_n_96__9_, r_n_96__8_, r_n_96__7_, r_n_96__6_, r_n_96__5_, r_n_96__4_, r_n_96__3_, r_n_96__2_, r_n_96__1_, r_n_96__0_ } = (N192)? { r_97__63_, r_97__62_, r_97__61_, r_97__60_, r_97__59_, r_97__58_, r_97__57_, r_97__56_, r_97__55_, r_97__54_, r_97__53_, r_97__52_, r_97__51_, r_97__50_, r_97__49_, r_97__48_, r_97__47_, r_97__46_, r_97__45_, r_97__44_, r_97__43_, r_97__42_, r_97__41_, r_97__40_, r_97__39_, r_97__38_, r_97__37_, r_97__36_, r_97__35_, r_97__34_, r_97__33_, r_97__32_, r_97__31_, r_97__30_, r_97__29_, r_97__28_, r_97__27_, r_97__26_, r_97__25_, r_97__24_, r_97__23_, r_97__22_, r_97__21_, r_97__20_, r_97__19_, r_97__18_, r_97__17_, r_97__16_, r_97__15_, r_97__14_, r_97__13_, r_97__12_, r_97__11_, r_97__10_, r_97__9_, r_97__8_, r_97__7_, r_97__6_, r_97__5_, r_97__4_, r_97__3_, r_97__2_, r_97__1_, r_97__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N193)? data_i : 1'b0;
  assign N192 = sel_i[192];
  assign N193 = N1508;
  assign { r_n_97__63_, r_n_97__62_, r_n_97__61_, r_n_97__60_, r_n_97__59_, r_n_97__58_, r_n_97__57_, r_n_97__56_, r_n_97__55_, r_n_97__54_, r_n_97__53_, r_n_97__52_, r_n_97__51_, r_n_97__50_, r_n_97__49_, r_n_97__48_, r_n_97__47_, r_n_97__46_, r_n_97__45_, r_n_97__44_, r_n_97__43_, r_n_97__42_, r_n_97__41_, r_n_97__40_, r_n_97__39_, r_n_97__38_, r_n_97__37_, r_n_97__36_, r_n_97__35_, r_n_97__34_, r_n_97__33_, r_n_97__32_, r_n_97__31_, r_n_97__30_, r_n_97__29_, r_n_97__28_, r_n_97__27_, r_n_97__26_, r_n_97__25_, r_n_97__24_, r_n_97__23_, r_n_97__22_, r_n_97__21_, r_n_97__20_, r_n_97__19_, r_n_97__18_, r_n_97__17_, r_n_97__16_, r_n_97__15_, r_n_97__14_, r_n_97__13_, r_n_97__12_, r_n_97__11_, r_n_97__10_, r_n_97__9_, r_n_97__8_, r_n_97__7_, r_n_97__6_, r_n_97__5_, r_n_97__4_, r_n_97__3_, r_n_97__2_, r_n_97__1_, r_n_97__0_ } = (N194)? { r_98__63_, r_98__62_, r_98__61_, r_98__60_, r_98__59_, r_98__58_, r_98__57_, r_98__56_, r_98__55_, r_98__54_, r_98__53_, r_98__52_, r_98__51_, r_98__50_, r_98__49_, r_98__48_, r_98__47_, r_98__46_, r_98__45_, r_98__44_, r_98__43_, r_98__42_, r_98__41_, r_98__40_, r_98__39_, r_98__38_, r_98__37_, r_98__36_, r_98__35_, r_98__34_, r_98__33_, r_98__32_, r_98__31_, r_98__30_, r_98__29_, r_98__28_, r_98__27_, r_98__26_, r_98__25_, r_98__24_, r_98__23_, r_98__22_, r_98__21_, r_98__20_, r_98__19_, r_98__18_, r_98__17_, r_98__16_, r_98__15_, r_98__14_, r_98__13_, r_98__12_, r_98__11_, r_98__10_, r_98__9_, r_98__8_, r_98__7_, r_98__6_, r_98__5_, r_98__4_, r_98__3_, r_98__2_, r_98__1_, r_98__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N195)? data_i : 1'b0;
  assign N194 = sel_i[194];
  assign N195 = N1513;
  assign { r_n_98__63_, r_n_98__62_, r_n_98__61_, r_n_98__60_, r_n_98__59_, r_n_98__58_, r_n_98__57_, r_n_98__56_, r_n_98__55_, r_n_98__54_, r_n_98__53_, r_n_98__52_, r_n_98__51_, r_n_98__50_, r_n_98__49_, r_n_98__48_, r_n_98__47_, r_n_98__46_, r_n_98__45_, r_n_98__44_, r_n_98__43_, r_n_98__42_, r_n_98__41_, r_n_98__40_, r_n_98__39_, r_n_98__38_, r_n_98__37_, r_n_98__36_, r_n_98__35_, r_n_98__34_, r_n_98__33_, r_n_98__32_, r_n_98__31_, r_n_98__30_, r_n_98__29_, r_n_98__28_, r_n_98__27_, r_n_98__26_, r_n_98__25_, r_n_98__24_, r_n_98__23_, r_n_98__22_, r_n_98__21_, r_n_98__20_, r_n_98__19_, r_n_98__18_, r_n_98__17_, r_n_98__16_, r_n_98__15_, r_n_98__14_, r_n_98__13_, r_n_98__12_, r_n_98__11_, r_n_98__10_, r_n_98__9_, r_n_98__8_, r_n_98__7_, r_n_98__6_, r_n_98__5_, r_n_98__4_, r_n_98__3_, r_n_98__2_, r_n_98__1_, r_n_98__0_ } = (N196)? { r_99__63_, r_99__62_, r_99__61_, r_99__60_, r_99__59_, r_99__58_, r_99__57_, r_99__56_, r_99__55_, r_99__54_, r_99__53_, r_99__52_, r_99__51_, r_99__50_, r_99__49_, r_99__48_, r_99__47_, r_99__46_, r_99__45_, r_99__44_, r_99__43_, r_99__42_, r_99__41_, r_99__40_, r_99__39_, r_99__38_, r_99__37_, r_99__36_, r_99__35_, r_99__34_, r_99__33_, r_99__32_, r_99__31_, r_99__30_, r_99__29_, r_99__28_, r_99__27_, r_99__26_, r_99__25_, r_99__24_, r_99__23_, r_99__22_, r_99__21_, r_99__20_, r_99__19_, r_99__18_, r_99__17_, r_99__16_, r_99__15_, r_99__14_, r_99__13_, r_99__12_, r_99__11_, r_99__10_, r_99__9_, r_99__8_, r_99__7_, r_99__6_, r_99__5_, r_99__4_, r_99__3_, r_99__2_, r_99__1_, r_99__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N197)? data_i : 1'b0;
  assign N196 = sel_i[196];
  assign N197 = N1518;
  assign { r_n_99__63_, r_n_99__62_, r_n_99__61_, r_n_99__60_, r_n_99__59_, r_n_99__58_, r_n_99__57_, r_n_99__56_, r_n_99__55_, r_n_99__54_, r_n_99__53_, r_n_99__52_, r_n_99__51_, r_n_99__50_, r_n_99__49_, r_n_99__48_, r_n_99__47_, r_n_99__46_, r_n_99__45_, r_n_99__44_, r_n_99__43_, r_n_99__42_, r_n_99__41_, r_n_99__40_, r_n_99__39_, r_n_99__38_, r_n_99__37_, r_n_99__36_, r_n_99__35_, r_n_99__34_, r_n_99__33_, r_n_99__32_, r_n_99__31_, r_n_99__30_, r_n_99__29_, r_n_99__28_, r_n_99__27_, r_n_99__26_, r_n_99__25_, r_n_99__24_, r_n_99__23_, r_n_99__22_, r_n_99__21_, r_n_99__20_, r_n_99__19_, r_n_99__18_, r_n_99__17_, r_n_99__16_, r_n_99__15_, r_n_99__14_, r_n_99__13_, r_n_99__12_, r_n_99__11_, r_n_99__10_, r_n_99__9_, r_n_99__8_, r_n_99__7_, r_n_99__6_, r_n_99__5_, r_n_99__4_, r_n_99__3_, r_n_99__2_, r_n_99__1_, r_n_99__0_ } = (N198)? { r_100__63_, r_100__62_, r_100__61_, r_100__60_, r_100__59_, r_100__58_, r_100__57_, r_100__56_, r_100__55_, r_100__54_, r_100__53_, r_100__52_, r_100__51_, r_100__50_, r_100__49_, r_100__48_, r_100__47_, r_100__46_, r_100__45_, r_100__44_, r_100__43_, r_100__42_, r_100__41_, r_100__40_, r_100__39_, r_100__38_, r_100__37_, r_100__36_, r_100__35_, r_100__34_, r_100__33_, r_100__32_, r_100__31_, r_100__30_, r_100__29_, r_100__28_, r_100__27_, r_100__26_, r_100__25_, r_100__24_, r_100__23_, r_100__22_, r_100__21_, r_100__20_, r_100__19_, r_100__18_, r_100__17_, r_100__16_, r_100__15_, r_100__14_, r_100__13_, r_100__12_, r_100__11_, r_100__10_, r_100__9_, r_100__8_, r_100__7_, r_100__6_, r_100__5_, r_100__4_, r_100__3_, r_100__2_, r_100__1_, r_100__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N199)? data_i : 1'b0;
  assign N198 = sel_i[198];
  assign N199 = N1523;
  assign { r_n_100__63_, r_n_100__62_, r_n_100__61_, r_n_100__60_, r_n_100__59_, r_n_100__58_, r_n_100__57_, r_n_100__56_, r_n_100__55_, r_n_100__54_, r_n_100__53_, r_n_100__52_, r_n_100__51_, r_n_100__50_, r_n_100__49_, r_n_100__48_, r_n_100__47_, r_n_100__46_, r_n_100__45_, r_n_100__44_, r_n_100__43_, r_n_100__42_, r_n_100__41_, r_n_100__40_, r_n_100__39_, r_n_100__38_, r_n_100__37_, r_n_100__36_, r_n_100__35_, r_n_100__34_, r_n_100__33_, r_n_100__32_, r_n_100__31_, r_n_100__30_, r_n_100__29_, r_n_100__28_, r_n_100__27_, r_n_100__26_, r_n_100__25_, r_n_100__24_, r_n_100__23_, r_n_100__22_, r_n_100__21_, r_n_100__20_, r_n_100__19_, r_n_100__18_, r_n_100__17_, r_n_100__16_, r_n_100__15_, r_n_100__14_, r_n_100__13_, r_n_100__12_, r_n_100__11_, r_n_100__10_, r_n_100__9_, r_n_100__8_, r_n_100__7_, r_n_100__6_, r_n_100__5_, r_n_100__4_, r_n_100__3_, r_n_100__2_, r_n_100__1_, r_n_100__0_ } = (N200)? { r_101__63_, r_101__62_, r_101__61_, r_101__60_, r_101__59_, r_101__58_, r_101__57_, r_101__56_, r_101__55_, r_101__54_, r_101__53_, r_101__52_, r_101__51_, r_101__50_, r_101__49_, r_101__48_, r_101__47_, r_101__46_, r_101__45_, r_101__44_, r_101__43_, r_101__42_, r_101__41_, r_101__40_, r_101__39_, r_101__38_, r_101__37_, r_101__36_, r_101__35_, r_101__34_, r_101__33_, r_101__32_, r_101__31_, r_101__30_, r_101__29_, r_101__28_, r_101__27_, r_101__26_, r_101__25_, r_101__24_, r_101__23_, r_101__22_, r_101__21_, r_101__20_, r_101__19_, r_101__18_, r_101__17_, r_101__16_, r_101__15_, r_101__14_, r_101__13_, r_101__12_, r_101__11_, r_101__10_, r_101__9_, r_101__8_, r_101__7_, r_101__6_, r_101__5_, r_101__4_, r_101__3_, r_101__2_, r_101__1_, r_101__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N201)? data_i : 1'b0;
  assign N200 = sel_i[200];
  assign N201 = N1528;
  assign { r_n_101__63_, r_n_101__62_, r_n_101__61_, r_n_101__60_, r_n_101__59_, r_n_101__58_, r_n_101__57_, r_n_101__56_, r_n_101__55_, r_n_101__54_, r_n_101__53_, r_n_101__52_, r_n_101__51_, r_n_101__50_, r_n_101__49_, r_n_101__48_, r_n_101__47_, r_n_101__46_, r_n_101__45_, r_n_101__44_, r_n_101__43_, r_n_101__42_, r_n_101__41_, r_n_101__40_, r_n_101__39_, r_n_101__38_, r_n_101__37_, r_n_101__36_, r_n_101__35_, r_n_101__34_, r_n_101__33_, r_n_101__32_, r_n_101__31_, r_n_101__30_, r_n_101__29_, r_n_101__28_, r_n_101__27_, r_n_101__26_, r_n_101__25_, r_n_101__24_, r_n_101__23_, r_n_101__22_, r_n_101__21_, r_n_101__20_, r_n_101__19_, r_n_101__18_, r_n_101__17_, r_n_101__16_, r_n_101__15_, r_n_101__14_, r_n_101__13_, r_n_101__12_, r_n_101__11_, r_n_101__10_, r_n_101__9_, r_n_101__8_, r_n_101__7_, r_n_101__6_, r_n_101__5_, r_n_101__4_, r_n_101__3_, r_n_101__2_, r_n_101__1_, r_n_101__0_ } = (N202)? { r_102__63_, r_102__62_, r_102__61_, r_102__60_, r_102__59_, r_102__58_, r_102__57_, r_102__56_, r_102__55_, r_102__54_, r_102__53_, r_102__52_, r_102__51_, r_102__50_, r_102__49_, r_102__48_, r_102__47_, r_102__46_, r_102__45_, r_102__44_, r_102__43_, r_102__42_, r_102__41_, r_102__40_, r_102__39_, r_102__38_, r_102__37_, r_102__36_, r_102__35_, r_102__34_, r_102__33_, r_102__32_, r_102__31_, r_102__30_, r_102__29_, r_102__28_, r_102__27_, r_102__26_, r_102__25_, r_102__24_, r_102__23_, r_102__22_, r_102__21_, r_102__20_, r_102__19_, r_102__18_, r_102__17_, r_102__16_, r_102__15_, r_102__14_, r_102__13_, r_102__12_, r_102__11_, r_102__10_, r_102__9_, r_102__8_, r_102__7_, r_102__6_, r_102__5_, r_102__4_, r_102__3_, r_102__2_, r_102__1_, r_102__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N203)? data_i : 1'b0;
  assign N202 = sel_i[202];
  assign N203 = N1533;
  assign { r_n_102__63_, r_n_102__62_, r_n_102__61_, r_n_102__60_, r_n_102__59_, r_n_102__58_, r_n_102__57_, r_n_102__56_, r_n_102__55_, r_n_102__54_, r_n_102__53_, r_n_102__52_, r_n_102__51_, r_n_102__50_, r_n_102__49_, r_n_102__48_, r_n_102__47_, r_n_102__46_, r_n_102__45_, r_n_102__44_, r_n_102__43_, r_n_102__42_, r_n_102__41_, r_n_102__40_, r_n_102__39_, r_n_102__38_, r_n_102__37_, r_n_102__36_, r_n_102__35_, r_n_102__34_, r_n_102__33_, r_n_102__32_, r_n_102__31_, r_n_102__30_, r_n_102__29_, r_n_102__28_, r_n_102__27_, r_n_102__26_, r_n_102__25_, r_n_102__24_, r_n_102__23_, r_n_102__22_, r_n_102__21_, r_n_102__20_, r_n_102__19_, r_n_102__18_, r_n_102__17_, r_n_102__16_, r_n_102__15_, r_n_102__14_, r_n_102__13_, r_n_102__12_, r_n_102__11_, r_n_102__10_, r_n_102__9_, r_n_102__8_, r_n_102__7_, r_n_102__6_, r_n_102__5_, r_n_102__4_, r_n_102__3_, r_n_102__2_, r_n_102__1_, r_n_102__0_ } = (N204)? { r_103__63_, r_103__62_, r_103__61_, r_103__60_, r_103__59_, r_103__58_, r_103__57_, r_103__56_, r_103__55_, r_103__54_, r_103__53_, r_103__52_, r_103__51_, r_103__50_, r_103__49_, r_103__48_, r_103__47_, r_103__46_, r_103__45_, r_103__44_, r_103__43_, r_103__42_, r_103__41_, r_103__40_, r_103__39_, r_103__38_, r_103__37_, r_103__36_, r_103__35_, r_103__34_, r_103__33_, r_103__32_, r_103__31_, r_103__30_, r_103__29_, r_103__28_, r_103__27_, r_103__26_, r_103__25_, r_103__24_, r_103__23_, r_103__22_, r_103__21_, r_103__20_, r_103__19_, r_103__18_, r_103__17_, r_103__16_, r_103__15_, r_103__14_, r_103__13_, r_103__12_, r_103__11_, r_103__10_, r_103__9_, r_103__8_, r_103__7_, r_103__6_, r_103__5_, r_103__4_, r_103__3_, r_103__2_, r_103__1_, r_103__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N205)? data_i : 1'b0;
  assign N204 = sel_i[204];
  assign N205 = N1538;
  assign { r_n_103__63_, r_n_103__62_, r_n_103__61_, r_n_103__60_, r_n_103__59_, r_n_103__58_, r_n_103__57_, r_n_103__56_, r_n_103__55_, r_n_103__54_, r_n_103__53_, r_n_103__52_, r_n_103__51_, r_n_103__50_, r_n_103__49_, r_n_103__48_, r_n_103__47_, r_n_103__46_, r_n_103__45_, r_n_103__44_, r_n_103__43_, r_n_103__42_, r_n_103__41_, r_n_103__40_, r_n_103__39_, r_n_103__38_, r_n_103__37_, r_n_103__36_, r_n_103__35_, r_n_103__34_, r_n_103__33_, r_n_103__32_, r_n_103__31_, r_n_103__30_, r_n_103__29_, r_n_103__28_, r_n_103__27_, r_n_103__26_, r_n_103__25_, r_n_103__24_, r_n_103__23_, r_n_103__22_, r_n_103__21_, r_n_103__20_, r_n_103__19_, r_n_103__18_, r_n_103__17_, r_n_103__16_, r_n_103__15_, r_n_103__14_, r_n_103__13_, r_n_103__12_, r_n_103__11_, r_n_103__10_, r_n_103__9_, r_n_103__8_, r_n_103__7_, r_n_103__6_, r_n_103__5_, r_n_103__4_, r_n_103__3_, r_n_103__2_, r_n_103__1_, r_n_103__0_ } = (N206)? { r_104__63_, r_104__62_, r_104__61_, r_104__60_, r_104__59_, r_104__58_, r_104__57_, r_104__56_, r_104__55_, r_104__54_, r_104__53_, r_104__52_, r_104__51_, r_104__50_, r_104__49_, r_104__48_, r_104__47_, r_104__46_, r_104__45_, r_104__44_, r_104__43_, r_104__42_, r_104__41_, r_104__40_, r_104__39_, r_104__38_, r_104__37_, r_104__36_, r_104__35_, r_104__34_, r_104__33_, r_104__32_, r_104__31_, r_104__30_, r_104__29_, r_104__28_, r_104__27_, r_104__26_, r_104__25_, r_104__24_, r_104__23_, r_104__22_, r_104__21_, r_104__20_, r_104__19_, r_104__18_, r_104__17_, r_104__16_, r_104__15_, r_104__14_, r_104__13_, r_104__12_, r_104__11_, r_104__10_, r_104__9_, r_104__8_, r_104__7_, r_104__6_, r_104__5_, r_104__4_, r_104__3_, r_104__2_, r_104__1_, r_104__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N207)? data_i : 1'b0;
  assign N206 = sel_i[206];
  assign N207 = N1543;
  assign { r_n_104__63_, r_n_104__62_, r_n_104__61_, r_n_104__60_, r_n_104__59_, r_n_104__58_, r_n_104__57_, r_n_104__56_, r_n_104__55_, r_n_104__54_, r_n_104__53_, r_n_104__52_, r_n_104__51_, r_n_104__50_, r_n_104__49_, r_n_104__48_, r_n_104__47_, r_n_104__46_, r_n_104__45_, r_n_104__44_, r_n_104__43_, r_n_104__42_, r_n_104__41_, r_n_104__40_, r_n_104__39_, r_n_104__38_, r_n_104__37_, r_n_104__36_, r_n_104__35_, r_n_104__34_, r_n_104__33_, r_n_104__32_, r_n_104__31_, r_n_104__30_, r_n_104__29_, r_n_104__28_, r_n_104__27_, r_n_104__26_, r_n_104__25_, r_n_104__24_, r_n_104__23_, r_n_104__22_, r_n_104__21_, r_n_104__20_, r_n_104__19_, r_n_104__18_, r_n_104__17_, r_n_104__16_, r_n_104__15_, r_n_104__14_, r_n_104__13_, r_n_104__12_, r_n_104__11_, r_n_104__10_, r_n_104__9_, r_n_104__8_, r_n_104__7_, r_n_104__6_, r_n_104__5_, r_n_104__4_, r_n_104__3_, r_n_104__2_, r_n_104__1_, r_n_104__0_ } = (N208)? { r_105__63_, r_105__62_, r_105__61_, r_105__60_, r_105__59_, r_105__58_, r_105__57_, r_105__56_, r_105__55_, r_105__54_, r_105__53_, r_105__52_, r_105__51_, r_105__50_, r_105__49_, r_105__48_, r_105__47_, r_105__46_, r_105__45_, r_105__44_, r_105__43_, r_105__42_, r_105__41_, r_105__40_, r_105__39_, r_105__38_, r_105__37_, r_105__36_, r_105__35_, r_105__34_, r_105__33_, r_105__32_, r_105__31_, r_105__30_, r_105__29_, r_105__28_, r_105__27_, r_105__26_, r_105__25_, r_105__24_, r_105__23_, r_105__22_, r_105__21_, r_105__20_, r_105__19_, r_105__18_, r_105__17_, r_105__16_, r_105__15_, r_105__14_, r_105__13_, r_105__12_, r_105__11_, r_105__10_, r_105__9_, r_105__8_, r_105__7_, r_105__6_, r_105__5_, r_105__4_, r_105__3_, r_105__2_, r_105__1_, r_105__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N209)? data_i : 1'b0;
  assign N208 = sel_i[208];
  assign N209 = N1548;
  assign { r_n_105__63_, r_n_105__62_, r_n_105__61_, r_n_105__60_, r_n_105__59_, r_n_105__58_, r_n_105__57_, r_n_105__56_, r_n_105__55_, r_n_105__54_, r_n_105__53_, r_n_105__52_, r_n_105__51_, r_n_105__50_, r_n_105__49_, r_n_105__48_, r_n_105__47_, r_n_105__46_, r_n_105__45_, r_n_105__44_, r_n_105__43_, r_n_105__42_, r_n_105__41_, r_n_105__40_, r_n_105__39_, r_n_105__38_, r_n_105__37_, r_n_105__36_, r_n_105__35_, r_n_105__34_, r_n_105__33_, r_n_105__32_, r_n_105__31_, r_n_105__30_, r_n_105__29_, r_n_105__28_, r_n_105__27_, r_n_105__26_, r_n_105__25_, r_n_105__24_, r_n_105__23_, r_n_105__22_, r_n_105__21_, r_n_105__20_, r_n_105__19_, r_n_105__18_, r_n_105__17_, r_n_105__16_, r_n_105__15_, r_n_105__14_, r_n_105__13_, r_n_105__12_, r_n_105__11_, r_n_105__10_, r_n_105__9_, r_n_105__8_, r_n_105__7_, r_n_105__6_, r_n_105__5_, r_n_105__4_, r_n_105__3_, r_n_105__2_, r_n_105__1_, r_n_105__0_ } = (N210)? { r_106__63_, r_106__62_, r_106__61_, r_106__60_, r_106__59_, r_106__58_, r_106__57_, r_106__56_, r_106__55_, r_106__54_, r_106__53_, r_106__52_, r_106__51_, r_106__50_, r_106__49_, r_106__48_, r_106__47_, r_106__46_, r_106__45_, r_106__44_, r_106__43_, r_106__42_, r_106__41_, r_106__40_, r_106__39_, r_106__38_, r_106__37_, r_106__36_, r_106__35_, r_106__34_, r_106__33_, r_106__32_, r_106__31_, r_106__30_, r_106__29_, r_106__28_, r_106__27_, r_106__26_, r_106__25_, r_106__24_, r_106__23_, r_106__22_, r_106__21_, r_106__20_, r_106__19_, r_106__18_, r_106__17_, r_106__16_, r_106__15_, r_106__14_, r_106__13_, r_106__12_, r_106__11_, r_106__10_, r_106__9_, r_106__8_, r_106__7_, r_106__6_, r_106__5_, r_106__4_, r_106__3_, r_106__2_, r_106__1_, r_106__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N211)? data_i : 1'b0;
  assign N210 = sel_i[210];
  assign N211 = N1553;
  assign { r_n_106__63_, r_n_106__62_, r_n_106__61_, r_n_106__60_, r_n_106__59_, r_n_106__58_, r_n_106__57_, r_n_106__56_, r_n_106__55_, r_n_106__54_, r_n_106__53_, r_n_106__52_, r_n_106__51_, r_n_106__50_, r_n_106__49_, r_n_106__48_, r_n_106__47_, r_n_106__46_, r_n_106__45_, r_n_106__44_, r_n_106__43_, r_n_106__42_, r_n_106__41_, r_n_106__40_, r_n_106__39_, r_n_106__38_, r_n_106__37_, r_n_106__36_, r_n_106__35_, r_n_106__34_, r_n_106__33_, r_n_106__32_, r_n_106__31_, r_n_106__30_, r_n_106__29_, r_n_106__28_, r_n_106__27_, r_n_106__26_, r_n_106__25_, r_n_106__24_, r_n_106__23_, r_n_106__22_, r_n_106__21_, r_n_106__20_, r_n_106__19_, r_n_106__18_, r_n_106__17_, r_n_106__16_, r_n_106__15_, r_n_106__14_, r_n_106__13_, r_n_106__12_, r_n_106__11_, r_n_106__10_, r_n_106__9_, r_n_106__8_, r_n_106__7_, r_n_106__6_, r_n_106__5_, r_n_106__4_, r_n_106__3_, r_n_106__2_, r_n_106__1_, r_n_106__0_ } = (N212)? { r_107__63_, r_107__62_, r_107__61_, r_107__60_, r_107__59_, r_107__58_, r_107__57_, r_107__56_, r_107__55_, r_107__54_, r_107__53_, r_107__52_, r_107__51_, r_107__50_, r_107__49_, r_107__48_, r_107__47_, r_107__46_, r_107__45_, r_107__44_, r_107__43_, r_107__42_, r_107__41_, r_107__40_, r_107__39_, r_107__38_, r_107__37_, r_107__36_, r_107__35_, r_107__34_, r_107__33_, r_107__32_, r_107__31_, r_107__30_, r_107__29_, r_107__28_, r_107__27_, r_107__26_, r_107__25_, r_107__24_, r_107__23_, r_107__22_, r_107__21_, r_107__20_, r_107__19_, r_107__18_, r_107__17_, r_107__16_, r_107__15_, r_107__14_, r_107__13_, r_107__12_, r_107__11_, r_107__10_, r_107__9_, r_107__8_, r_107__7_, r_107__6_, r_107__5_, r_107__4_, r_107__3_, r_107__2_, r_107__1_, r_107__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N213)? data_i : 1'b0;
  assign N212 = sel_i[212];
  assign N213 = N1558;
  assign { r_n_107__63_, r_n_107__62_, r_n_107__61_, r_n_107__60_, r_n_107__59_, r_n_107__58_, r_n_107__57_, r_n_107__56_, r_n_107__55_, r_n_107__54_, r_n_107__53_, r_n_107__52_, r_n_107__51_, r_n_107__50_, r_n_107__49_, r_n_107__48_, r_n_107__47_, r_n_107__46_, r_n_107__45_, r_n_107__44_, r_n_107__43_, r_n_107__42_, r_n_107__41_, r_n_107__40_, r_n_107__39_, r_n_107__38_, r_n_107__37_, r_n_107__36_, r_n_107__35_, r_n_107__34_, r_n_107__33_, r_n_107__32_, r_n_107__31_, r_n_107__30_, r_n_107__29_, r_n_107__28_, r_n_107__27_, r_n_107__26_, r_n_107__25_, r_n_107__24_, r_n_107__23_, r_n_107__22_, r_n_107__21_, r_n_107__20_, r_n_107__19_, r_n_107__18_, r_n_107__17_, r_n_107__16_, r_n_107__15_, r_n_107__14_, r_n_107__13_, r_n_107__12_, r_n_107__11_, r_n_107__10_, r_n_107__9_, r_n_107__8_, r_n_107__7_, r_n_107__6_, r_n_107__5_, r_n_107__4_, r_n_107__3_, r_n_107__2_, r_n_107__1_, r_n_107__0_ } = (N214)? { r_108__63_, r_108__62_, r_108__61_, r_108__60_, r_108__59_, r_108__58_, r_108__57_, r_108__56_, r_108__55_, r_108__54_, r_108__53_, r_108__52_, r_108__51_, r_108__50_, r_108__49_, r_108__48_, r_108__47_, r_108__46_, r_108__45_, r_108__44_, r_108__43_, r_108__42_, r_108__41_, r_108__40_, r_108__39_, r_108__38_, r_108__37_, r_108__36_, r_108__35_, r_108__34_, r_108__33_, r_108__32_, r_108__31_, r_108__30_, r_108__29_, r_108__28_, r_108__27_, r_108__26_, r_108__25_, r_108__24_, r_108__23_, r_108__22_, r_108__21_, r_108__20_, r_108__19_, r_108__18_, r_108__17_, r_108__16_, r_108__15_, r_108__14_, r_108__13_, r_108__12_, r_108__11_, r_108__10_, r_108__9_, r_108__8_, r_108__7_, r_108__6_, r_108__5_, r_108__4_, r_108__3_, r_108__2_, r_108__1_, r_108__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N215)? data_i : 1'b0;
  assign N214 = sel_i[214];
  assign N215 = N1563;
  assign { r_n_108__63_, r_n_108__62_, r_n_108__61_, r_n_108__60_, r_n_108__59_, r_n_108__58_, r_n_108__57_, r_n_108__56_, r_n_108__55_, r_n_108__54_, r_n_108__53_, r_n_108__52_, r_n_108__51_, r_n_108__50_, r_n_108__49_, r_n_108__48_, r_n_108__47_, r_n_108__46_, r_n_108__45_, r_n_108__44_, r_n_108__43_, r_n_108__42_, r_n_108__41_, r_n_108__40_, r_n_108__39_, r_n_108__38_, r_n_108__37_, r_n_108__36_, r_n_108__35_, r_n_108__34_, r_n_108__33_, r_n_108__32_, r_n_108__31_, r_n_108__30_, r_n_108__29_, r_n_108__28_, r_n_108__27_, r_n_108__26_, r_n_108__25_, r_n_108__24_, r_n_108__23_, r_n_108__22_, r_n_108__21_, r_n_108__20_, r_n_108__19_, r_n_108__18_, r_n_108__17_, r_n_108__16_, r_n_108__15_, r_n_108__14_, r_n_108__13_, r_n_108__12_, r_n_108__11_, r_n_108__10_, r_n_108__9_, r_n_108__8_, r_n_108__7_, r_n_108__6_, r_n_108__5_, r_n_108__4_, r_n_108__3_, r_n_108__2_, r_n_108__1_, r_n_108__0_ } = (N216)? { r_109__63_, r_109__62_, r_109__61_, r_109__60_, r_109__59_, r_109__58_, r_109__57_, r_109__56_, r_109__55_, r_109__54_, r_109__53_, r_109__52_, r_109__51_, r_109__50_, r_109__49_, r_109__48_, r_109__47_, r_109__46_, r_109__45_, r_109__44_, r_109__43_, r_109__42_, r_109__41_, r_109__40_, r_109__39_, r_109__38_, r_109__37_, r_109__36_, r_109__35_, r_109__34_, r_109__33_, r_109__32_, r_109__31_, r_109__30_, r_109__29_, r_109__28_, r_109__27_, r_109__26_, r_109__25_, r_109__24_, r_109__23_, r_109__22_, r_109__21_, r_109__20_, r_109__19_, r_109__18_, r_109__17_, r_109__16_, r_109__15_, r_109__14_, r_109__13_, r_109__12_, r_109__11_, r_109__10_, r_109__9_, r_109__8_, r_109__7_, r_109__6_, r_109__5_, r_109__4_, r_109__3_, r_109__2_, r_109__1_, r_109__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N217)? data_i : 1'b0;
  assign N216 = sel_i[216];
  assign N217 = N1568;
  assign { r_n_109__63_, r_n_109__62_, r_n_109__61_, r_n_109__60_, r_n_109__59_, r_n_109__58_, r_n_109__57_, r_n_109__56_, r_n_109__55_, r_n_109__54_, r_n_109__53_, r_n_109__52_, r_n_109__51_, r_n_109__50_, r_n_109__49_, r_n_109__48_, r_n_109__47_, r_n_109__46_, r_n_109__45_, r_n_109__44_, r_n_109__43_, r_n_109__42_, r_n_109__41_, r_n_109__40_, r_n_109__39_, r_n_109__38_, r_n_109__37_, r_n_109__36_, r_n_109__35_, r_n_109__34_, r_n_109__33_, r_n_109__32_, r_n_109__31_, r_n_109__30_, r_n_109__29_, r_n_109__28_, r_n_109__27_, r_n_109__26_, r_n_109__25_, r_n_109__24_, r_n_109__23_, r_n_109__22_, r_n_109__21_, r_n_109__20_, r_n_109__19_, r_n_109__18_, r_n_109__17_, r_n_109__16_, r_n_109__15_, r_n_109__14_, r_n_109__13_, r_n_109__12_, r_n_109__11_, r_n_109__10_, r_n_109__9_, r_n_109__8_, r_n_109__7_, r_n_109__6_, r_n_109__5_, r_n_109__4_, r_n_109__3_, r_n_109__2_, r_n_109__1_, r_n_109__0_ } = (N218)? { r_110__63_, r_110__62_, r_110__61_, r_110__60_, r_110__59_, r_110__58_, r_110__57_, r_110__56_, r_110__55_, r_110__54_, r_110__53_, r_110__52_, r_110__51_, r_110__50_, r_110__49_, r_110__48_, r_110__47_, r_110__46_, r_110__45_, r_110__44_, r_110__43_, r_110__42_, r_110__41_, r_110__40_, r_110__39_, r_110__38_, r_110__37_, r_110__36_, r_110__35_, r_110__34_, r_110__33_, r_110__32_, r_110__31_, r_110__30_, r_110__29_, r_110__28_, r_110__27_, r_110__26_, r_110__25_, r_110__24_, r_110__23_, r_110__22_, r_110__21_, r_110__20_, r_110__19_, r_110__18_, r_110__17_, r_110__16_, r_110__15_, r_110__14_, r_110__13_, r_110__12_, r_110__11_, r_110__10_, r_110__9_, r_110__8_, r_110__7_, r_110__6_, r_110__5_, r_110__4_, r_110__3_, r_110__2_, r_110__1_, r_110__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N219)? data_i : 1'b0;
  assign N218 = sel_i[218];
  assign N219 = N1573;
  assign { r_n_110__63_, r_n_110__62_, r_n_110__61_, r_n_110__60_, r_n_110__59_, r_n_110__58_, r_n_110__57_, r_n_110__56_, r_n_110__55_, r_n_110__54_, r_n_110__53_, r_n_110__52_, r_n_110__51_, r_n_110__50_, r_n_110__49_, r_n_110__48_, r_n_110__47_, r_n_110__46_, r_n_110__45_, r_n_110__44_, r_n_110__43_, r_n_110__42_, r_n_110__41_, r_n_110__40_, r_n_110__39_, r_n_110__38_, r_n_110__37_, r_n_110__36_, r_n_110__35_, r_n_110__34_, r_n_110__33_, r_n_110__32_, r_n_110__31_, r_n_110__30_, r_n_110__29_, r_n_110__28_, r_n_110__27_, r_n_110__26_, r_n_110__25_, r_n_110__24_, r_n_110__23_, r_n_110__22_, r_n_110__21_, r_n_110__20_, r_n_110__19_, r_n_110__18_, r_n_110__17_, r_n_110__16_, r_n_110__15_, r_n_110__14_, r_n_110__13_, r_n_110__12_, r_n_110__11_, r_n_110__10_, r_n_110__9_, r_n_110__8_, r_n_110__7_, r_n_110__6_, r_n_110__5_, r_n_110__4_, r_n_110__3_, r_n_110__2_, r_n_110__1_, r_n_110__0_ } = (N220)? { r_111__63_, r_111__62_, r_111__61_, r_111__60_, r_111__59_, r_111__58_, r_111__57_, r_111__56_, r_111__55_, r_111__54_, r_111__53_, r_111__52_, r_111__51_, r_111__50_, r_111__49_, r_111__48_, r_111__47_, r_111__46_, r_111__45_, r_111__44_, r_111__43_, r_111__42_, r_111__41_, r_111__40_, r_111__39_, r_111__38_, r_111__37_, r_111__36_, r_111__35_, r_111__34_, r_111__33_, r_111__32_, r_111__31_, r_111__30_, r_111__29_, r_111__28_, r_111__27_, r_111__26_, r_111__25_, r_111__24_, r_111__23_, r_111__22_, r_111__21_, r_111__20_, r_111__19_, r_111__18_, r_111__17_, r_111__16_, r_111__15_, r_111__14_, r_111__13_, r_111__12_, r_111__11_, r_111__10_, r_111__9_, r_111__8_, r_111__7_, r_111__6_, r_111__5_, r_111__4_, r_111__3_, r_111__2_, r_111__1_, r_111__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N221)? data_i : 1'b0;
  assign N220 = sel_i[220];
  assign N221 = N1578;
  assign { r_n_111__63_, r_n_111__62_, r_n_111__61_, r_n_111__60_, r_n_111__59_, r_n_111__58_, r_n_111__57_, r_n_111__56_, r_n_111__55_, r_n_111__54_, r_n_111__53_, r_n_111__52_, r_n_111__51_, r_n_111__50_, r_n_111__49_, r_n_111__48_, r_n_111__47_, r_n_111__46_, r_n_111__45_, r_n_111__44_, r_n_111__43_, r_n_111__42_, r_n_111__41_, r_n_111__40_, r_n_111__39_, r_n_111__38_, r_n_111__37_, r_n_111__36_, r_n_111__35_, r_n_111__34_, r_n_111__33_, r_n_111__32_, r_n_111__31_, r_n_111__30_, r_n_111__29_, r_n_111__28_, r_n_111__27_, r_n_111__26_, r_n_111__25_, r_n_111__24_, r_n_111__23_, r_n_111__22_, r_n_111__21_, r_n_111__20_, r_n_111__19_, r_n_111__18_, r_n_111__17_, r_n_111__16_, r_n_111__15_, r_n_111__14_, r_n_111__13_, r_n_111__12_, r_n_111__11_, r_n_111__10_, r_n_111__9_, r_n_111__8_, r_n_111__7_, r_n_111__6_, r_n_111__5_, r_n_111__4_, r_n_111__3_, r_n_111__2_, r_n_111__1_, r_n_111__0_ } = (N222)? { r_112__63_, r_112__62_, r_112__61_, r_112__60_, r_112__59_, r_112__58_, r_112__57_, r_112__56_, r_112__55_, r_112__54_, r_112__53_, r_112__52_, r_112__51_, r_112__50_, r_112__49_, r_112__48_, r_112__47_, r_112__46_, r_112__45_, r_112__44_, r_112__43_, r_112__42_, r_112__41_, r_112__40_, r_112__39_, r_112__38_, r_112__37_, r_112__36_, r_112__35_, r_112__34_, r_112__33_, r_112__32_, r_112__31_, r_112__30_, r_112__29_, r_112__28_, r_112__27_, r_112__26_, r_112__25_, r_112__24_, r_112__23_, r_112__22_, r_112__21_, r_112__20_, r_112__19_, r_112__18_, r_112__17_, r_112__16_, r_112__15_, r_112__14_, r_112__13_, r_112__12_, r_112__11_, r_112__10_, r_112__9_, r_112__8_, r_112__7_, r_112__6_, r_112__5_, r_112__4_, r_112__3_, r_112__2_, r_112__1_, r_112__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N223)? data_i : 1'b0;
  assign N222 = sel_i[222];
  assign N223 = N1583;
  assign { r_n_112__63_, r_n_112__62_, r_n_112__61_, r_n_112__60_, r_n_112__59_, r_n_112__58_, r_n_112__57_, r_n_112__56_, r_n_112__55_, r_n_112__54_, r_n_112__53_, r_n_112__52_, r_n_112__51_, r_n_112__50_, r_n_112__49_, r_n_112__48_, r_n_112__47_, r_n_112__46_, r_n_112__45_, r_n_112__44_, r_n_112__43_, r_n_112__42_, r_n_112__41_, r_n_112__40_, r_n_112__39_, r_n_112__38_, r_n_112__37_, r_n_112__36_, r_n_112__35_, r_n_112__34_, r_n_112__33_, r_n_112__32_, r_n_112__31_, r_n_112__30_, r_n_112__29_, r_n_112__28_, r_n_112__27_, r_n_112__26_, r_n_112__25_, r_n_112__24_, r_n_112__23_, r_n_112__22_, r_n_112__21_, r_n_112__20_, r_n_112__19_, r_n_112__18_, r_n_112__17_, r_n_112__16_, r_n_112__15_, r_n_112__14_, r_n_112__13_, r_n_112__12_, r_n_112__11_, r_n_112__10_, r_n_112__9_, r_n_112__8_, r_n_112__7_, r_n_112__6_, r_n_112__5_, r_n_112__4_, r_n_112__3_, r_n_112__2_, r_n_112__1_, r_n_112__0_ } = (N224)? { r_113__63_, r_113__62_, r_113__61_, r_113__60_, r_113__59_, r_113__58_, r_113__57_, r_113__56_, r_113__55_, r_113__54_, r_113__53_, r_113__52_, r_113__51_, r_113__50_, r_113__49_, r_113__48_, r_113__47_, r_113__46_, r_113__45_, r_113__44_, r_113__43_, r_113__42_, r_113__41_, r_113__40_, r_113__39_, r_113__38_, r_113__37_, r_113__36_, r_113__35_, r_113__34_, r_113__33_, r_113__32_, r_113__31_, r_113__30_, r_113__29_, r_113__28_, r_113__27_, r_113__26_, r_113__25_, r_113__24_, r_113__23_, r_113__22_, r_113__21_, r_113__20_, r_113__19_, r_113__18_, r_113__17_, r_113__16_, r_113__15_, r_113__14_, r_113__13_, r_113__12_, r_113__11_, r_113__10_, r_113__9_, r_113__8_, r_113__7_, r_113__6_, r_113__5_, r_113__4_, r_113__3_, r_113__2_, r_113__1_, r_113__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N225)? data_i : 1'b0;
  assign N224 = sel_i[224];
  assign N225 = N1588;
  assign { r_n_113__63_, r_n_113__62_, r_n_113__61_, r_n_113__60_, r_n_113__59_, r_n_113__58_, r_n_113__57_, r_n_113__56_, r_n_113__55_, r_n_113__54_, r_n_113__53_, r_n_113__52_, r_n_113__51_, r_n_113__50_, r_n_113__49_, r_n_113__48_, r_n_113__47_, r_n_113__46_, r_n_113__45_, r_n_113__44_, r_n_113__43_, r_n_113__42_, r_n_113__41_, r_n_113__40_, r_n_113__39_, r_n_113__38_, r_n_113__37_, r_n_113__36_, r_n_113__35_, r_n_113__34_, r_n_113__33_, r_n_113__32_, r_n_113__31_, r_n_113__30_, r_n_113__29_, r_n_113__28_, r_n_113__27_, r_n_113__26_, r_n_113__25_, r_n_113__24_, r_n_113__23_, r_n_113__22_, r_n_113__21_, r_n_113__20_, r_n_113__19_, r_n_113__18_, r_n_113__17_, r_n_113__16_, r_n_113__15_, r_n_113__14_, r_n_113__13_, r_n_113__12_, r_n_113__11_, r_n_113__10_, r_n_113__9_, r_n_113__8_, r_n_113__7_, r_n_113__6_, r_n_113__5_, r_n_113__4_, r_n_113__3_, r_n_113__2_, r_n_113__1_, r_n_113__0_ } = (N226)? { r_114__63_, r_114__62_, r_114__61_, r_114__60_, r_114__59_, r_114__58_, r_114__57_, r_114__56_, r_114__55_, r_114__54_, r_114__53_, r_114__52_, r_114__51_, r_114__50_, r_114__49_, r_114__48_, r_114__47_, r_114__46_, r_114__45_, r_114__44_, r_114__43_, r_114__42_, r_114__41_, r_114__40_, r_114__39_, r_114__38_, r_114__37_, r_114__36_, r_114__35_, r_114__34_, r_114__33_, r_114__32_, r_114__31_, r_114__30_, r_114__29_, r_114__28_, r_114__27_, r_114__26_, r_114__25_, r_114__24_, r_114__23_, r_114__22_, r_114__21_, r_114__20_, r_114__19_, r_114__18_, r_114__17_, r_114__16_, r_114__15_, r_114__14_, r_114__13_, r_114__12_, r_114__11_, r_114__10_, r_114__9_, r_114__8_, r_114__7_, r_114__6_, r_114__5_, r_114__4_, r_114__3_, r_114__2_, r_114__1_, r_114__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N227)? data_i : 1'b0;
  assign N226 = sel_i[226];
  assign N227 = N1593;
  assign { r_n_114__63_, r_n_114__62_, r_n_114__61_, r_n_114__60_, r_n_114__59_, r_n_114__58_, r_n_114__57_, r_n_114__56_, r_n_114__55_, r_n_114__54_, r_n_114__53_, r_n_114__52_, r_n_114__51_, r_n_114__50_, r_n_114__49_, r_n_114__48_, r_n_114__47_, r_n_114__46_, r_n_114__45_, r_n_114__44_, r_n_114__43_, r_n_114__42_, r_n_114__41_, r_n_114__40_, r_n_114__39_, r_n_114__38_, r_n_114__37_, r_n_114__36_, r_n_114__35_, r_n_114__34_, r_n_114__33_, r_n_114__32_, r_n_114__31_, r_n_114__30_, r_n_114__29_, r_n_114__28_, r_n_114__27_, r_n_114__26_, r_n_114__25_, r_n_114__24_, r_n_114__23_, r_n_114__22_, r_n_114__21_, r_n_114__20_, r_n_114__19_, r_n_114__18_, r_n_114__17_, r_n_114__16_, r_n_114__15_, r_n_114__14_, r_n_114__13_, r_n_114__12_, r_n_114__11_, r_n_114__10_, r_n_114__9_, r_n_114__8_, r_n_114__7_, r_n_114__6_, r_n_114__5_, r_n_114__4_, r_n_114__3_, r_n_114__2_, r_n_114__1_, r_n_114__0_ } = (N228)? { r_115__63_, r_115__62_, r_115__61_, r_115__60_, r_115__59_, r_115__58_, r_115__57_, r_115__56_, r_115__55_, r_115__54_, r_115__53_, r_115__52_, r_115__51_, r_115__50_, r_115__49_, r_115__48_, r_115__47_, r_115__46_, r_115__45_, r_115__44_, r_115__43_, r_115__42_, r_115__41_, r_115__40_, r_115__39_, r_115__38_, r_115__37_, r_115__36_, r_115__35_, r_115__34_, r_115__33_, r_115__32_, r_115__31_, r_115__30_, r_115__29_, r_115__28_, r_115__27_, r_115__26_, r_115__25_, r_115__24_, r_115__23_, r_115__22_, r_115__21_, r_115__20_, r_115__19_, r_115__18_, r_115__17_, r_115__16_, r_115__15_, r_115__14_, r_115__13_, r_115__12_, r_115__11_, r_115__10_, r_115__9_, r_115__8_, r_115__7_, r_115__6_, r_115__5_, r_115__4_, r_115__3_, r_115__2_, r_115__1_, r_115__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N229)? data_i : 1'b0;
  assign N228 = sel_i[228];
  assign N229 = N1598;
  assign { r_n_115__63_, r_n_115__62_, r_n_115__61_, r_n_115__60_, r_n_115__59_, r_n_115__58_, r_n_115__57_, r_n_115__56_, r_n_115__55_, r_n_115__54_, r_n_115__53_, r_n_115__52_, r_n_115__51_, r_n_115__50_, r_n_115__49_, r_n_115__48_, r_n_115__47_, r_n_115__46_, r_n_115__45_, r_n_115__44_, r_n_115__43_, r_n_115__42_, r_n_115__41_, r_n_115__40_, r_n_115__39_, r_n_115__38_, r_n_115__37_, r_n_115__36_, r_n_115__35_, r_n_115__34_, r_n_115__33_, r_n_115__32_, r_n_115__31_, r_n_115__30_, r_n_115__29_, r_n_115__28_, r_n_115__27_, r_n_115__26_, r_n_115__25_, r_n_115__24_, r_n_115__23_, r_n_115__22_, r_n_115__21_, r_n_115__20_, r_n_115__19_, r_n_115__18_, r_n_115__17_, r_n_115__16_, r_n_115__15_, r_n_115__14_, r_n_115__13_, r_n_115__12_, r_n_115__11_, r_n_115__10_, r_n_115__9_, r_n_115__8_, r_n_115__7_, r_n_115__6_, r_n_115__5_, r_n_115__4_, r_n_115__3_, r_n_115__2_, r_n_115__1_, r_n_115__0_ } = (N230)? { r_116__63_, r_116__62_, r_116__61_, r_116__60_, r_116__59_, r_116__58_, r_116__57_, r_116__56_, r_116__55_, r_116__54_, r_116__53_, r_116__52_, r_116__51_, r_116__50_, r_116__49_, r_116__48_, r_116__47_, r_116__46_, r_116__45_, r_116__44_, r_116__43_, r_116__42_, r_116__41_, r_116__40_, r_116__39_, r_116__38_, r_116__37_, r_116__36_, r_116__35_, r_116__34_, r_116__33_, r_116__32_, r_116__31_, r_116__30_, r_116__29_, r_116__28_, r_116__27_, r_116__26_, r_116__25_, r_116__24_, r_116__23_, r_116__22_, r_116__21_, r_116__20_, r_116__19_, r_116__18_, r_116__17_, r_116__16_, r_116__15_, r_116__14_, r_116__13_, r_116__12_, r_116__11_, r_116__10_, r_116__9_, r_116__8_, r_116__7_, r_116__6_, r_116__5_, r_116__4_, r_116__3_, r_116__2_, r_116__1_, r_116__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N231)? data_i : 1'b0;
  assign N230 = sel_i[230];
  assign N231 = N1603;
  assign { r_n_116__63_, r_n_116__62_, r_n_116__61_, r_n_116__60_, r_n_116__59_, r_n_116__58_, r_n_116__57_, r_n_116__56_, r_n_116__55_, r_n_116__54_, r_n_116__53_, r_n_116__52_, r_n_116__51_, r_n_116__50_, r_n_116__49_, r_n_116__48_, r_n_116__47_, r_n_116__46_, r_n_116__45_, r_n_116__44_, r_n_116__43_, r_n_116__42_, r_n_116__41_, r_n_116__40_, r_n_116__39_, r_n_116__38_, r_n_116__37_, r_n_116__36_, r_n_116__35_, r_n_116__34_, r_n_116__33_, r_n_116__32_, r_n_116__31_, r_n_116__30_, r_n_116__29_, r_n_116__28_, r_n_116__27_, r_n_116__26_, r_n_116__25_, r_n_116__24_, r_n_116__23_, r_n_116__22_, r_n_116__21_, r_n_116__20_, r_n_116__19_, r_n_116__18_, r_n_116__17_, r_n_116__16_, r_n_116__15_, r_n_116__14_, r_n_116__13_, r_n_116__12_, r_n_116__11_, r_n_116__10_, r_n_116__9_, r_n_116__8_, r_n_116__7_, r_n_116__6_, r_n_116__5_, r_n_116__4_, r_n_116__3_, r_n_116__2_, r_n_116__1_, r_n_116__0_ } = (N232)? { r_117__63_, r_117__62_, r_117__61_, r_117__60_, r_117__59_, r_117__58_, r_117__57_, r_117__56_, r_117__55_, r_117__54_, r_117__53_, r_117__52_, r_117__51_, r_117__50_, r_117__49_, r_117__48_, r_117__47_, r_117__46_, r_117__45_, r_117__44_, r_117__43_, r_117__42_, r_117__41_, r_117__40_, r_117__39_, r_117__38_, r_117__37_, r_117__36_, r_117__35_, r_117__34_, r_117__33_, r_117__32_, r_117__31_, r_117__30_, r_117__29_, r_117__28_, r_117__27_, r_117__26_, r_117__25_, r_117__24_, r_117__23_, r_117__22_, r_117__21_, r_117__20_, r_117__19_, r_117__18_, r_117__17_, r_117__16_, r_117__15_, r_117__14_, r_117__13_, r_117__12_, r_117__11_, r_117__10_, r_117__9_, r_117__8_, r_117__7_, r_117__6_, r_117__5_, r_117__4_, r_117__3_, r_117__2_, r_117__1_, r_117__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N233)? data_i : 1'b0;
  assign N232 = sel_i[232];
  assign N233 = N1608;
  assign { r_n_117__63_, r_n_117__62_, r_n_117__61_, r_n_117__60_, r_n_117__59_, r_n_117__58_, r_n_117__57_, r_n_117__56_, r_n_117__55_, r_n_117__54_, r_n_117__53_, r_n_117__52_, r_n_117__51_, r_n_117__50_, r_n_117__49_, r_n_117__48_, r_n_117__47_, r_n_117__46_, r_n_117__45_, r_n_117__44_, r_n_117__43_, r_n_117__42_, r_n_117__41_, r_n_117__40_, r_n_117__39_, r_n_117__38_, r_n_117__37_, r_n_117__36_, r_n_117__35_, r_n_117__34_, r_n_117__33_, r_n_117__32_, r_n_117__31_, r_n_117__30_, r_n_117__29_, r_n_117__28_, r_n_117__27_, r_n_117__26_, r_n_117__25_, r_n_117__24_, r_n_117__23_, r_n_117__22_, r_n_117__21_, r_n_117__20_, r_n_117__19_, r_n_117__18_, r_n_117__17_, r_n_117__16_, r_n_117__15_, r_n_117__14_, r_n_117__13_, r_n_117__12_, r_n_117__11_, r_n_117__10_, r_n_117__9_, r_n_117__8_, r_n_117__7_, r_n_117__6_, r_n_117__5_, r_n_117__4_, r_n_117__3_, r_n_117__2_, r_n_117__1_, r_n_117__0_ } = (N234)? { r_118__63_, r_118__62_, r_118__61_, r_118__60_, r_118__59_, r_118__58_, r_118__57_, r_118__56_, r_118__55_, r_118__54_, r_118__53_, r_118__52_, r_118__51_, r_118__50_, r_118__49_, r_118__48_, r_118__47_, r_118__46_, r_118__45_, r_118__44_, r_118__43_, r_118__42_, r_118__41_, r_118__40_, r_118__39_, r_118__38_, r_118__37_, r_118__36_, r_118__35_, r_118__34_, r_118__33_, r_118__32_, r_118__31_, r_118__30_, r_118__29_, r_118__28_, r_118__27_, r_118__26_, r_118__25_, r_118__24_, r_118__23_, r_118__22_, r_118__21_, r_118__20_, r_118__19_, r_118__18_, r_118__17_, r_118__16_, r_118__15_, r_118__14_, r_118__13_, r_118__12_, r_118__11_, r_118__10_, r_118__9_, r_118__8_, r_118__7_, r_118__6_, r_118__5_, r_118__4_, r_118__3_, r_118__2_, r_118__1_, r_118__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N235)? data_i : 1'b0;
  assign N234 = sel_i[234];
  assign N235 = N1613;
  assign { r_n_118__63_, r_n_118__62_, r_n_118__61_, r_n_118__60_, r_n_118__59_, r_n_118__58_, r_n_118__57_, r_n_118__56_, r_n_118__55_, r_n_118__54_, r_n_118__53_, r_n_118__52_, r_n_118__51_, r_n_118__50_, r_n_118__49_, r_n_118__48_, r_n_118__47_, r_n_118__46_, r_n_118__45_, r_n_118__44_, r_n_118__43_, r_n_118__42_, r_n_118__41_, r_n_118__40_, r_n_118__39_, r_n_118__38_, r_n_118__37_, r_n_118__36_, r_n_118__35_, r_n_118__34_, r_n_118__33_, r_n_118__32_, r_n_118__31_, r_n_118__30_, r_n_118__29_, r_n_118__28_, r_n_118__27_, r_n_118__26_, r_n_118__25_, r_n_118__24_, r_n_118__23_, r_n_118__22_, r_n_118__21_, r_n_118__20_, r_n_118__19_, r_n_118__18_, r_n_118__17_, r_n_118__16_, r_n_118__15_, r_n_118__14_, r_n_118__13_, r_n_118__12_, r_n_118__11_, r_n_118__10_, r_n_118__9_, r_n_118__8_, r_n_118__7_, r_n_118__6_, r_n_118__5_, r_n_118__4_, r_n_118__3_, r_n_118__2_, r_n_118__1_, r_n_118__0_ } = (N236)? { r_119__63_, r_119__62_, r_119__61_, r_119__60_, r_119__59_, r_119__58_, r_119__57_, r_119__56_, r_119__55_, r_119__54_, r_119__53_, r_119__52_, r_119__51_, r_119__50_, r_119__49_, r_119__48_, r_119__47_, r_119__46_, r_119__45_, r_119__44_, r_119__43_, r_119__42_, r_119__41_, r_119__40_, r_119__39_, r_119__38_, r_119__37_, r_119__36_, r_119__35_, r_119__34_, r_119__33_, r_119__32_, r_119__31_, r_119__30_, r_119__29_, r_119__28_, r_119__27_, r_119__26_, r_119__25_, r_119__24_, r_119__23_, r_119__22_, r_119__21_, r_119__20_, r_119__19_, r_119__18_, r_119__17_, r_119__16_, r_119__15_, r_119__14_, r_119__13_, r_119__12_, r_119__11_, r_119__10_, r_119__9_, r_119__8_, r_119__7_, r_119__6_, r_119__5_, r_119__4_, r_119__3_, r_119__2_, r_119__1_, r_119__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N237)? data_i : 1'b0;
  assign N236 = sel_i[236];
  assign N237 = N1618;
  assign { r_n_119__63_, r_n_119__62_, r_n_119__61_, r_n_119__60_, r_n_119__59_, r_n_119__58_, r_n_119__57_, r_n_119__56_, r_n_119__55_, r_n_119__54_, r_n_119__53_, r_n_119__52_, r_n_119__51_, r_n_119__50_, r_n_119__49_, r_n_119__48_, r_n_119__47_, r_n_119__46_, r_n_119__45_, r_n_119__44_, r_n_119__43_, r_n_119__42_, r_n_119__41_, r_n_119__40_, r_n_119__39_, r_n_119__38_, r_n_119__37_, r_n_119__36_, r_n_119__35_, r_n_119__34_, r_n_119__33_, r_n_119__32_, r_n_119__31_, r_n_119__30_, r_n_119__29_, r_n_119__28_, r_n_119__27_, r_n_119__26_, r_n_119__25_, r_n_119__24_, r_n_119__23_, r_n_119__22_, r_n_119__21_, r_n_119__20_, r_n_119__19_, r_n_119__18_, r_n_119__17_, r_n_119__16_, r_n_119__15_, r_n_119__14_, r_n_119__13_, r_n_119__12_, r_n_119__11_, r_n_119__10_, r_n_119__9_, r_n_119__8_, r_n_119__7_, r_n_119__6_, r_n_119__5_, r_n_119__4_, r_n_119__3_, r_n_119__2_, r_n_119__1_, r_n_119__0_ } = (N238)? { r_120__63_, r_120__62_, r_120__61_, r_120__60_, r_120__59_, r_120__58_, r_120__57_, r_120__56_, r_120__55_, r_120__54_, r_120__53_, r_120__52_, r_120__51_, r_120__50_, r_120__49_, r_120__48_, r_120__47_, r_120__46_, r_120__45_, r_120__44_, r_120__43_, r_120__42_, r_120__41_, r_120__40_, r_120__39_, r_120__38_, r_120__37_, r_120__36_, r_120__35_, r_120__34_, r_120__33_, r_120__32_, r_120__31_, r_120__30_, r_120__29_, r_120__28_, r_120__27_, r_120__26_, r_120__25_, r_120__24_, r_120__23_, r_120__22_, r_120__21_, r_120__20_, r_120__19_, r_120__18_, r_120__17_, r_120__16_, r_120__15_, r_120__14_, r_120__13_, r_120__12_, r_120__11_, r_120__10_, r_120__9_, r_120__8_, r_120__7_, r_120__6_, r_120__5_, r_120__4_, r_120__3_, r_120__2_, r_120__1_, r_120__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N239)? data_i : 1'b0;
  assign N238 = sel_i[238];
  assign N239 = N1623;
  assign { r_n_120__63_, r_n_120__62_, r_n_120__61_, r_n_120__60_, r_n_120__59_, r_n_120__58_, r_n_120__57_, r_n_120__56_, r_n_120__55_, r_n_120__54_, r_n_120__53_, r_n_120__52_, r_n_120__51_, r_n_120__50_, r_n_120__49_, r_n_120__48_, r_n_120__47_, r_n_120__46_, r_n_120__45_, r_n_120__44_, r_n_120__43_, r_n_120__42_, r_n_120__41_, r_n_120__40_, r_n_120__39_, r_n_120__38_, r_n_120__37_, r_n_120__36_, r_n_120__35_, r_n_120__34_, r_n_120__33_, r_n_120__32_, r_n_120__31_, r_n_120__30_, r_n_120__29_, r_n_120__28_, r_n_120__27_, r_n_120__26_, r_n_120__25_, r_n_120__24_, r_n_120__23_, r_n_120__22_, r_n_120__21_, r_n_120__20_, r_n_120__19_, r_n_120__18_, r_n_120__17_, r_n_120__16_, r_n_120__15_, r_n_120__14_, r_n_120__13_, r_n_120__12_, r_n_120__11_, r_n_120__10_, r_n_120__9_, r_n_120__8_, r_n_120__7_, r_n_120__6_, r_n_120__5_, r_n_120__4_, r_n_120__3_, r_n_120__2_, r_n_120__1_, r_n_120__0_ } = (N240)? { r_121__63_, r_121__62_, r_121__61_, r_121__60_, r_121__59_, r_121__58_, r_121__57_, r_121__56_, r_121__55_, r_121__54_, r_121__53_, r_121__52_, r_121__51_, r_121__50_, r_121__49_, r_121__48_, r_121__47_, r_121__46_, r_121__45_, r_121__44_, r_121__43_, r_121__42_, r_121__41_, r_121__40_, r_121__39_, r_121__38_, r_121__37_, r_121__36_, r_121__35_, r_121__34_, r_121__33_, r_121__32_, r_121__31_, r_121__30_, r_121__29_, r_121__28_, r_121__27_, r_121__26_, r_121__25_, r_121__24_, r_121__23_, r_121__22_, r_121__21_, r_121__20_, r_121__19_, r_121__18_, r_121__17_, r_121__16_, r_121__15_, r_121__14_, r_121__13_, r_121__12_, r_121__11_, r_121__10_, r_121__9_, r_121__8_, r_121__7_, r_121__6_, r_121__5_, r_121__4_, r_121__3_, r_121__2_, r_121__1_, r_121__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N241)? data_i : 1'b0;
  assign N240 = sel_i[240];
  assign N241 = N1628;
  assign { r_n_121__63_, r_n_121__62_, r_n_121__61_, r_n_121__60_, r_n_121__59_, r_n_121__58_, r_n_121__57_, r_n_121__56_, r_n_121__55_, r_n_121__54_, r_n_121__53_, r_n_121__52_, r_n_121__51_, r_n_121__50_, r_n_121__49_, r_n_121__48_, r_n_121__47_, r_n_121__46_, r_n_121__45_, r_n_121__44_, r_n_121__43_, r_n_121__42_, r_n_121__41_, r_n_121__40_, r_n_121__39_, r_n_121__38_, r_n_121__37_, r_n_121__36_, r_n_121__35_, r_n_121__34_, r_n_121__33_, r_n_121__32_, r_n_121__31_, r_n_121__30_, r_n_121__29_, r_n_121__28_, r_n_121__27_, r_n_121__26_, r_n_121__25_, r_n_121__24_, r_n_121__23_, r_n_121__22_, r_n_121__21_, r_n_121__20_, r_n_121__19_, r_n_121__18_, r_n_121__17_, r_n_121__16_, r_n_121__15_, r_n_121__14_, r_n_121__13_, r_n_121__12_, r_n_121__11_, r_n_121__10_, r_n_121__9_, r_n_121__8_, r_n_121__7_, r_n_121__6_, r_n_121__5_, r_n_121__4_, r_n_121__3_, r_n_121__2_, r_n_121__1_, r_n_121__0_ } = (N242)? { r_122__63_, r_122__62_, r_122__61_, r_122__60_, r_122__59_, r_122__58_, r_122__57_, r_122__56_, r_122__55_, r_122__54_, r_122__53_, r_122__52_, r_122__51_, r_122__50_, r_122__49_, r_122__48_, r_122__47_, r_122__46_, r_122__45_, r_122__44_, r_122__43_, r_122__42_, r_122__41_, r_122__40_, r_122__39_, r_122__38_, r_122__37_, r_122__36_, r_122__35_, r_122__34_, r_122__33_, r_122__32_, r_122__31_, r_122__30_, r_122__29_, r_122__28_, r_122__27_, r_122__26_, r_122__25_, r_122__24_, r_122__23_, r_122__22_, r_122__21_, r_122__20_, r_122__19_, r_122__18_, r_122__17_, r_122__16_, r_122__15_, r_122__14_, r_122__13_, r_122__12_, r_122__11_, r_122__10_, r_122__9_, r_122__8_, r_122__7_, r_122__6_, r_122__5_, r_122__4_, r_122__3_, r_122__2_, r_122__1_, r_122__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N243)? data_i : 1'b0;
  assign N242 = sel_i[242];
  assign N243 = N1633;
  assign { r_n_122__63_, r_n_122__62_, r_n_122__61_, r_n_122__60_, r_n_122__59_, r_n_122__58_, r_n_122__57_, r_n_122__56_, r_n_122__55_, r_n_122__54_, r_n_122__53_, r_n_122__52_, r_n_122__51_, r_n_122__50_, r_n_122__49_, r_n_122__48_, r_n_122__47_, r_n_122__46_, r_n_122__45_, r_n_122__44_, r_n_122__43_, r_n_122__42_, r_n_122__41_, r_n_122__40_, r_n_122__39_, r_n_122__38_, r_n_122__37_, r_n_122__36_, r_n_122__35_, r_n_122__34_, r_n_122__33_, r_n_122__32_, r_n_122__31_, r_n_122__30_, r_n_122__29_, r_n_122__28_, r_n_122__27_, r_n_122__26_, r_n_122__25_, r_n_122__24_, r_n_122__23_, r_n_122__22_, r_n_122__21_, r_n_122__20_, r_n_122__19_, r_n_122__18_, r_n_122__17_, r_n_122__16_, r_n_122__15_, r_n_122__14_, r_n_122__13_, r_n_122__12_, r_n_122__11_, r_n_122__10_, r_n_122__9_, r_n_122__8_, r_n_122__7_, r_n_122__6_, r_n_122__5_, r_n_122__4_, r_n_122__3_, r_n_122__2_, r_n_122__1_, r_n_122__0_ } = (N244)? { r_123__63_, r_123__62_, r_123__61_, r_123__60_, r_123__59_, r_123__58_, r_123__57_, r_123__56_, r_123__55_, r_123__54_, r_123__53_, r_123__52_, r_123__51_, r_123__50_, r_123__49_, r_123__48_, r_123__47_, r_123__46_, r_123__45_, r_123__44_, r_123__43_, r_123__42_, r_123__41_, r_123__40_, r_123__39_, r_123__38_, r_123__37_, r_123__36_, r_123__35_, r_123__34_, r_123__33_, r_123__32_, r_123__31_, r_123__30_, r_123__29_, r_123__28_, r_123__27_, r_123__26_, r_123__25_, r_123__24_, r_123__23_, r_123__22_, r_123__21_, r_123__20_, r_123__19_, r_123__18_, r_123__17_, r_123__16_, r_123__15_, r_123__14_, r_123__13_, r_123__12_, r_123__11_, r_123__10_, r_123__9_, r_123__8_, r_123__7_, r_123__6_, r_123__5_, r_123__4_, r_123__3_, r_123__2_, r_123__1_, r_123__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N245)? data_i : 1'b0;
  assign N244 = sel_i[244];
  assign N245 = N1638;
  assign { r_n_123__63_, r_n_123__62_, r_n_123__61_, r_n_123__60_, r_n_123__59_, r_n_123__58_, r_n_123__57_, r_n_123__56_, r_n_123__55_, r_n_123__54_, r_n_123__53_, r_n_123__52_, r_n_123__51_, r_n_123__50_, r_n_123__49_, r_n_123__48_, r_n_123__47_, r_n_123__46_, r_n_123__45_, r_n_123__44_, r_n_123__43_, r_n_123__42_, r_n_123__41_, r_n_123__40_, r_n_123__39_, r_n_123__38_, r_n_123__37_, r_n_123__36_, r_n_123__35_, r_n_123__34_, r_n_123__33_, r_n_123__32_, r_n_123__31_, r_n_123__30_, r_n_123__29_, r_n_123__28_, r_n_123__27_, r_n_123__26_, r_n_123__25_, r_n_123__24_, r_n_123__23_, r_n_123__22_, r_n_123__21_, r_n_123__20_, r_n_123__19_, r_n_123__18_, r_n_123__17_, r_n_123__16_, r_n_123__15_, r_n_123__14_, r_n_123__13_, r_n_123__12_, r_n_123__11_, r_n_123__10_, r_n_123__9_, r_n_123__8_, r_n_123__7_, r_n_123__6_, r_n_123__5_, r_n_123__4_, r_n_123__3_, r_n_123__2_, r_n_123__1_, r_n_123__0_ } = (N246)? { r_124__63_, r_124__62_, r_124__61_, r_124__60_, r_124__59_, r_124__58_, r_124__57_, r_124__56_, r_124__55_, r_124__54_, r_124__53_, r_124__52_, r_124__51_, r_124__50_, r_124__49_, r_124__48_, r_124__47_, r_124__46_, r_124__45_, r_124__44_, r_124__43_, r_124__42_, r_124__41_, r_124__40_, r_124__39_, r_124__38_, r_124__37_, r_124__36_, r_124__35_, r_124__34_, r_124__33_, r_124__32_, r_124__31_, r_124__30_, r_124__29_, r_124__28_, r_124__27_, r_124__26_, r_124__25_, r_124__24_, r_124__23_, r_124__22_, r_124__21_, r_124__20_, r_124__19_, r_124__18_, r_124__17_, r_124__16_, r_124__15_, r_124__14_, r_124__13_, r_124__12_, r_124__11_, r_124__10_, r_124__9_, r_124__8_, r_124__7_, r_124__6_, r_124__5_, r_124__4_, r_124__3_, r_124__2_, r_124__1_, r_124__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N247)? data_i : 1'b0;
  assign N246 = sel_i[246];
  assign N247 = N1643;
  assign { r_n_124__63_, r_n_124__62_, r_n_124__61_, r_n_124__60_, r_n_124__59_, r_n_124__58_, r_n_124__57_, r_n_124__56_, r_n_124__55_, r_n_124__54_, r_n_124__53_, r_n_124__52_, r_n_124__51_, r_n_124__50_, r_n_124__49_, r_n_124__48_, r_n_124__47_, r_n_124__46_, r_n_124__45_, r_n_124__44_, r_n_124__43_, r_n_124__42_, r_n_124__41_, r_n_124__40_, r_n_124__39_, r_n_124__38_, r_n_124__37_, r_n_124__36_, r_n_124__35_, r_n_124__34_, r_n_124__33_, r_n_124__32_, r_n_124__31_, r_n_124__30_, r_n_124__29_, r_n_124__28_, r_n_124__27_, r_n_124__26_, r_n_124__25_, r_n_124__24_, r_n_124__23_, r_n_124__22_, r_n_124__21_, r_n_124__20_, r_n_124__19_, r_n_124__18_, r_n_124__17_, r_n_124__16_, r_n_124__15_, r_n_124__14_, r_n_124__13_, r_n_124__12_, r_n_124__11_, r_n_124__10_, r_n_124__9_, r_n_124__8_, r_n_124__7_, r_n_124__6_, r_n_124__5_, r_n_124__4_, r_n_124__3_, r_n_124__2_, r_n_124__1_, r_n_124__0_ } = (N248)? { r_125__63_, r_125__62_, r_125__61_, r_125__60_, r_125__59_, r_125__58_, r_125__57_, r_125__56_, r_125__55_, r_125__54_, r_125__53_, r_125__52_, r_125__51_, r_125__50_, r_125__49_, r_125__48_, r_125__47_, r_125__46_, r_125__45_, r_125__44_, r_125__43_, r_125__42_, r_125__41_, r_125__40_, r_125__39_, r_125__38_, r_125__37_, r_125__36_, r_125__35_, r_125__34_, r_125__33_, r_125__32_, r_125__31_, r_125__30_, r_125__29_, r_125__28_, r_125__27_, r_125__26_, r_125__25_, r_125__24_, r_125__23_, r_125__22_, r_125__21_, r_125__20_, r_125__19_, r_125__18_, r_125__17_, r_125__16_, r_125__15_, r_125__14_, r_125__13_, r_125__12_, r_125__11_, r_125__10_, r_125__9_, r_125__8_, r_125__7_, r_125__6_, r_125__5_, r_125__4_, r_125__3_, r_125__2_, r_125__1_, r_125__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N249)? data_i : 1'b0;
  assign N248 = sel_i[248];
  assign N249 = N1648;
  assign { r_n_125__63_, r_n_125__62_, r_n_125__61_, r_n_125__60_, r_n_125__59_, r_n_125__58_, r_n_125__57_, r_n_125__56_, r_n_125__55_, r_n_125__54_, r_n_125__53_, r_n_125__52_, r_n_125__51_, r_n_125__50_, r_n_125__49_, r_n_125__48_, r_n_125__47_, r_n_125__46_, r_n_125__45_, r_n_125__44_, r_n_125__43_, r_n_125__42_, r_n_125__41_, r_n_125__40_, r_n_125__39_, r_n_125__38_, r_n_125__37_, r_n_125__36_, r_n_125__35_, r_n_125__34_, r_n_125__33_, r_n_125__32_, r_n_125__31_, r_n_125__30_, r_n_125__29_, r_n_125__28_, r_n_125__27_, r_n_125__26_, r_n_125__25_, r_n_125__24_, r_n_125__23_, r_n_125__22_, r_n_125__21_, r_n_125__20_, r_n_125__19_, r_n_125__18_, r_n_125__17_, r_n_125__16_, r_n_125__15_, r_n_125__14_, r_n_125__13_, r_n_125__12_, r_n_125__11_, r_n_125__10_, r_n_125__9_, r_n_125__8_, r_n_125__7_, r_n_125__6_, r_n_125__5_, r_n_125__4_, r_n_125__3_, r_n_125__2_, r_n_125__1_, r_n_125__0_ } = (N250)? { r_126__63_, r_126__62_, r_126__61_, r_126__60_, r_126__59_, r_126__58_, r_126__57_, r_126__56_, r_126__55_, r_126__54_, r_126__53_, r_126__52_, r_126__51_, r_126__50_, r_126__49_, r_126__48_, r_126__47_, r_126__46_, r_126__45_, r_126__44_, r_126__43_, r_126__42_, r_126__41_, r_126__40_, r_126__39_, r_126__38_, r_126__37_, r_126__36_, r_126__35_, r_126__34_, r_126__33_, r_126__32_, r_126__31_, r_126__30_, r_126__29_, r_126__28_, r_126__27_, r_126__26_, r_126__25_, r_126__24_, r_126__23_, r_126__22_, r_126__21_, r_126__20_, r_126__19_, r_126__18_, r_126__17_, r_126__16_, r_126__15_, r_126__14_, r_126__13_, r_126__12_, r_126__11_, r_126__10_, r_126__9_, r_126__8_, r_126__7_, r_126__6_, r_126__5_, r_126__4_, r_126__3_, r_126__2_, r_126__1_, r_126__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N251)? data_i : 1'b0;
  assign N250 = sel_i[250];
  assign N251 = N1653;
  assign { r_n_126__63_, r_n_126__62_, r_n_126__61_, r_n_126__60_, r_n_126__59_, r_n_126__58_, r_n_126__57_, r_n_126__56_, r_n_126__55_, r_n_126__54_, r_n_126__53_, r_n_126__52_, r_n_126__51_, r_n_126__50_, r_n_126__49_, r_n_126__48_, r_n_126__47_, r_n_126__46_, r_n_126__45_, r_n_126__44_, r_n_126__43_, r_n_126__42_, r_n_126__41_, r_n_126__40_, r_n_126__39_, r_n_126__38_, r_n_126__37_, r_n_126__36_, r_n_126__35_, r_n_126__34_, r_n_126__33_, r_n_126__32_, r_n_126__31_, r_n_126__30_, r_n_126__29_, r_n_126__28_, r_n_126__27_, r_n_126__26_, r_n_126__25_, r_n_126__24_, r_n_126__23_, r_n_126__22_, r_n_126__21_, r_n_126__20_, r_n_126__19_, r_n_126__18_, r_n_126__17_, r_n_126__16_, r_n_126__15_, r_n_126__14_, r_n_126__13_, r_n_126__12_, r_n_126__11_, r_n_126__10_, r_n_126__9_, r_n_126__8_, r_n_126__7_, r_n_126__6_, r_n_126__5_, r_n_126__4_, r_n_126__3_, r_n_126__2_, r_n_126__1_, r_n_126__0_ } = (N252)? { r_127__63_, r_127__62_, r_127__61_, r_127__60_, r_127__59_, r_127__58_, r_127__57_, r_127__56_, r_127__55_, r_127__54_, r_127__53_, r_127__52_, r_127__51_, r_127__50_, r_127__49_, r_127__48_, r_127__47_, r_127__46_, r_127__45_, r_127__44_, r_127__43_, r_127__42_, r_127__41_, r_127__40_, r_127__39_, r_127__38_, r_127__37_, r_127__36_, r_127__35_, r_127__34_, r_127__33_, r_127__32_, r_127__31_, r_127__30_, r_127__29_, r_127__28_, r_127__27_, r_127__26_, r_127__25_, r_127__24_, r_127__23_, r_127__22_, r_127__21_, r_127__20_, r_127__19_, r_127__18_, r_127__17_, r_127__16_, r_127__15_, r_127__14_, r_127__13_, r_127__12_, r_127__11_, r_127__10_, r_127__9_, r_127__8_, r_127__7_, r_127__6_, r_127__5_, r_127__4_, r_127__3_, r_127__2_, r_127__1_, r_127__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N253)? data_i : 1'b0;
  assign N252 = sel_i[252];
  assign N253 = N1658;
  assign { r_n_127__63_, r_n_127__62_, r_n_127__61_, r_n_127__60_, r_n_127__59_, r_n_127__58_, r_n_127__57_, r_n_127__56_, r_n_127__55_, r_n_127__54_, r_n_127__53_, r_n_127__52_, r_n_127__51_, r_n_127__50_, r_n_127__49_, r_n_127__48_, r_n_127__47_, r_n_127__46_, r_n_127__45_, r_n_127__44_, r_n_127__43_, r_n_127__42_, r_n_127__41_, r_n_127__40_, r_n_127__39_, r_n_127__38_, r_n_127__37_, r_n_127__36_, r_n_127__35_, r_n_127__34_, r_n_127__33_, r_n_127__32_, r_n_127__31_, r_n_127__30_, r_n_127__29_, r_n_127__28_, r_n_127__27_, r_n_127__26_, r_n_127__25_, r_n_127__24_, r_n_127__23_, r_n_127__22_, r_n_127__21_, r_n_127__20_, r_n_127__19_, r_n_127__18_, r_n_127__17_, r_n_127__16_, r_n_127__15_, r_n_127__14_, r_n_127__13_, r_n_127__12_, r_n_127__11_, r_n_127__10_, r_n_127__9_, r_n_127__8_, r_n_127__7_, r_n_127__6_, r_n_127__5_, r_n_127__4_, r_n_127__3_, r_n_127__2_, r_n_127__1_, r_n_127__0_ } = (N254)? { r_128__63_, r_128__62_, r_128__61_, r_128__60_, r_128__59_, r_128__58_, r_128__57_, r_128__56_, r_128__55_, r_128__54_, r_128__53_, r_128__52_, r_128__51_, r_128__50_, r_128__49_, r_128__48_, r_128__47_, r_128__46_, r_128__45_, r_128__44_, r_128__43_, r_128__42_, r_128__41_, r_128__40_, r_128__39_, r_128__38_, r_128__37_, r_128__36_, r_128__35_, r_128__34_, r_128__33_, r_128__32_, r_128__31_, r_128__30_, r_128__29_, r_128__28_, r_128__27_, r_128__26_, r_128__25_, r_128__24_, r_128__23_, r_128__22_, r_128__21_, r_128__20_, r_128__19_, r_128__18_, r_128__17_, r_128__16_, r_128__15_, r_128__14_, r_128__13_, r_128__12_, r_128__11_, r_128__10_, r_128__9_, r_128__8_, r_128__7_, r_128__6_, r_128__5_, r_128__4_, r_128__3_, r_128__2_, r_128__1_, r_128__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N255)? data_i : 1'b0;
  assign N254 = sel_i[254];
  assign N255 = N1663;
  assign { r_n_128__63_, r_n_128__62_, r_n_128__61_, r_n_128__60_, r_n_128__59_, r_n_128__58_, r_n_128__57_, r_n_128__56_, r_n_128__55_, r_n_128__54_, r_n_128__53_, r_n_128__52_, r_n_128__51_, r_n_128__50_, r_n_128__49_, r_n_128__48_, r_n_128__47_, r_n_128__46_, r_n_128__45_, r_n_128__44_, r_n_128__43_, r_n_128__42_, r_n_128__41_, r_n_128__40_, r_n_128__39_, r_n_128__38_, r_n_128__37_, r_n_128__36_, r_n_128__35_, r_n_128__34_, r_n_128__33_, r_n_128__32_, r_n_128__31_, r_n_128__30_, r_n_128__29_, r_n_128__28_, r_n_128__27_, r_n_128__26_, r_n_128__25_, r_n_128__24_, r_n_128__23_, r_n_128__22_, r_n_128__21_, r_n_128__20_, r_n_128__19_, r_n_128__18_, r_n_128__17_, r_n_128__16_, r_n_128__15_, r_n_128__14_, r_n_128__13_, r_n_128__12_, r_n_128__11_, r_n_128__10_, r_n_128__9_, r_n_128__8_, r_n_128__7_, r_n_128__6_, r_n_128__5_, r_n_128__4_, r_n_128__3_, r_n_128__2_, r_n_128__1_, r_n_128__0_ } = (N256)? { r_129__63_, r_129__62_, r_129__61_, r_129__60_, r_129__59_, r_129__58_, r_129__57_, r_129__56_, r_129__55_, r_129__54_, r_129__53_, r_129__52_, r_129__51_, r_129__50_, r_129__49_, r_129__48_, r_129__47_, r_129__46_, r_129__45_, r_129__44_, r_129__43_, r_129__42_, r_129__41_, r_129__40_, r_129__39_, r_129__38_, r_129__37_, r_129__36_, r_129__35_, r_129__34_, r_129__33_, r_129__32_, r_129__31_, r_129__30_, r_129__29_, r_129__28_, r_129__27_, r_129__26_, r_129__25_, r_129__24_, r_129__23_, r_129__22_, r_129__21_, r_129__20_, r_129__19_, r_129__18_, r_129__17_, r_129__16_, r_129__15_, r_129__14_, r_129__13_, r_129__12_, r_129__11_, r_129__10_, r_129__9_, r_129__8_, r_129__7_, r_129__6_, r_129__5_, r_129__4_, r_129__3_, r_129__2_, r_129__1_, r_129__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N257)? data_i : 1'b0;
  assign N256 = sel_i[256];
  assign N257 = N1668;
  assign { r_n_129__63_, r_n_129__62_, r_n_129__61_, r_n_129__60_, r_n_129__59_, r_n_129__58_, r_n_129__57_, r_n_129__56_, r_n_129__55_, r_n_129__54_, r_n_129__53_, r_n_129__52_, r_n_129__51_, r_n_129__50_, r_n_129__49_, r_n_129__48_, r_n_129__47_, r_n_129__46_, r_n_129__45_, r_n_129__44_, r_n_129__43_, r_n_129__42_, r_n_129__41_, r_n_129__40_, r_n_129__39_, r_n_129__38_, r_n_129__37_, r_n_129__36_, r_n_129__35_, r_n_129__34_, r_n_129__33_, r_n_129__32_, r_n_129__31_, r_n_129__30_, r_n_129__29_, r_n_129__28_, r_n_129__27_, r_n_129__26_, r_n_129__25_, r_n_129__24_, r_n_129__23_, r_n_129__22_, r_n_129__21_, r_n_129__20_, r_n_129__19_, r_n_129__18_, r_n_129__17_, r_n_129__16_, r_n_129__15_, r_n_129__14_, r_n_129__13_, r_n_129__12_, r_n_129__11_, r_n_129__10_, r_n_129__9_, r_n_129__8_, r_n_129__7_, r_n_129__6_, r_n_129__5_, r_n_129__4_, r_n_129__3_, r_n_129__2_, r_n_129__1_, r_n_129__0_ } = (N258)? { r_130__63_, r_130__62_, r_130__61_, r_130__60_, r_130__59_, r_130__58_, r_130__57_, r_130__56_, r_130__55_, r_130__54_, r_130__53_, r_130__52_, r_130__51_, r_130__50_, r_130__49_, r_130__48_, r_130__47_, r_130__46_, r_130__45_, r_130__44_, r_130__43_, r_130__42_, r_130__41_, r_130__40_, r_130__39_, r_130__38_, r_130__37_, r_130__36_, r_130__35_, r_130__34_, r_130__33_, r_130__32_, r_130__31_, r_130__30_, r_130__29_, r_130__28_, r_130__27_, r_130__26_, r_130__25_, r_130__24_, r_130__23_, r_130__22_, r_130__21_, r_130__20_, r_130__19_, r_130__18_, r_130__17_, r_130__16_, r_130__15_, r_130__14_, r_130__13_, r_130__12_, r_130__11_, r_130__10_, r_130__9_, r_130__8_, r_130__7_, r_130__6_, r_130__5_, r_130__4_, r_130__3_, r_130__2_, r_130__1_, r_130__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N259)? data_i : 1'b0;
  assign N258 = sel_i[258];
  assign N259 = N1673;
  assign { r_n_130__63_, r_n_130__62_, r_n_130__61_, r_n_130__60_, r_n_130__59_, r_n_130__58_, r_n_130__57_, r_n_130__56_, r_n_130__55_, r_n_130__54_, r_n_130__53_, r_n_130__52_, r_n_130__51_, r_n_130__50_, r_n_130__49_, r_n_130__48_, r_n_130__47_, r_n_130__46_, r_n_130__45_, r_n_130__44_, r_n_130__43_, r_n_130__42_, r_n_130__41_, r_n_130__40_, r_n_130__39_, r_n_130__38_, r_n_130__37_, r_n_130__36_, r_n_130__35_, r_n_130__34_, r_n_130__33_, r_n_130__32_, r_n_130__31_, r_n_130__30_, r_n_130__29_, r_n_130__28_, r_n_130__27_, r_n_130__26_, r_n_130__25_, r_n_130__24_, r_n_130__23_, r_n_130__22_, r_n_130__21_, r_n_130__20_, r_n_130__19_, r_n_130__18_, r_n_130__17_, r_n_130__16_, r_n_130__15_, r_n_130__14_, r_n_130__13_, r_n_130__12_, r_n_130__11_, r_n_130__10_, r_n_130__9_, r_n_130__8_, r_n_130__7_, r_n_130__6_, r_n_130__5_, r_n_130__4_, r_n_130__3_, r_n_130__2_, r_n_130__1_, r_n_130__0_ } = (N260)? { r_131__63_, r_131__62_, r_131__61_, r_131__60_, r_131__59_, r_131__58_, r_131__57_, r_131__56_, r_131__55_, r_131__54_, r_131__53_, r_131__52_, r_131__51_, r_131__50_, r_131__49_, r_131__48_, r_131__47_, r_131__46_, r_131__45_, r_131__44_, r_131__43_, r_131__42_, r_131__41_, r_131__40_, r_131__39_, r_131__38_, r_131__37_, r_131__36_, r_131__35_, r_131__34_, r_131__33_, r_131__32_, r_131__31_, r_131__30_, r_131__29_, r_131__28_, r_131__27_, r_131__26_, r_131__25_, r_131__24_, r_131__23_, r_131__22_, r_131__21_, r_131__20_, r_131__19_, r_131__18_, r_131__17_, r_131__16_, r_131__15_, r_131__14_, r_131__13_, r_131__12_, r_131__11_, r_131__10_, r_131__9_, r_131__8_, r_131__7_, r_131__6_, r_131__5_, r_131__4_, r_131__3_, r_131__2_, r_131__1_, r_131__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N261)? data_i : 1'b0;
  assign N260 = sel_i[260];
  assign N261 = N1678;
  assign { r_n_131__63_, r_n_131__62_, r_n_131__61_, r_n_131__60_, r_n_131__59_, r_n_131__58_, r_n_131__57_, r_n_131__56_, r_n_131__55_, r_n_131__54_, r_n_131__53_, r_n_131__52_, r_n_131__51_, r_n_131__50_, r_n_131__49_, r_n_131__48_, r_n_131__47_, r_n_131__46_, r_n_131__45_, r_n_131__44_, r_n_131__43_, r_n_131__42_, r_n_131__41_, r_n_131__40_, r_n_131__39_, r_n_131__38_, r_n_131__37_, r_n_131__36_, r_n_131__35_, r_n_131__34_, r_n_131__33_, r_n_131__32_, r_n_131__31_, r_n_131__30_, r_n_131__29_, r_n_131__28_, r_n_131__27_, r_n_131__26_, r_n_131__25_, r_n_131__24_, r_n_131__23_, r_n_131__22_, r_n_131__21_, r_n_131__20_, r_n_131__19_, r_n_131__18_, r_n_131__17_, r_n_131__16_, r_n_131__15_, r_n_131__14_, r_n_131__13_, r_n_131__12_, r_n_131__11_, r_n_131__10_, r_n_131__9_, r_n_131__8_, r_n_131__7_, r_n_131__6_, r_n_131__5_, r_n_131__4_, r_n_131__3_, r_n_131__2_, r_n_131__1_, r_n_131__0_ } = (N262)? { r_132__63_, r_132__62_, r_132__61_, r_132__60_, r_132__59_, r_132__58_, r_132__57_, r_132__56_, r_132__55_, r_132__54_, r_132__53_, r_132__52_, r_132__51_, r_132__50_, r_132__49_, r_132__48_, r_132__47_, r_132__46_, r_132__45_, r_132__44_, r_132__43_, r_132__42_, r_132__41_, r_132__40_, r_132__39_, r_132__38_, r_132__37_, r_132__36_, r_132__35_, r_132__34_, r_132__33_, r_132__32_, r_132__31_, r_132__30_, r_132__29_, r_132__28_, r_132__27_, r_132__26_, r_132__25_, r_132__24_, r_132__23_, r_132__22_, r_132__21_, r_132__20_, r_132__19_, r_132__18_, r_132__17_, r_132__16_, r_132__15_, r_132__14_, r_132__13_, r_132__12_, r_132__11_, r_132__10_, r_132__9_, r_132__8_, r_132__7_, r_132__6_, r_132__5_, r_132__4_, r_132__3_, r_132__2_, r_132__1_, r_132__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N263)? data_i : 1'b0;
  assign N262 = sel_i[262];
  assign N263 = N1683;
  assign { r_n_132__63_, r_n_132__62_, r_n_132__61_, r_n_132__60_, r_n_132__59_, r_n_132__58_, r_n_132__57_, r_n_132__56_, r_n_132__55_, r_n_132__54_, r_n_132__53_, r_n_132__52_, r_n_132__51_, r_n_132__50_, r_n_132__49_, r_n_132__48_, r_n_132__47_, r_n_132__46_, r_n_132__45_, r_n_132__44_, r_n_132__43_, r_n_132__42_, r_n_132__41_, r_n_132__40_, r_n_132__39_, r_n_132__38_, r_n_132__37_, r_n_132__36_, r_n_132__35_, r_n_132__34_, r_n_132__33_, r_n_132__32_, r_n_132__31_, r_n_132__30_, r_n_132__29_, r_n_132__28_, r_n_132__27_, r_n_132__26_, r_n_132__25_, r_n_132__24_, r_n_132__23_, r_n_132__22_, r_n_132__21_, r_n_132__20_, r_n_132__19_, r_n_132__18_, r_n_132__17_, r_n_132__16_, r_n_132__15_, r_n_132__14_, r_n_132__13_, r_n_132__12_, r_n_132__11_, r_n_132__10_, r_n_132__9_, r_n_132__8_, r_n_132__7_, r_n_132__6_, r_n_132__5_, r_n_132__4_, r_n_132__3_, r_n_132__2_, r_n_132__1_, r_n_132__0_ } = (N264)? { r_133__63_, r_133__62_, r_133__61_, r_133__60_, r_133__59_, r_133__58_, r_133__57_, r_133__56_, r_133__55_, r_133__54_, r_133__53_, r_133__52_, r_133__51_, r_133__50_, r_133__49_, r_133__48_, r_133__47_, r_133__46_, r_133__45_, r_133__44_, r_133__43_, r_133__42_, r_133__41_, r_133__40_, r_133__39_, r_133__38_, r_133__37_, r_133__36_, r_133__35_, r_133__34_, r_133__33_, r_133__32_, r_133__31_, r_133__30_, r_133__29_, r_133__28_, r_133__27_, r_133__26_, r_133__25_, r_133__24_, r_133__23_, r_133__22_, r_133__21_, r_133__20_, r_133__19_, r_133__18_, r_133__17_, r_133__16_, r_133__15_, r_133__14_, r_133__13_, r_133__12_, r_133__11_, r_133__10_, r_133__9_, r_133__8_, r_133__7_, r_133__6_, r_133__5_, r_133__4_, r_133__3_, r_133__2_, r_133__1_, r_133__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N265)? data_i : 1'b0;
  assign N264 = sel_i[264];
  assign N265 = N1688;
  assign { r_n_133__63_, r_n_133__62_, r_n_133__61_, r_n_133__60_, r_n_133__59_, r_n_133__58_, r_n_133__57_, r_n_133__56_, r_n_133__55_, r_n_133__54_, r_n_133__53_, r_n_133__52_, r_n_133__51_, r_n_133__50_, r_n_133__49_, r_n_133__48_, r_n_133__47_, r_n_133__46_, r_n_133__45_, r_n_133__44_, r_n_133__43_, r_n_133__42_, r_n_133__41_, r_n_133__40_, r_n_133__39_, r_n_133__38_, r_n_133__37_, r_n_133__36_, r_n_133__35_, r_n_133__34_, r_n_133__33_, r_n_133__32_, r_n_133__31_, r_n_133__30_, r_n_133__29_, r_n_133__28_, r_n_133__27_, r_n_133__26_, r_n_133__25_, r_n_133__24_, r_n_133__23_, r_n_133__22_, r_n_133__21_, r_n_133__20_, r_n_133__19_, r_n_133__18_, r_n_133__17_, r_n_133__16_, r_n_133__15_, r_n_133__14_, r_n_133__13_, r_n_133__12_, r_n_133__11_, r_n_133__10_, r_n_133__9_, r_n_133__8_, r_n_133__7_, r_n_133__6_, r_n_133__5_, r_n_133__4_, r_n_133__3_, r_n_133__2_, r_n_133__1_, r_n_133__0_ } = (N266)? { r_134__63_, r_134__62_, r_134__61_, r_134__60_, r_134__59_, r_134__58_, r_134__57_, r_134__56_, r_134__55_, r_134__54_, r_134__53_, r_134__52_, r_134__51_, r_134__50_, r_134__49_, r_134__48_, r_134__47_, r_134__46_, r_134__45_, r_134__44_, r_134__43_, r_134__42_, r_134__41_, r_134__40_, r_134__39_, r_134__38_, r_134__37_, r_134__36_, r_134__35_, r_134__34_, r_134__33_, r_134__32_, r_134__31_, r_134__30_, r_134__29_, r_134__28_, r_134__27_, r_134__26_, r_134__25_, r_134__24_, r_134__23_, r_134__22_, r_134__21_, r_134__20_, r_134__19_, r_134__18_, r_134__17_, r_134__16_, r_134__15_, r_134__14_, r_134__13_, r_134__12_, r_134__11_, r_134__10_, r_134__9_, r_134__8_, r_134__7_, r_134__6_, r_134__5_, r_134__4_, r_134__3_, r_134__2_, r_134__1_, r_134__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N267)? data_i : 1'b0;
  assign N266 = sel_i[266];
  assign N267 = N1693;
  assign { r_n_134__63_, r_n_134__62_, r_n_134__61_, r_n_134__60_, r_n_134__59_, r_n_134__58_, r_n_134__57_, r_n_134__56_, r_n_134__55_, r_n_134__54_, r_n_134__53_, r_n_134__52_, r_n_134__51_, r_n_134__50_, r_n_134__49_, r_n_134__48_, r_n_134__47_, r_n_134__46_, r_n_134__45_, r_n_134__44_, r_n_134__43_, r_n_134__42_, r_n_134__41_, r_n_134__40_, r_n_134__39_, r_n_134__38_, r_n_134__37_, r_n_134__36_, r_n_134__35_, r_n_134__34_, r_n_134__33_, r_n_134__32_, r_n_134__31_, r_n_134__30_, r_n_134__29_, r_n_134__28_, r_n_134__27_, r_n_134__26_, r_n_134__25_, r_n_134__24_, r_n_134__23_, r_n_134__22_, r_n_134__21_, r_n_134__20_, r_n_134__19_, r_n_134__18_, r_n_134__17_, r_n_134__16_, r_n_134__15_, r_n_134__14_, r_n_134__13_, r_n_134__12_, r_n_134__11_, r_n_134__10_, r_n_134__9_, r_n_134__8_, r_n_134__7_, r_n_134__6_, r_n_134__5_, r_n_134__4_, r_n_134__3_, r_n_134__2_, r_n_134__1_, r_n_134__0_ } = (N268)? { r_135__63_, r_135__62_, r_135__61_, r_135__60_, r_135__59_, r_135__58_, r_135__57_, r_135__56_, r_135__55_, r_135__54_, r_135__53_, r_135__52_, r_135__51_, r_135__50_, r_135__49_, r_135__48_, r_135__47_, r_135__46_, r_135__45_, r_135__44_, r_135__43_, r_135__42_, r_135__41_, r_135__40_, r_135__39_, r_135__38_, r_135__37_, r_135__36_, r_135__35_, r_135__34_, r_135__33_, r_135__32_, r_135__31_, r_135__30_, r_135__29_, r_135__28_, r_135__27_, r_135__26_, r_135__25_, r_135__24_, r_135__23_, r_135__22_, r_135__21_, r_135__20_, r_135__19_, r_135__18_, r_135__17_, r_135__16_, r_135__15_, r_135__14_, r_135__13_, r_135__12_, r_135__11_, r_135__10_, r_135__9_, r_135__8_, r_135__7_, r_135__6_, r_135__5_, r_135__4_, r_135__3_, r_135__2_, r_135__1_, r_135__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N269)? data_i : 1'b0;
  assign N268 = sel_i[268];
  assign N269 = N1698;
  assign { r_n_135__63_, r_n_135__62_, r_n_135__61_, r_n_135__60_, r_n_135__59_, r_n_135__58_, r_n_135__57_, r_n_135__56_, r_n_135__55_, r_n_135__54_, r_n_135__53_, r_n_135__52_, r_n_135__51_, r_n_135__50_, r_n_135__49_, r_n_135__48_, r_n_135__47_, r_n_135__46_, r_n_135__45_, r_n_135__44_, r_n_135__43_, r_n_135__42_, r_n_135__41_, r_n_135__40_, r_n_135__39_, r_n_135__38_, r_n_135__37_, r_n_135__36_, r_n_135__35_, r_n_135__34_, r_n_135__33_, r_n_135__32_, r_n_135__31_, r_n_135__30_, r_n_135__29_, r_n_135__28_, r_n_135__27_, r_n_135__26_, r_n_135__25_, r_n_135__24_, r_n_135__23_, r_n_135__22_, r_n_135__21_, r_n_135__20_, r_n_135__19_, r_n_135__18_, r_n_135__17_, r_n_135__16_, r_n_135__15_, r_n_135__14_, r_n_135__13_, r_n_135__12_, r_n_135__11_, r_n_135__10_, r_n_135__9_, r_n_135__8_, r_n_135__7_, r_n_135__6_, r_n_135__5_, r_n_135__4_, r_n_135__3_, r_n_135__2_, r_n_135__1_, r_n_135__0_ } = (N270)? { r_136__63_, r_136__62_, r_136__61_, r_136__60_, r_136__59_, r_136__58_, r_136__57_, r_136__56_, r_136__55_, r_136__54_, r_136__53_, r_136__52_, r_136__51_, r_136__50_, r_136__49_, r_136__48_, r_136__47_, r_136__46_, r_136__45_, r_136__44_, r_136__43_, r_136__42_, r_136__41_, r_136__40_, r_136__39_, r_136__38_, r_136__37_, r_136__36_, r_136__35_, r_136__34_, r_136__33_, r_136__32_, r_136__31_, r_136__30_, r_136__29_, r_136__28_, r_136__27_, r_136__26_, r_136__25_, r_136__24_, r_136__23_, r_136__22_, r_136__21_, r_136__20_, r_136__19_, r_136__18_, r_136__17_, r_136__16_, r_136__15_, r_136__14_, r_136__13_, r_136__12_, r_136__11_, r_136__10_, r_136__9_, r_136__8_, r_136__7_, r_136__6_, r_136__5_, r_136__4_, r_136__3_, r_136__2_, r_136__1_, r_136__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N271)? data_i : 1'b0;
  assign N270 = sel_i[270];
  assign N271 = N1703;
  assign { r_n_136__63_, r_n_136__62_, r_n_136__61_, r_n_136__60_, r_n_136__59_, r_n_136__58_, r_n_136__57_, r_n_136__56_, r_n_136__55_, r_n_136__54_, r_n_136__53_, r_n_136__52_, r_n_136__51_, r_n_136__50_, r_n_136__49_, r_n_136__48_, r_n_136__47_, r_n_136__46_, r_n_136__45_, r_n_136__44_, r_n_136__43_, r_n_136__42_, r_n_136__41_, r_n_136__40_, r_n_136__39_, r_n_136__38_, r_n_136__37_, r_n_136__36_, r_n_136__35_, r_n_136__34_, r_n_136__33_, r_n_136__32_, r_n_136__31_, r_n_136__30_, r_n_136__29_, r_n_136__28_, r_n_136__27_, r_n_136__26_, r_n_136__25_, r_n_136__24_, r_n_136__23_, r_n_136__22_, r_n_136__21_, r_n_136__20_, r_n_136__19_, r_n_136__18_, r_n_136__17_, r_n_136__16_, r_n_136__15_, r_n_136__14_, r_n_136__13_, r_n_136__12_, r_n_136__11_, r_n_136__10_, r_n_136__9_, r_n_136__8_, r_n_136__7_, r_n_136__6_, r_n_136__5_, r_n_136__4_, r_n_136__3_, r_n_136__2_, r_n_136__1_, r_n_136__0_ } = (N272)? { r_137__63_, r_137__62_, r_137__61_, r_137__60_, r_137__59_, r_137__58_, r_137__57_, r_137__56_, r_137__55_, r_137__54_, r_137__53_, r_137__52_, r_137__51_, r_137__50_, r_137__49_, r_137__48_, r_137__47_, r_137__46_, r_137__45_, r_137__44_, r_137__43_, r_137__42_, r_137__41_, r_137__40_, r_137__39_, r_137__38_, r_137__37_, r_137__36_, r_137__35_, r_137__34_, r_137__33_, r_137__32_, r_137__31_, r_137__30_, r_137__29_, r_137__28_, r_137__27_, r_137__26_, r_137__25_, r_137__24_, r_137__23_, r_137__22_, r_137__21_, r_137__20_, r_137__19_, r_137__18_, r_137__17_, r_137__16_, r_137__15_, r_137__14_, r_137__13_, r_137__12_, r_137__11_, r_137__10_, r_137__9_, r_137__8_, r_137__7_, r_137__6_, r_137__5_, r_137__4_, r_137__3_, r_137__2_, r_137__1_, r_137__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N273)? data_i : 1'b0;
  assign N272 = sel_i[272];
  assign N273 = N1708;
  assign { r_n_137__63_, r_n_137__62_, r_n_137__61_, r_n_137__60_, r_n_137__59_, r_n_137__58_, r_n_137__57_, r_n_137__56_, r_n_137__55_, r_n_137__54_, r_n_137__53_, r_n_137__52_, r_n_137__51_, r_n_137__50_, r_n_137__49_, r_n_137__48_, r_n_137__47_, r_n_137__46_, r_n_137__45_, r_n_137__44_, r_n_137__43_, r_n_137__42_, r_n_137__41_, r_n_137__40_, r_n_137__39_, r_n_137__38_, r_n_137__37_, r_n_137__36_, r_n_137__35_, r_n_137__34_, r_n_137__33_, r_n_137__32_, r_n_137__31_, r_n_137__30_, r_n_137__29_, r_n_137__28_, r_n_137__27_, r_n_137__26_, r_n_137__25_, r_n_137__24_, r_n_137__23_, r_n_137__22_, r_n_137__21_, r_n_137__20_, r_n_137__19_, r_n_137__18_, r_n_137__17_, r_n_137__16_, r_n_137__15_, r_n_137__14_, r_n_137__13_, r_n_137__12_, r_n_137__11_, r_n_137__10_, r_n_137__9_, r_n_137__8_, r_n_137__7_, r_n_137__6_, r_n_137__5_, r_n_137__4_, r_n_137__3_, r_n_137__2_, r_n_137__1_, r_n_137__0_ } = (N274)? { r_138__63_, r_138__62_, r_138__61_, r_138__60_, r_138__59_, r_138__58_, r_138__57_, r_138__56_, r_138__55_, r_138__54_, r_138__53_, r_138__52_, r_138__51_, r_138__50_, r_138__49_, r_138__48_, r_138__47_, r_138__46_, r_138__45_, r_138__44_, r_138__43_, r_138__42_, r_138__41_, r_138__40_, r_138__39_, r_138__38_, r_138__37_, r_138__36_, r_138__35_, r_138__34_, r_138__33_, r_138__32_, r_138__31_, r_138__30_, r_138__29_, r_138__28_, r_138__27_, r_138__26_, r_138__25_, r_138__24_, r_138__23_, r_138__22_, r_138__21_, r_138__20_, r_138__19_, r_138__18_, r_138__17_, r_138__16_, r_138__15_, r_138__14_, r_138__13_, r_138__12_, r_138__11_, r_138__10_, r_138__9_, r_138__8_, r_138__7_, r_138__6_, r_138__5_, r_138__4_, r_138__3_, r_138__2_, r_138__1_, r_138__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N275)? data_i : 1'b0;
  assign N274 = sel_i[274];
  assign N275 = N1713;
  assign { r_n_138__63_, r_n_138__62_, r_n_138__61_, r_n_138__60_, r_n_138__59_, r_n_138__58_, r_n_138__57_, r_n_138__56_, r_n_138__55_, r_n_138__54_, r_n_138__53_, r_n_138__52_, r_n_138__51_, r_n_138__50_, r_n_138__49_, r_n_138__48_, r_n_138__47_, r_n_138__46_, r_n_138__45_, r_n_138__44_, r_n_138__43_, r_n_138__42_, r_n_138__41_, r_n_138__40_, r_n_138__39_, r_n_138__38_, r_n_138__37_, r_n_138__36_, r_n_138__35_, r_n_138__34_, r_n_138__33_, r_n_138__32_, r_n_138__31_, r_n_138__30_, r_n_138__29_, r_n_138__28_, r_n_138__27_, r_n_138__26_, r_n_138__25_, r_n_138__24_, r_n_138__23_, r_n_138__22_, r_n_138__21_, r_n_138__20_, r_n_138__19_, r_n_138__18_, r_n_138__17_, r_n_138__16_, r_n_138__15_, r_n_138__14_, r_n_138__13_, r_n_138__12_, r_n_138__11_, r_n_138__10_, r_n_138__9_, r_n_138__8_, r_n_138__7_, r_n_138__6_, r_n_138__5_, r_n_138__4_, r_n_138__3_, r_n_138__2_, r_n_138__1_, r_n_138__0_ } = (N276)? { r_139__63_, r_139__62_, r_139__61_, r_139__60_, r_139__59_, r_139__58_, r_139__57_, r_139__56_, r_139__55_, r_139__54_, r_139__53_, r_139__52_, r_139__51_, r_139__50_, r_139__49_, r_139__48_, r_139__47_, r_139__46_, r_139__45_, r_139__44_, r_139__43_, r_139__42_, r_139__41_, r_139__40_, r_139__39_, r_139__38_, r_139__37_, r_139__36_, r_139__35_, r_139__34_, r_139__33_, r_139__32_, r_139__31_, r_139__30_, r_139__29_, r_139__28_, r_139__27_, r_139__26_, r_139__25_, r_139__24_, r_139__23_, r_139__22_, r_139__21_, r_139__20_, r_139__19_, r_139__18_, r_139__17_, r_139__16_, r_139__15_, r_139__14_, r_139__13_, r_139__12_, r_139__11_, r_139__10_, r_139__9_, r_139__8_, r_139__7_, r_139__6_, r_139__5_, r_139__4_, r_139__3_, r_139__2_, r_139__1_, r_139__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N277)? data_i : 1'b0;
  assign N276 = sel_i[276];
  assign N277 = N1718;
  assign { r_n_139__63_, r_n_139__62_, r_n_139__61_, r_n_139__60_, r_n_139__59_, r_n_139__58_, r_n_139__57_, r_n_139__56_, r_n_139__55_, r_n_139__54_, r_n_139__53_, r_n_139__52_, r_n_139__51_, r_n_139__50_, r_n_139__49_, r_n_139__48_, r_n_139__47_, r_n_139__46_, r_n_139__45_, r_n_139__44_, r_n_139__43_, r_n_139__42_, r_n_139__41_, r_n_139__40_, r_n_139__39_, r_n_139__38_, r_n_139__37_, r_n_139__36_, r_n_139__35_, r_n_139__34_, r_n_139__33_, r_n_139__32_, r_n_139__31_, r_n_139__30_, r_n_139__29_, r_n_139__28_, r_n_139__27_, r_n_139__26_, r_n_139__25_, r_n_139__24_, r_n_139__23_, r_n_139__22_, r_n_139__21_, r_n_139__20_, r_n_139__19_, r_n_139__18_, r_n_139__17_, r_n_139__16_, r_n_139__15_, r_n_139__14_, r_n_139__13_, r_n_139__12_, r_n_139__11_, r_n_139__10_, r_n_139__9_, r_n_139__8_, r_n_139__7_, r_n_139__6_, r_n_139__5_, r_n_139__4_, r_n_139__3_, r_n_139__2_, r_n_139__1_, r_n_139__0_ } = (N278)? { r_140__63_, r_140__62_, r_140__61_, r_140__60_, r_140__59_, r_140__58_, r_140__57_, r_140__56_, r_140__55_, r_140__54_, r_140__53_, r_140__52_, r_140__51_, r_140__50_, r_140__49_, r_140__48_, r_140__47_, r_140__46_, r_140__45_, r_140__44_, r_140__43_, r_140__42_, r_140__41_, r_140__40_, r_140__39_, r_140__38_, r_140__37_, r_140__36_, r_140__35_, r_140__34_, r_140__33_, r_140__32_, r_140__31_, r_140__30_, r_140__29_, r_140__28_, r_140__27_, r_140__26_, r_140__25_, r_140__24_, r_140__23_, r_140__22_, r_140__21_, r_140__20_, r_140__19_, r_140__18_, r_140__17_, r_140__16_, r_140__15_, r_140__14_, r_140__13_, r_140__12_, r_140__11_, r_140__10_, r_140__9_, r_140__8_, r_140__7_, r_140__6_, r_140__5_, r_140__4_, r_140__3_, r_140__2_, r_140__1_, r_140__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N279)? data_i : 1'b0;
  assign N278 = sel_i[278];
  assign N279 = N1723;
  assign { r_n_140__63_, r_n_140__62_, r_n_140__61_, r_n_140__60_, r_n_140__59_, r_n_140__58_, r_n_140__57_, r_n_140__56_, r_n_140__55_, r_n_140__54_, r_n_140__53_, r_n_140__52_, r_n_140__51_, r_n_140__50_, r_n_140__49_, r_n_140__48_, r_n_140__47_, r_n_140__46_, r_n_140__45_, r_n_140__44_, r_n_140__43_, r_n_140__42_, r_n_140__41_, r_n_140__40_, r_n_140__39_, r_n_140__38_, r_n_140__37_, r_n_140__36_, r_n_140__35_, r_n_140__34_, r_n_140__33_, r_n_140__32_, r_n_140__31_, r_n_140__30_, r_n_140__29_, r_n_140__28_, r_n_140__27_, r_n_140__26_, r_n_140__25_, r_n_140__24_, r_n_140__23_, r_n_140__22_, r_n_140__21_, r_n_140__20_, r_n_140__19_, r_n_140__18_, r_n_140__17_, r_n_140__16_, r_n_140__15_, r_n_140__14_, r_n_140__13_, r_n_140__12_, r_n_140__11_, r_n_140__10_, r_n_140__9_, r_n_140__8_, r_n_140__7_, r_n_140__6_, r_n_140__5_, r_n_140__4_, r_n_140__3_, r_n_140__2_, r_n_140__1_, r_n_140__0_ } = (N280)? { r_141__63_, r_141__62_, r_141__61_, r_141__60_, r_141__59_, r_141__58_, r_141__57_, r_141__56_, r_141__55_, r_141__54_, r_141__53_, r_141__52_, r_141__51_, r_141__50_, r_141__49_, r_141__48_, r_141__47_, r_141__46_, r_141__45_, r_141__44_, r_141__43_, r_141__42_, r_141__41_, r_141__40_, r_141__39_, r_141__38_, r_141__37_, r_141__36_, r_141__35_, r_141__34_, r_141__33_, r_141__32_, r_141__31_, r_141__30_, r_141__29_, r_141__28_, r_141__27_, r_141__26_, r_141__25_, r_141__24_, r_141__23_, r_141__22_, r_141__21_, r_141__20_, r_141__19_, r_141__18_, r_141__17_, r_141__16_, r_141__15_, r_141__14_, r_141__13_, r_141__12_, r_141__11_, r_141__10_, r_141__9_, r_141__8_, r_141__7_, r_141__6_, r_141__5_, r_141__4_, r_141__3_, r_141__2_, r_141__1_, r_141__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N281)? data_i : 1'b0;
  assign N280 = sel_i[280];
  assign N281 = N1728;
  assign { r_n_141__63_, r_n_141__62_, r_n_141__61_, r_n_141__60_, r_n_141__59_, r_n_141__58_, r_n_141__57_, r_n_141__56_, r_n_141__55_, r_n_141__54_, r_n_141__53_, r_n_141__52_, r_n_141__51_, r_n_141__50_, r_n_141__49_, r_n_141__48_, r_n_141__47_, r_n_141__46_, r_n_141__45_, r_n_141__44_, r_n_141__43_, r_n_141__42_, r_n_141__41_, r_n_141__40_, r_n_141__39_, r_n_141__38_, r_n_141__37_, r_n_141__36_, r_n_141__35_, r_n_141__34_, r_n_141__33_, r_n_141__32_, r_n_141__31_, r_n_141__30_, r_n_141__29_, r_n_141__28_, r_n_141__27_, r_n_141__26_, r_n_141__25_, r_n_141__24_, r_n_141__23_, r_n_141__22_, r_n_141__21_, r_n_141__20_, r_n_141__19_, r_n_141__18_, r_n_141__17_, r_n_141__16_, r_n_141__15_, r_n_141__14_, r_n_141__13_, r_n_141__12_, r_n_141__11_, r_n_141__10_, r_n_141__9_, r_n_141__8_, r_n_141__7_, r_n_141__6_, r_n_141__5_, r_n_141__4_, r_n_141__3_, r_n_141__2_, r_n_141__1_, r_n_141__0_ } = (N282)? { r_142__63_, r_142__62_, r_142__61_, r_142__60_, r_142__59_, r_142__58_, r_142__57_, r_142__56_, r_142__55_, r_142__54_, r_142__53_, r_142__52_, r_142__51_, r_142__50_, r_142__49_, r_142__48_, r_142__47_, r_142__46_, r_142__45_, r_142__44_, r_142__43_, r_142__42_, r_142__41_, r_142__40_, r_142__39_, r_142__38_, r_142__37_, r_142__36_, r_142__35_, r_142__34_, r_142__33_, r_142__32_, r_142__31_, r_142__30_, r_142__29_, r_142__28_, r_142__27_, r_142__26_, r_142__25_, r_142__24_, r_142__23_, r_142__22_, r_142__21_, r_142__20_, r_142__19_, r_142__18_, r_142__17_, r_142__16_, r_142__15_, r_142__14_, r_142__13_, r_142__12_, r_142__11_, r_142__10_, r_142__9_, r_142__8_, r_142__7_, r_142__6_, r_142__5_, r_142__4_, r_142__3_, r_142__2_, r_142__1_, r_142__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N283)? data_i : 1'b0;
  assign N282 = sel_i[282];
  assign N283 = N1733;
  assign { r_n_142__63_, r_n_142__62_, r_n_142__61_, r_n_142__60_, r_n_142__59_, r_n_142__58_, r_n_142__57_, r_n_142__56_, r_n_142__55_, r_n_142__54_, r_n_142__53_, r_n_142__52_, r_n_142__51_, r_n_142__50_, r_n_142__49_, r_n_142__48_, r_n_142__47_, r_n_142__46_, r_n_142__45_, r_n_142__44_, r_n_142__43_, r_n_142__42_, r_n_142__41_, r_n_142__40_, r_n_142__39_, r_n_142__38_, r_n_142__37_, r_n_142__36_, r_n_142__35_, r_n_142__34_, r_n_142__33_, r_n_142__32_, r_n_142__31_, r_n_142__30_, r_n_142__29_, r_n_142__28_, r_n_142__27_, r_n_142__26_, r_n_142__25_, r_n_142__24_, r_n_142__23_, r_n_142__22_, r_n_142__21_, r_n_142__20_, r_n_142__19_, r_n_142__18_, r_n_142__17_, r_n_142__16_, r_n_142__15_, r_n_142__14_, r_n_142__13_, r_n_142__12_, r_n_142__11_, r_n_142__10_, r_n_142__9_, r_n_142__8_, r_n_142__7_, r_n_142__6_, r_n_142__5_, r_n_142__4_, r_n_142__3_, r_n_142__2_, r_n_142__1_, r_n_142__0_ } = (N284)? { r_143__63_, r_143__62_, r_143__61_, r_143__60_, r_143__59_, r_143__58_, r_143__57_, r_143__56_, r_143__55_, r_143__54_, r_143__53_, r_143__52_, r_143__51_, r_143__50_, r_143__49_, r_143__48_, r_143__47_, r_143__46_, r_143__45_, r_143__44_, r_143__43_, r_143__42_, r_143__41_, r_143__40_, r_143__39_, r_143__38_, r_143__37_, r_143__36_, r_143__35_, r_143__34_, r_143__33_, r_143__32_, r_143__31_, r_143__30_, r_143__29_, r_143__28_, r_143__27_, r_143__26_, r_143__25_, r_143__24_, r_143__23_, r_143__22_, r_143__21_, r_143__20_, r_143__19_, r_143__18_, r_143__17_, r_143__16_, r_143__15_, r_143__14_, r_143__13_, r_143__12_, r_143__11_, r_143__10_, r_143__9_, r_143__8_, r_143__7_, r_143__6_, r_143__5_, r_143__4_, r_143__3_, r_143__2_, r_143__1_, r_143__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N285)? data_i : 1'b0;
  assign N284 = sel_i[284];
  assign N285 = N1738;
  assign { r_n_143__63_, r_n_143__62_, r_n_143__61_, r_n_143__60_, r_n_143__59_, r_n_143__58_, r_n_143__57_, r_n_143__56_, r_n_143__55_, r_n_143__54_, r_n_143__53_, r_n_143__52_, r_n_143__51_, r_n_143__50_, r_n_143__49_, r_n_143__48_, r_n_143__47_, r_n_143__46_, r_n_143__45_, r_n_143__44_, r_n_143__43_, r_n_143__42_, r_n_143__41_, r_n_143__40_, r_n_143__39_, r_n_143__38_, r_n_143__37_, r_n_143__36_, r_n_143__35_, r_n_143__34_, r_n_143__33_, r_n_143__32_, r_n_143__31_, r_n_143__30_, r_n_143__29_, r_n_143__28_, r_n_143__27_, r_n_143__26_, r_n_143__25_, r_n_143__24_, r_n_143__23_, r_n_143__22_, r_n_143__21_, r_n_143__20_, r_n_143__19_, r_n_143__18_, r_n_143__17_, r_n_143__16_, r_n_143__15_, r_n_143__14_, r_n_143__13_, r_n_143__12_, r_n_143__11_, r_n_143__10_, r_n_143__9_, r_n_143__8_, r_n_143__7_, r_n_143__6_, r_n_143__5_, r_n_143__4_, r_n_143__3_, r_n_143__2_, r_n_143__1_, r_n_143__0_ } = (N286)? { r_144__63_, r_144__62_, r_144__61_, r_144__60_, r_144__59_, r_144__58_, r_144__57_, r_144__56_, r_144__55_, r_144__54_, r_144__53_, r_144__52_, r_144__51_, r_144__50_, r_144__49_, r_144__48_, r_144__47_, r_144__46_, r_144__45_, r_144__44_, r_144__43_, r_144__42_, r_144__41_, r_144__40_, r_144__39_, r_144__38_, r_144__37_, r_144__36_, r_144__35_, r_144__34_, r_144__33_, r_144__32_, r_144__31_, r_144__30_, r_144__29_, r_144__28_, r_144__27_, r_144__26_, r_144__25_, r_144__24_, r_144__23_, r_144__22_, r_144__21_, r_144__20_, r_144__19_, r_144__18_, r_144__17_, r_144__16_, r_144__15_, r_144__14_, r_144__13_, r_144__12_, r_144__11_, r_144__10_, r_144__9_, r_144__8_, r_144__7_, r_144__6_, r_144__5_, r_144__4_, r_144__3_, r_144__2_, r_144__1_, r_144__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N287)? data_i : 1'b0;
  assign N286 = sel_i[286];
  assign N287 = N1743;
  assign { r_n_144__63_, r_n_144__62_, r_n_144__61_, r_n_144__60_, r_n_144__59_, r_n_144__58_, r_n_144__57_, r_n_144__56_, r_n_144__55_, r_n_144__54_, r_n_144__53_, r_n_144__52_, r_n_144__51_, r_n_144__50_, r_n_144__49_, r_n_144__48_, r_n_144__47_, r_n_144__46_, r_n_144__45_, r_n_144__44_, r_n_144__43_, r_n_144__42_, r_n_144__41_, r_n_144__40_, r_n_144__39_, r_n_144__38_, r_n_144__37_, r_n_144__36_, r_n_144__35_, r_n_144__34_, r_n_144__33_, r_n_144__32_, r_n_144__31_, r_n_144__30_, r_n_144__29_, r_n_144__28_, r_n_144__27_, r_n_144__26_, r_n_144__25_, r_n_144__24_, r_n_144__23_, r_n_144__22_, r_n_144__21_, r_n_144__20_, r_n_144__19_, r_n_144__18_, r_n_144__17_, r_n_144__16_, r_n_144__15_, r_n_144__14_, r_n_144__13_, r_n_144__12_, r_n_144__11_, r_n_144__10_, r_n_144__9_, r_n_144__8_, r_n_144__7_, r_n_144__6_, r_n_144__5_, r_n_144__4_, r_n_144__3_, r_n_144__2_, r_n_144__1_, r_n_144__0_ } = (N288)? { r_145__63_, r_145__62_, r_145__61_, r_145__60_, r_145__59_, r_145__58_, r_145__57_, r_145__56_, r_145__55_, r_145__54_, r_145__53_, r_145__52_, r_145__51_, r_145__50_, r_145__49_, r_145__48_, r_145__47_, r_145__46_, r_145__45_, r_145__44_, r_145__43_, r_145__42_, r_145__41_, r_145__40_, r_145__39_, r_145__38_, r_145__37_, r_145__36_, r_145__35_, r_145__34_, r_145__33_, r_145__32_, r_145__31_, r_145__30_, r_145__29_, r_145__28_, r_145__27_, r_145__26_, r_145__25_, r_145__24_, r_145__23_, r_145__22_, r_145__21_, r_145__20_, r_145__19_, r_145__18_, r_145__17_, r_145__16_, r_145__15_, r_145__14_, r_145__13_, r_145__12_, r_145__11_, r_145__10_, r_145__9_, r_145__8_, r_145__7_, r_145__6_, r_145__5_, r_145__4_, r_145__3_, r_145__2_, r_145__1_, r_145__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N289)? data_i : 1'b0;
  assign N288 = sel_i[288];
  assign N289 = N1748;
  assign { r_n_145__63_, r_n_145__62_, r_n_145__61_, r_n_145__60_, r_n_145__59_, r_n_145__58_, r_n_145__57_, r_n_145__56_, r_n_145__55_, r_n_145__54_, r_n_145__53_, r_n_145__52_, r_n_145__51_, r_n_145__50_, r_n_145__49_, r_n_145__48_, r_n_145__47_, r_n_145__46_, r_n_145__45_, r_n_145__44_, r_n_145__43_, r_n_145__42_, r_n_145__41_, r_n_145__40_, r_n_145__39_, r_n_145__38_, r_n_145__37_, r_n_145__36_, r_n_145__35_, r_n_145__34_, r_n_145__33_, r_n_145__32_, r_n_145__31_, r_n_145__30_, r_n_145__29_, r_n_145__28_, r_n_145__27_, r_n_145__26_, r_n_145__25_, r_n_145__24_, r_n_145__23_, r_n_145__22_, r_n_145__21_, r_n_145__20_, r_n_145__19_, r_n_145__18_, r_n_145__17_, r_n_145__16_, r_n_145__15_, r_n_145__14_, r_n_145__13_, r_n_145__12_, r_n_145__11_, r_n_145__10_, r_n_145__9_, r_n_145__8_, r_n_145__7_, r_n_145__6_, r_n_145__5_, r_n_145__4_, r_n_145__3_, r_n_145__2_, r_n_145__1_, r_n_145__0_ } = (N290)? { r_146__63_, r_146__62_, r_146__61_, r_146__60_, r_146__59_, r_146__58_, r_146__57_, r_146__56_, r_146__55_, r_146__54_, r_146__53_, r_146__52_, r_146__51_, r_146__50_, r_146__49_, r_146__48_, r_146__47_, r_146__46_, r_146__45_, r_146__44_, r_146__43_, r_146__42_, r_146__41_, r_146__40_, r_146__39_, r_146__38_, r_146__37_, r_146__36_, r_146__35_, r_146__34_, r_146__33_, r_146__32_, r_146__31_, r_146__30_, r_146__29_, r_146__28_, r_146__27_, r_146__26_, r_146__25_, r_146__24_, r_146__23_, r_146__22_, r_146__21_, r_146__20_, r_146__19_, r_146__18_, r_146__17_, r_146__16_, r_146__15_, r_146__14_, r_146__13_, r_146__12_, r_146__11_, r_146__10_, r_146__9_, r_146__8_, r_146__7_, r_146__6_, r_146__5_, r_146__4_, r_146__3_, r_146__2_, r_146__1_, r_146__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N291)? data_i : 1'b0;
  assign N290 = sel_i[290];
  assign N291 = N1753;
  assign { r_n_146__63_, r_n_146__62_, r_n_146__61_, r_n_146__60_, r_n_146__59_, r_n_146__58_, r_n_146__57_, r_n_146__56_, r_n_146__55_, r_n_146__54_, r_n_146__53_, r_n_146__52_, r_n_146__51_, r_n_146__50_, r_n_146__49_, r_n_146__48_, r_n_146__47_, r_n_146__46_, r_n_146__45_, r_n_146__44_, r_n_146__43_, r_n_146__42_, r_n_146__41_, r_n_146__40_, r_n_146__39_, r_n_146__38_, r_n_146__37_, r_n_146__36_, r_n_146__35_, r_n_146__34_, r_n_146__33_, r_n_146__32_, r_n_146__31_, r_n_146__30_, r_n_146__29_, r_n_146__28_, r_n_146__27_, r_n_146__26_, r_n_146__25_, r_n_146__24_, r_n_146__23_, r_n_146__22_, r_n_146__21_, r_n_146__20_, r_n_146__19_, r_n_146__18_, r_n_146__17_, r_n_146__16_, r_n_146__15_, r_n_146__14_, r_n_146__13_, r_n_146__12_, r_n_146__11_, r_n_146__10_, r_n_146__9_, r_n_146__8_, r_n_146__7_, r_n_146__6_, r_n_146__5_, r_n_146__4_, r_n_146__3_, r_n_146__2_, r_n_146__1_, r_n_146__0_ } = (N292)? { r_147__63_, r_147__62_, r_147__61_, r_147__60_, r_147__59_, r_147__58_, r_147__57_, r_147__56_, r_147__55_, r_147__54_, r_147__53_, r_147__52_, r_147__51_, r_147__50_, r_147__49_, r_147__48_, r_147__47_, r_147__46_, r_147__45_, r_147__44_, r_147__43_, r_147__42_, r_147__41_, r_147__40_, r_147__39_, r_147__38_, r_147__37_, r_147__36_, r_147__35_, r_147__34_, r_147__33_, r_147__32_, r_147__31_, r_147__30_, r_147__29_, r_147__28_, r_147__27_, r_147__26_, r_147__25_, r_147__24_, r_147__23_, r_147__22_, r_147__21_, r_147__20_, r_147__19_, r_147__18_, r_147__17_, r_147__16_, r_147__15_, r_147__14_, r_147__13_, r_147__12_, r_147__11_, r_147__10_, r_147__9_, r_147__8_, r_147__7_, r_147__6_, r_147__5_, r_147__4_, r_147__3_, r_147__2_, r_147__1_, r_147__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N293)? data_i : 1'b0;
  assign N292 = sel_i[292];
  assign N293 = N1758;
  assign { r_n_147__63_, r_n_147__62_, r_n_147__61_, r_n_147__60_, r_n_147__59_, r_n_147__58_, r_n_147__57_, r_n_147__56_, r_n_147__55_, r_n_147__54_, r_n_147__53_, r_n_147__52_, r_n_147__51_, r_n_147__50_, r_n_147__49_, r_n_147__48_, r_n_147__47_, r_n_147__46_, r_n_147__45_, r_n_147__44_, r_n_147__43_, r_n_147__42_, r_n_147__41_, r_n_147__40_, r_n_147__39_, r_n_147__38_, r_n_147__37_, r_n_147__36_, r_n_147__35_, r_n_147__34_, r_n_147__33_, r_n_147__32_, r_n_147__31_, r_n_147__30_, r_n_147__29_, r_n_147__28_, r_n_147__27_, r_n_147__26_, r_n_147__25_, r_n_147__24_, r_n_147__23_, r_n_147__22_, r_n_147__21_, r_n_147__20_, r_n_147__19_, r_n_147__18_, r_n_147__17_, r_n_147__16_, r_n_147__15_, r_n_147__14_, r_n_147__13_, r_n_147__12_, r_n_147__11_, r_n_147__10_, r_n_147__9_, r_n_147__8_, r_n_147__7_, r_n_147__6_, r_n_147__5_, r_n_147__4_, r_n_147__3_, r_n_147__2_, r_n_147__1_, r_n_147__0_ } = (N294)? { r_148__63_, r_148__62_, r_148__61_, r_148__60_, r_148__59_, r_148__58_, r_148__57_, r_148__56_, r_148__55_, r_148__54_, r_148__53_, r_148__52_, r_148__51_, r_148__50_, r_148__49_, r_148__48_, r_148__47_, r_148__46_, r_148__45_, r_148__44_, r_148__43_, r_148__42_, r_148__41_, r_148__40_, r_148__39_, r_148__38_, r_148__37_, r_148__36_, r_148__35_, r_148__34_, r_148__33_, r_148__32_, r_148__31_, r_148__30_, r_148__29_, r_148__28_, r_148__27_, r_148__26_, r_148__25_, r_148__24_, r_148__23_, r_148__22_, r_148__21_, r_148__20_, r_148__19_, r_148__18_, r_148__17_, r_148__16_, r_148__15_, r_148__14_, r_148__13_, r_148__12_, r_148__11_, r_148__10_, r_148__9_, r_148__8_, r_148__7_, r_148__6_, r_148__5_, r_148__4_, r_148__3_, r_148__2_, r_148__1_, r_148__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N295)? data_i : 1'b0;
  assign N294 = sel_i[294];
  assign N295 = N1763;
  assign { r_n_148__63_, r_n_148__62_, r_n_148__61_, r_n_148__60_, r_n_148__59_, r_n_148__58_, r_n_148__57_, r_n_148__56_, r_n_148__55_, r_n_148__54_, r_n_148__53_, r_n_148__52_, r_n_148__51_, r_n_148__50_, r_n_148__49_, r_n_148__48_, r_n_148__47_, r_n_148__46_, r_n_148__45_, r_n_148__44_, r_n_148__43_, r_n_148__42_, r_n_148__41_, r_n_148__40_, r_n_148__39_, r_n_148__38_, r_n_148__37_, r_n_148__36_, r_n_148__35_, r_n_148__34_, r_n_148__33_, r_n_148__32_, r_n_148__31_, r_n_148__30_, r_n_148__29_, r_n_148__28_, r_n_148__27_, r_n_148__26_, r_n_148__25_, r_n_148__24_, r_n_148__23_, r_n_148__22_, r_n_148__21_, r_n_148__20_, r_n_148__19_, r_n_148__18_, r_n_148__17_, r_n_148__16_, r_n_148__15_, r_n_148__14_, r_n_148__13_, r_n_148__12_, r_n_148__11_, r_n_148__10_, r_n_148__9_, r_n_148__8_, r_n_148__7_, r_n_148__6_, r_n_148__5_, r_n_148__4_, r_n_148__3_, r_n_148__2_, r_n_148__1_, r_n_148__0_ } = (N296)? { r_149__63_, r_149__62_, r_149__61_, r_149__60_, r_149__59_, r_149__58_, r_149__57_, r_149__56_, r_149__55_, r_149__54_, r_149__53_, r_149__52_, r_149__51_, r_149__50_, r_149__49_, r_149__48_, r_149__47_, r_149__46_, r_149__45_, r_149__44_, r_149__43_, r_149__42_, r_149__41_, r_149__40_, r_149__39_, r_149__38_, r_149__37_, r_149__36_, r_149__35_, r_149__34_, r_149__33_, r_149__32_, r_149__31_, r_149__30_, r_149__29_, r_149__28_, r_149__27_, r_149__26_, r_149__25_, r_149__24_, r_149__23_, r_149__22_, r_149__21_, r_149__20_, r_149__19_, r_149__18_, r_149__17_, r_149__16_, r_149__15_, r_149__14_, r_149__13_, r_149__12_, r_149__11_, r_149__10_, r_149__9_, r_149__8_, r_149__7_, r_149__6_, r_149__5_, r_149__4_, r_149__3_, r_149__2_, r_149__1_, r_149__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N297)? data_i : 1'b0;
  assign N296 = sel_i[296];
  assign N297 = N1768;
  assign { r_n_149__63_, r_n_149__62_, r_n_149__61_, r_n_149__60_, r_n_149__59_, r_n_149__58_, r_n_149__57_, r_n_149__56_, r_n_149__55_, r_n_149__54_, r_n_149__53_, r_n_149__52_, r_n_149__51_, r_n_149__50_, r_n_149__49_, r_n_149__48_, r_n_149__47_, r_n_149__46_, r_n_149__45_, r_n_149__44_, r_n_149__43_, r_n_149__42_, r_n_149__41_, r_n_149__40_, r_n_149__39_, r_n_149__38_, r_n_149__37_, r_n_149__36_, r_n_149__35_, r_n_149__34_, r_n_149__33_, r_n_149__32_, r_n_149__31_, r_n_149__30_, r_n_149__29_, r_n_149__28_, r_n_149__27_, r_n_149__26_, r_n_149__25_, r_n_149__24_, r_n_149__23_, r_n_149__22_, r_n_149__21_, r_n_149__20_, r_n_149__19_, r_n_149__18_, r_n_149__17_, r_n_149__16_, r_n_149__15_, r_n_149__14_, r_n_149__13_, r_n_149__12_, r_n_149__11_, r_n_149__10_, r_n_149__9_, r_n_149__8_, r_n_149__7_, r_n_149__6_, r_n_149__5_, r_n_149__4_, r_n_149__3_, r_n_149__2_, r_n_149__1_, r_n_149__0_ } = (N298)? { r_150__63_, r_150__62_, r_150__61_, r_150__60_, r_150__59_, r_150__58_, r_150__57_, r_150__56_, r_150__55_, r_150__54_, r_150__53_, r_150__52_, r_150__51_, r_150__50_, r_150__49_, r_150__48_, r_150__47_, r_150__46_, r_150__45_, r_150__44_, r_150__43_, r_150__42_, r_150__41_, r_150__40_, r_150__39_, r_150__38_, r_150__37_, r_150__36_, r_150__35_, r_150__34_, r_150__33_, r_150__32_, r_150__31_, r_150__30_, r_150__29_, r_150__28_, r_150__27_, r_150__26_, r_150__25_, r_150__24_, r_150__23_, r_150__22_, r_150__21_, r_150__20_, r_150__19_, r_150__18_, r_150__17_, r_150__16_, r_150__15_, r_150__14_, r_150__13_, r_150__12_, r_150__11_, r_150__10_, r_150__9_, r_150__8_, r_150__7_, r_150__6_, r_150__5_, r_150__4_, r_150__3_, r_150__2_, r_150__1_, r_150__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N299)? data_i : 1'b0;
  assign N298 = sel_i[298];
  assign N299 = N1773;
  assign { r_n_150__63_, r_n_150__62_, r_n_150__61_, r_n_150__60_, r_n_150__59_, r_n_150__58_, r_n_150__57_, r_n_150__56_, r_n_150__55_, r_n_150__54_, r_n_150__53_, r_n_150__52_, r_n_150__51_, r_n_150__50_, r_n_150__49_, r_n_150__48_, r_n_150__47_, r_n_150__46_, r_n_150__45_, r_n_150__44_, r_n_150__43_, r_n_150__42_, r_n_150__41_, r_n_150__40_, r_n_150__39_, r_n_150__38_, r_n_150__37_, r_n_150__36_, r_n_150__35_, r_n_150__34_, r_n_150__33_, r_n_150__32_, r_n_150__31_, r_n_150__30_, r_n_150__29_, r_n_150__28_, r_n_150__27_, r_n_150__26_, r_n_150__25_, r_n_150__24_, r_n_150__23_, r_n_150__22_, r_n_150__21_, r_n_150__20_, r_n_150__19_, r_n_150__18_, r_n_150__17_, r_n_150__16_, r_n_150__15_, r_n_150__14_, r_n_150__13_, r_n_150__12_, r_n_150__11_, r_n_150__10_, r_n_150__9_, r_n_150__8_, r_n_150__7_, r_n_150__6_, r_n_150__5_, r_n_150__4_, r_n_150__3_, r_n_150__2_, r_n_150__1_, r_n_150__0_ } = (N300)? { r_151__63_, r_151__62_, r_151__61_, r_151__60_, r_151__59_, r_151__58_, r_151__57_, r_151__56_, r_151__55_, r_151__54_, r_151__53_, r_151__52_, r_151__51_, r_151__50_, r_151__49_, r_151__48_, r_151__47_, r_151__46_, r_151__45_, r_151__44_, r_151__43_, r_151__42_, r_151__41_, r_151__40_, r_151__39_, r_151__38_, r_151__37_, r_151__36_, r_151__35_, r_151__34_, r_151__33_, r_151__32_, r_151__31_, r_151__30_, r_151__29_, r_151__28_, r_151__27_, r_151__26_, r_151__25_, r_151__24_, r_151__23_, r_151__22_, r_151__21_, r_151__20_, r_151__19_, r_151__18_, r_151__17_, r_151__16_, r_151__15_, r_151__14_, r_151__13_, r_151__12_, r_151__11_, r_151__10_, r_151__9_, r_151__8_, r_151__7_, r_151__6_, r_151__5_, r_151__4_, r_151__3_, r_151__2_, r_151__1_, r_151__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N301)? data_i : 1'b0;
  assign N300 = sel_i[300];
  assign N301 = N1778;
  assign { r_n_151__63_, r_n_151__62_, r_n_151__61_, r_n_151__60_, r_n_151__59_, r_n_151__58_, r_n_151__57_, r_n_151__56_, r_n_151__55_, r_n_151__54_, r_n_151__53_, r_n_151__52_, r_n_151__51_, r_n_151__50_, r_n_151__49_, r_n_151__48_, r_n_151__47_, r_n_151__46_, r_n_151__45_, r_n_151__44_, r_n_151__43_, r_n_151__42_, r_n_151__41_, r_n_151__40_, r_n_151__39_, r_n_151__38_, r_n_151__37_, r_n_151__36_, r_n_151__35_, r_n_151__34_, r_n_151__33_, r_n_151__32_, r_n_151__31_, r_n_151__30_, r_n_151__29_, r_n_151__28_, r_n_151__27_, r_n_151__26_, r_n_151__25_, r_n_151__24_, r_n_151__23_, r_n_151__22_, r_n_151__21_, r_n_151__20_, r_n_151__19_, r_n_151__18_, r_n_151__17_, r_n_151__16_, r_n_151__15_, r_n_151__14_, r_n_151__13_, r_n_151__12_, r_n_151__11_, r_n_151__10_, r_n_151__9_, r_n_151__8_, r_n_151__7_, r_n_151__6_, r_n_151__5_, r_n_151__4_, r_n_151__3_, r_n_151__2_, r_n_151__1_, r_n_151__0_ } = (N302)? { r_152__63_, r_152__62_, r_152__61_, r_152__60_, r_152__59_, r_152__58_, r_152__57_, r_152__56_, r_152__55_, r_152__54_, r_152__53_, r_152__52_, r_152__51_, r_152__50_, r_152__49_, r_152__48_, r_152__47_, r_152__46_, r_152__45_, r_152__44_, r_152__43_, r_152__42_, r_152__41_, r_152__40_, r_152__39_, r_152__38_, r_152__37_, r_152__36_, r_152__35_, r_152__34_, r_152__33_, r_152__32_, r_152__31_, r_152__30_, r_152__29_, r_152__28_, r_152__27_, r_152__26_, r_152__25_, r_152__24_, r_152__23_, r_152__22_, r_152__21_, r_152__20_, r_152__19_, r_152__18_, r_152__17_, r_152__16_, r_152__15_, r_152__14_, r_152__13_, r_152__12_, r_152__11_, r_152__10_, r_152__9_, r_152__8_, r_152__7_, r_152__6_, r_152__5_, r_152__4_, r_152__3_, r_152__2_, r_152__1_, r_152__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N303)? data_i : 1'b0;
  assign N302 = sel_i[302];
  assign N303 = N1783;
  assign { r_n_152__63_, r_n_152__62_, r_n_152__61_, r_n_152__60_, r_n_152__59_, r_n_152__58_, r_n_152__57_, r_n_152__56_, r_n_152__55_, r_n_152__54_, r_n_152__53_, r_n_152__52_, r_n_152__51_, r_n_152__50_, r_n_152__49_, r_n_152__48_, r_n_152__47_, r_n_152__46_, r_n_152__45_, r_n_152__44_, r_n_152__43_, r_n_152__42_, r_n_152__41_, r_n_152__40_, r_n_152__39_, r_n_152__38_, r_n_152__37_, r_n_152__36_, r_n_152__35_, r_n_152__34_, r_n_152__33_, r_n_152__32_, r_n_152__31_, r_n_152__30_, r_n_152__29_, r_n_152__28_, r_n_152__27_, r_n_152__26_, r_n_152__25_, r_n_152__24_, r_n_152__23_, r_n_152__22_, r_n_152__21_, r_n_152__20_, r_n_152__19_, r_n_152__18_, r_n_152__17_, r_n_152__16_, r_n_152__15_, r_n_152__14_, r_n_152__13_, r_n_152__12_, r_n_152__11_, r_n_152__10_, r_n_152__9_, r_n_152__8_, r_n_152__7_, r_n_152__6_, r_n_152__5_, r_n_152__4_, r_n_152__3_, r_n_152__2_, r_n_152__1_, r_n_152__0_ } = (N304)? { r_153__63_, r_153__62_, r_153__61_, r_153__60_, r_153__59_, r_153__58_, r_153__57_, r_153__56_, r_153__55_, r_153__54_, r_153__53_, r_153__52_, r_153__51_, r_153__50_, r_153__49_, r_153__48_, r_153__47_, r_153__46_, r_153__45_, r_153__44_, r_153__43_, r_153__42_, r_153__41_, r_153__40_, r_153__39_, r_153__38_, r_153__37_, r_153__36_, r_153__35_, r_153__34_, r_153__33_, r_153__32_, r_153__31_, r_153__30_, r_153__29_, r_153__28_, r_153__27_, r_153__26_, r_153__25_, r_153__24_, r_153__23_, r_153__22_, r_153__21_, r_153__20_, r_153__19_, r_153__18_, r_153__17_, r_153__16_, r_153__15_, r_153__14_, r_153__13_, r_153__12_, r_153__11_, r_153__10_, r_153__9_, r_153__8_, r_153__7_, r_153__6_, r_153__5_, r_153__4_, r_153__3_, r_153__2_, r_153__1_, r_153__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N305)? data_i : 1'b0;
  assign N304 = sel_i[304];
  assign N305 = N1788;
  assign { r_n_153__63_, r_n_153__62_, r_n_153__61_, r_n_153__60_, r_n_153__59_, r_n_153__58_, r_n_153__57_, r_n_153__56_, r_n_153__55_, r_n_153__54_, r_n_153__53_, r_n_153__52_, r_n_153__51_, r_n_153__50_, r_n_153__49_, r_n_153__48_, r_n_153__47_, r_n_153__46_, r_n_153__45_, r_n_153__44_, r_n_153__43_, r_n_153__42_, r_n_153__41_, r_n_153__40_, r_n_153__39_, r_n_153__38_, r_n_153__37_, r_n_153__36_, r_n_153__35_, r_n_153__34_, r_n_153__33_, r_n_153__32_, r_n_153__31_, r_n_153__30_, r_n_153__29_, r_n_153__28_, r_n_153__27_, r_n_153__26_, r_n_153__25_, r_n_153__24_, r_n_153__23_, r_n_153__22_, r_n_153__21_, r_n_153__20_, r_n_153__19_, r_n_153__18_, r_n_153__17_, r_n_153__16_, r_n_153__15_, r_n_153__14_, r_n_153__13_, r_n_153__12_, r_n_153__11_, r_n_153__10_, r_n_153__9_, r_n_153__8_, r_n_153__7_, r_n_153__6_, r_n_153__5_, r_n_153__4_, r_n_153__3_, r_n_153__2_, r_n_153__1_, r_n_153__0_ } = (N306)? { r_154__63_, r_154__62_, r_154__61_, r_154__60_, r_154__59_, r_154__58_, r_154__57_, r_154__56_, r_154__55_, r_154__54_, r_154__53_, r_154__52_, r_154__51_, r_154__50_, r_154__49_, r_154__48_, r_154__47_, r_154__46_, r_154__45_, r_154__44_, r_154__43_, r_154__42_, r_154__41_, r_154__40_, r_154__39_, r_154__38_, r_154__37_, r_154__36_, r_154__35_, r_154__34_, r_154__33_, r_154__32_, r_154__31_, r_154__30_, r_154__29_, r_154__28_, r_154__27_, r_154__26_, r_154__25_, r_154__24_, r_154__23_, r_154__22_, r_154__21_, r_154__20_, r_154__19_, r_154__18_, r_154__17_, r_154__16_, r_154__15_, r_154__14_, r_154__13_, r_154__12_, r_154__11_, r_154__10_, r_154__9_, r_154__8_, r_154__7_, r_154__6_, r_154__5_, r_154__4_, r_154__3_, r_154__2_, r_154__1_, r_154__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N307)? data_i : 1'b0;
  assign N306 = sel_i[306];
  assign N307 = N1793;
  assign { r_n_154__63_, r_n_154__62_, r_n_154__61_, r_n_154__60_, r_n_154__59_, r_n_154__58_, r_n_154__57_, r_n_154__56_, r_n_154__55_, r_n_154__54_, r_n_154__53_, r_n_154__52_, r_n_154__51_, r_n_154__50_, r_n_154__49_, r_n_154__48_, r_n_154__47_, r_n_154__46_, r_n_154__45_, r_n_154__44_, r_n_154__43_, r_n_154__42_, r_n_154__41_, r_n_154__40_, r_n_154__39_, r_n_154__38_, r_n_154__37_, r_n_154__36_, r_n_154__35_, r_n_154__34_, r_n_154__33_, r_n_154__32_, r_n_154__31_, r_n_154__30_, r_n_154__29_, r_n_154__28_, r_n_154__27_, r_n_154__26_, r_n_154__25_, r_n_154__24_, r_n_154__23_, r_n_154__22_, r_n_154__21_, r_n_154__20_, r_n_154__19_, r_n_154__18_, r_n_154__17_, r_n_154__16_, r_n_154__15_, r_n_154__14_, r_n_154__13_, r_n_154__12_, r_n_154__11_, r_n_154__10_, r_n_154__9_, r_n_154__8_, r_n_154__7_, r_n_154__6_, r_n_154__5_, r_n_154__4_, r_n_154__3_, r_n_154__2_, r_n_154__1_, r_n_154__0_ } = (N308)? { r_155__63_, r_155__62_, r_155__61_, r_155__60_, r_155__59_, r_155__58_, r_155__57_, r_155__56_, r_155__55_, r_155__54_, r_155__53_, r_155__52_, r_155__51_, r_155__50_, r_155__49_, r_155__48_, r_155__47_, r_155__46_, r_155__45_, r_155__44_, r_155__43_, r_155__42_, r_155__41_, r_155__40_, r_155__39_, r_155__38_, r_155__37_, r_155__36_, r_155__35_, r_155__34_, r_155__33_, r_155__32_, r_155__31_, r_155__30_, r_155__29_, r_155__28_, r_155__27_, r_155__26_, r_155__25_, r_155__24_, r_155__23_, r_155__22_, r_155__21_, r_155__20_, r_155__19_, r_155__18_, r_155__17_, r_155__16_, r_155__15_, r_155__14_, r_155__13_, r_155__12_, r_155__11_, r_155__10_, r_155__9_, r_155__8_, r_155__7_, r_155__6_, r_155__5_, r_155__4_, r_155__3_, r_155__2_, r_155__1_, r_155__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N309)? data_i : 1'b0;
  assign N308 = sel_i[308];
  assign N309 = N1798;
  assign { r_n_155__63_, r_n_155__62_, r_n_155__61_, r_n_155__60_, r_n_155__59_, r_n_155__58_, r_n_155__57_, r_n_155__56_, r_n_155__55_, r_n_155__54_, r_n_155__53_, r_n_155__52_, r_n_155__51_, r_n_155__50_, r_n_155__49_, r_n_155__48_, r_n_155__47_, r_n_155__46_, r_n_155__45_, r_n_155__44_, r_n_155__43_, r_n_155__42_, r_n_155__41_, r_n_155__40_, r_n_155__39_, r_n_155__38_, r_n_155__37_, r_n_155__36_, r_n_155__35_, r_n_155__34_, r_n_155__33_, r_n_155__32_, r_n_155__31_, r_n_155__30_, r_n_155__29_, r_n_155__28_, r_n_155__27_, r_n_155__26_, r_n_155__25_, r_n_155__24_, r_n_155__23_, r_n_155__22_, r_n_155__21_, r_n_155__20_, r_n_155__19_, r_n_155__18_, r_n_155__17_, r_n_155__16_, r_n_155__15_, r_n_155__14_, r_n_155__13_, r_n_155__12_, r_n_155__11_, r_n_155__10_, r_n_155__9_, r_n_155__8_, r_n_155__7_, r_n_155__6_, r_n_155__5_, r_n_155__4_, r_n_155__3_, r_n_155__2_, r_n_155__1_, r_n_155__0_ } = (N310)? { r_156__63_, r_156__62_, r_156__61_, r_156__60_, r_156__59_, r_156__58_, r_156__57_, r_156__56_, r_156__55_, r_156__54_, r_156__53_, r_156__52_, r_156__51_, r_156__50_, r_156__49_, r_156__48_, r_156__47_, r_156__46_, r_156__45_, r_156__44_, r_156__43_, r_156__42_, r_156__41_, r_156__40_, r_156__39_, r_156__38_, r_156__37_, r_156__36_, r_156__35_, r_156__34_, r_156__33_, r_156__32_, r_156__31_, r_156__30_, r_156__29_, r_156__28_, r_156__27_, r_156__26_, r_156__25_, r_156__24_, r_156__23_, r_156__22_, r_156__21_, r_156__20_, r_156__19_, r_156__18_, r_156__17_, r_156__16_, r_156__15_, r_156__14_, r_156__13_, r_156__12_, r_156__11_, r_156__10_, r_156__9_, r_156__8_, r_156__7_, r_156__6_, r_156__5_, r_156__4_, r_156__3_, r_156__2_, r_156__1_, r_156__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N311)? data_i : 1'b0;
  assign N310 = sel_i[310];
  assign N311 = N1803;
  assign { r_n_156__63_, r_n_156__62_, r_n_156__61_, r_n_156__60_, r_n_156__59_, r_n_156__58_, r_n_156__57_, r_n_156__56_, r_n_156__55_, r_n_156__54_, r_n_156__53_, r_n_156__52_, r_n_156__51_, r_n_156__50_, r_n_156__49_, r_n_156__48_, r_n_156__47_, r_n_156__46_, r_n_156__45_, r_n_156__44_, r_n_156__43_, r_n_156__42_, r_n_156__41_, r_n_156__40_, r_n_156__39_, r_n_156__38_, r_n_156__37_, r_n_156__36_, r_n_156__35_, r_n_156__34_, r_n_156__33_, r_n_156__32_, r_n_156__31_, r_n_156__30_, r_n_156__29_, r_n_156__28_, r_n_156__27_, r_n_156__26_, r_n_156__25_, r_n_156__24_, r_n_156__23_, r_n_156__22_, r_n_156__21_, r_n_156__20_, r_n_156__19_, r_n_156__18_, r_n_156__17_, r_n_156__16_, r_n_156__15_, r_n_156__14_, r_n_156__13_, r_n_156__12_, r_n_156__11_, r_n_156__10_, r_n_156__9_, r_n_156__8_, r_n_156__7_, r_n_156__6_, r_n_156__5_, r_n_156__4_, r_n_156__3_, r_n_156__2_, r_n_156__1_, r_n_156__0_ } = (N312)? { r_157__63_, r_157__62_, r_157__61_, r_157__60_, r_157__59_, r_157__58_, r_157__57_, r_157__56_, r_157__55_, r_157__54_, r_157__53_, r_157__52_, r_157__51_, r_157__50_, r_157__49_, r_157__48_, r_157__47_, r_157__46_, r_157__45_, r_157__44_, r_157__43_, r_157__42_, r_157__41_, r_157__40_, r_157__39_, r_157__38_, r_157__37_, r_157__36_, r_157__35_, r_157__34_, r_157__33_, r_157__32_, r_157__31_, r_157__30_, r_157__29_, r_157__28_, r_157__27_, r_157__26_, r_157__25_, r_157__24_, r_157__23_, r_157__22_, r_157__21_, r_157__20_, r_157__19_, r_157__18_, r_157__17_, r_157__16_, r_157__15_, r_157__14_, r_157__13_, r_157__12_, r_157__11_, r_157__10_, r_157__9_, r_157__8_, r_157__7_, r_157__6_, r_157__5_, r_157__4_, r_157__3_, r_157__2_, r_157__1_, r_157__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N313)? data_i : 1'b0;
  assign N312 = sel_i[312];
  assign N313 = N1808;
  assign { r_n_157__63_, r_n_157__62_, r_n_157__61_, r_n_157__60_, r_n_157__59_, r_n_157__58_, r_n_157__57_, r_n_157__56_, r_n_157__55_, r_n_157__54_, r_n_157__53_, r_n_157__52_, r_n_157__51_, r_n_157__50_, r_n_157__49_, r_n_157__48_, r_n_157__47_, r_n_157__46_, r_n_157__45_, r_n_157__44_, r_n_157__43_, r_n_157__42_, r_n_157__41_, r_n_157__40_, r_n_157__39_, r_n_157__38_, r_n_157__37_, r_n_157__36_, r_n_157__35_, r_n_157__34_, r_n_157__33_, r_n_157__32_, r_n_157__31_, r_n_157__30_, r_n_157__29_, r_n_157__28_, r_n_157__27_, r_n_157__26_, r_n_157__25_, r_n_157__24_, r_n_157__23_, r_n_157__22_, r_n_157__21_, r_n_157__20_, r_n_157__19_, r_n_157__18_, r_n_157__17_, r_n_157__16_, r_n_157__15_, r_n_157__14_, r_n_157__13_, r_n_157__12_, r_n_157__11_, r_n_157__10_, r_n_157__9_, r_n_157__8_, r_n_157__7_, r_n_157__6_, r_n_157__5_, r_n_157__4_, r_n_157__3_, r_n_157__2_, r_n_157__1_, r_n_157__0_ } = (N314)? { r_158__63_, r_158__62_, r_158__61_, r_158__60_, r_158__59_, r_158__58_, r_158__57_, r_158__56_, r_158__55_, r_158__54_, r_158__53_, r_158__52_, r_158__51_, r_158__50_, r_158__49_, r_158__48_, r_158__47_, r_158__46_, r_158__45_, r_158__44_, r_158__43_, r_158__42_, r_158__41_, r_158__40_, r_158__39_, r_158__38_, r_158__37_, r_158__36_, r_158__35_, r_158__34_, r_158__33_, r_158__32_, r_158__31_, r_158__30_, r_158__29_, r_158__28_, r_158__27_, r_158__26_, r_158__25_, r_158__24_, r_158__23_, r_158__22_, r_158__21_, r_158__20_, r_158__19_, r_158__18_, r_158__17_, r_158__16_, r_158__15_, r_158__14_, r_158__13_, r_158__12_, r_158__11_, r_158__10_, r_158__9_, r_158__8_, r_158__7_, r_158__6_, r_158__5_, r_158__4_, r_158__3_, r_158__2_, r_158__1_, r_158__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N315)? data_i : 1'b0;
  assign N314 = sel_i[314];
  assign N315 = N1813;
  assign { r_n_158__63_, r_n_158__62_, r_n_158__61_, r_n_158__60_, r_n_158__59_, r_n_158__58_, r_n_158__57_, r_n_158__56_, r_n_158__55_, r_n_158__54_, r_n_158__53_, r_n_158__52_, r_n_158__51_, r_n_158__50_, r_n_158__49_, r_n_158__48_, r_n_158__47_, r_n_158__46_, r_n_158__45_, r_n_158__44_, r_n_158__43_, r_n_158__42_, r_n_158__41_, r_n_158__40_, r_n_158__39_, r_n_158__38_, r_n_158__37_, r_n_158__36_, r_n_158__35_, r_n_158__34_, r_n_158__33_, r_n_158__32_, r_n_158__31_, r_n_158__30_, r_n_158__29_, r_n_158__28_, r_n_158__27_, r_n_158__26_, r_n_158__25_, r_n_158__24_, r_n_158__23_, r_n_158__22_, r_n_158__21_, r_n_158__20_, r_n_158__19_, r_n_158__18_, r_n_158__17_, r_n_158__16_, r_n_158__15_, r_n_158__14_, r_n_158__13_, r_n_158__12_, r_n_158__11_, r_n_158__10_, r_n_158__9_, r_n_158__8_, r_n_158__7_, r_n_158__6_, r_n_158__5_, r_n_158__4_, r_n_158__3_, r_n_158__2_, r_n_158__1_, r_n_158__0_ } = (N316)? { r_159__63_, r_159__62_, r_159__61_, r_159__60_, r_159__59_, r_159__58_, r_159__57_, r_159__56_, r_159__55_, r_159__54_, r_159__53_, r_159__52_, r_159__51_, r_159__50_, r_159__49_, r_159__48_, r_159__47_, r_159__46_, r_159__45_, r_159__44_, r_159__43_, r_159__42_, r_159__41_, r_159__40_, r_159__39_, r_159__38_, r_159__37_, r_159__36_, r_159__35_, r_159__34_, r_159__33_, r_159__32_, r_159__31_, r_159__30_, r_159__29_, r_159__28_, r_159__27_, r_159__26_, r_159__25_, r_159__24_, r_159__23_, r_159__22_, r_159__21_, r_159__20_, r_159__19_, r_159__18_, r_159__17_, r_159__16_, r_159__15_, r_159__14_, r_159__13_, r_159__12_, r_159__11_, r_159__10_, r_159__9_, r_159__8_, r_159__7_, r_159__6_, r_159__5_, r_159__4_, r_159__3_, r_159__2_, r_159__1_, r_159__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N317)? data_i : 1'b0;
  assign N316 = sel_i[316];
  assign N317 = N1818;
  assign { r_n_159__63_, r_n_159__62_, r_n_159__61_, r_n_159__60_, r_n_159__59_, r_n_159__58_, r_n_159__57_, r_n_159__56_, r_n_159__55_, r_n_159__54_, r_n_159__53_, r_n_159__52_, r_n_159__51_, r_n_159__50_, r_n_159__49_, r_n_159__48_, r_n_159__47_, r_n_159__46_, r_n_159__45_, r_n_159__44_, r_n_159__43_, r_n_159__42_, r_n_159__41_, r_n_159__40_, r_n_159__39_, r_n_159__38_, r_n_159__37_, r_n_159__36_, r_n_159__35_, r_n_159__34_, r_n_159__33_, r_n_159__32_, r_n_159__31_, r_n_159__30_, r_n_159__29_, r_n_159__28_, r_n_159__27_, r_n_159__26_, r_n_159__25_, r_n_159__24_, r_n_159__23_, r_n_159__22_, r_n_159__21_, r_n_159__20_, r_n_159__19_, r_n_159__18_, r_n_159__17_, r_n_159__16_, r_n_159__15_, r_n_159__14_, r_n_159__13_, r_n_159__12_, r_n_159__11_, r_n_159__10_, r_n_159__9_, r_n_159__8_, r_n_159__7_, r_n_159__6_, r_n_159__5_, r_n_159__4_, r_n_159__3_, r_n_159__2_, r_n_159__1_, r_n_159__0_ } = (N318)? { r_160__63_, r_160__62_, r_160__61_, r_160__60_, r_160__59_, r_160__58_, r_160__57_, r_160__56_, r_160__55_, r_160__54_, r_160__53_, r_160__52_, r_160__51_, r_160__50_, r_160__49_, r_160__48_, r_160__47_, r_160__46_, r_160__45_, r_160__44_, r_160__43_, r_160__42_, r_160__41_, r_160__40_, r_160__39_, r_160__38_, r_160__37_, r_160__36_, r_160__35_, r_160__34_, r_160__33_, r_160__32_, r_160__31_, r_160__30_, r_160__29_, r_160__28_, r_160__27_, r_160__26_, r_160__25_, r_160__24_, r_160__23_, r_160__22_, r_160__21_, r_160__20_, r_160__19_, r_160__18_, r_160__17_, r_160__16_, r_160__15_, r_160__14_, r_160__13_, r_160__12_, r_160__11_, r_160__10_, r_160__9_, r_160__8_, r_160__7_, r_160__6_, r_160__5_, r_160__4_, r_160__3_, r_160__2_, r_160__1_, r_160__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N319)? data_i : 1'b0;
  assign N318 = sel_i[318];
  assign N319 = N1823;
  assign { r_n_160__63_, r_n_160__62_, r_n_160__61_, r_n_160__60_, r_n_160__59_, r_n_160__58_, r_n_160__57_, r_n_160__56_, r_n_160__55_, r_n_160__54_, r_n_160__53_, r_n_160__52_, r_n_160__51_, r_n_160__50_, r_n_160__49_, r_n_160__48_, r_n_160__47_, r_n_160__46_, r_n_160__45_, r_n_160__44_, r_n_160__43_, r_n_160__42_, r_n_160__41_, r_n_160__40_, r_n_160__39_, r_n_160__38_, r_n_160__37_, r_n_160__36_, r_n_160__35_, r_n_160__34_, r_n_160__33_, r_n_160__32_, r_n_160__31_, r_n_160__30_, r_n_160__29_, r_n_160__28_, r_n_160__27_, r_n_160__26_, r_n_160__25_, r_n_160__24_, r_n_160__23_, r_n_160__22_, r_n_160__21_, r_n_160__20_, r_n_160__19_, r_n_160__18_, r_n_160__17_, r_n_160__16_, r_n_160__15_, r_n_160__14_, r_n_160__13_, r_n_160__12_, r_n_160__11_, r_n_160__10_, r_n_160__9_, r_n_160__8_, r_n_160__7_, r_n_160__6_, r_n_160__5_, r_n_160__4_, r_n_160__3_, r_n_160__2_, r_n_160__1_, r_n_160__0_ } = (N320)? { r_161__63_, r_161__62_, r_161__61_, r_161__60_, r_161__59_, r_161__58_, r_161__57_, r_161__56_, r_161__55_, r_161__54_, r_161__53_, r_161__52_, r_161__51_, r_161__50_, r_161__49_, r_161__48_, r_161__47_, r_161__46_, r_161__45_, r_161__44_, r_161__43_, r_161__42_, r_161__41_, r_161__40_, r_161__39_, r_161__38_, r_161__37_, r_161__36_, r_161__35_, r_161__34_, r_161__33_, r_161__32_, r_161__31_, r_161__30_, r_161__29_, r_161__28_, r_161__27_, r_161__26_, r_161__25_, r_161__24_, r_161__23_, r_161__22_, r_161__21_, r_161__20_, r_161__19_, r_161__18_, r_161__17_, r_161__16_, r_161__15_, r_161__14_, r_161__13_, r_161__12_, r_161__11_, r_161__10_, r_161__9_, r_161__8_, r_161__7_, r_161__6_, r_161__5_, r_161__4_, r_161__3_, r_161__2_, r_161__1_, r_161__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N321)? data_i : 1'b0;
  assign N320 = sel_i[320];
  assign N321 = N1828;
  assign { r_n_161__63_, r_n_161__62_, r_n_161__61_, r_n_161__60_, r_n_161__59_, r_n_161__58_, r_n_161__57_, r_n_161__56_, r_n_161__55_, r_n_161__54_, r_n_161__53_, r_n_161__52_, r_n_161__51_, r_n_161__50_, r_n_161__49_, r_n_161__48_, r_n_161__47_, r_n_161__46_, r_n_161__45_, r_n_161__44_, r_n_161__43_, r_n_161__42_, r_n_161__41_, r_n_161__40_, r_n_161__39_, r_n_161__38_, r_n_161__37_, r_n_161__36_, r_n_161__35_, r_n_161__34_, r_n_161__33_, r_n_161__32_, r_n_161__31_, r_n_161__30_, r_n_161__29_, r_n_161__28_, r_n_161__27_, r_n_161__26_, r_n_161__25_, r_n_161__24_, r_n_161__23_, r_n_161__22_, r_n_161__21_, r_n_161__20_, r_n_161__19_, r_n_161__18_, r_n_161__17_, r_n_161__16_, r_n_161__15_, r_n_161__14_, r_n_161__13_, r_n_161__12_, r_n_161__11_, r_n_161__10_, r_n_161__9_, r_n_161__8_, r_n_161__7_, r_n_161__6_, r_n_161__5_, r_n_161__4_, r_n_161__3_, r_n_161__2_, r_n_161__1_, r_n_161__0_ } = (N322)? { r_162__63_, r_162__62_, r_162__61_, r_162__60_, r_162__59_, r_162__58_, r_162__57_, r_162__56_, r_162__55_, r_162__54_, r_162__53_, r_162__52_, r_162__51_, r_162__50_, r_162__49_, r_162__48_, r_162__47_, r_162__46_, r_162__45_, r_162__44_, r_162__43_, r_162__42_, r_162__41_, r_162__40_, r_162__39_, r_162__38_, r_162__37_, r_162__36_, r_162__35_, r_162__34_, r_162__33_, r_162__32_, r_162__31_, r_162__30_, r_162__29_, r_162__28_, r_162__27_, r_162__26_, r_162__25_, r_162__24_, r_162__23_, r_162__22_, r_162__21_, r_162__20_, r_162__19_, r_162__18_, r_162__17_, r_162__16_, r_162__15_, r_162__14_, r_162__13_, r_162__12_, r_162__11_, r_162__10_, r_162__9_, r_162__8_, r_162__7_, r_162__6_, r_162__5_, r_162__4_, r_162__3_, r_162__2_, r_162__1_, r_162__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N323)? data_i : 1'b0;
  assign N322 = sel_i[322];
  assign N323 = N1833;
  assign { r_n_162__63_, r_n_162__62_, r_n_162__61_, r_n_162__60_, r_n_162__59_, r_n_162__58_, r_n_162__57_, r_n_162__56_, r_n_162__55_, r_n_162__54_, r_n_162__53_, r_n_162__52_, r_n_162__51_, r_n_162__50_, r_n_162__49_, r_n_162__48_, r_n_162__47_, r_n_162__46_, r_n_162__45_, r_n_162__44_, r_n_162__43_, r_n_162__42_, r_n_162__41_, r_n_162__40_, r_n_162__39_, r_n_162__38_, r_n_162__37_, r_n_162__36_, r_n_162__35_, r_n_162__34_, r_n_162__33_, r_n_162__32_, r_n_162__31_, r_n_162__30_, r_n_162__29_, r_n_162__28_, r_n_162__27_, r_n_162__26_, r_n_162__25_, r_n_162__24_, r_n_162__23_, r_n_162__22_, r_n_162__21_, r_n_162__20_, r_n_162__19_, r_n_162__18_, r_n_162__17_, r_n_162__16_, r_n_162__15_, r_n_162__14_, r_n_162__13_, r_n_162__12_, r_n_162__11_, r_n_162__10_, r_n_162__9_, r_n_162__8_, r_n_162__7_, r_n_162__6_, r_n_162__5_, r_n_162__4_, r_n_162__3_, r_n_162__2_, r_n_162__1_, r_n_162__0_ } = (N324)? { r_163__63_, r_163__62_, r_163__61_, r_163__60_, r_163__59_, r_163__58_, r_163__57_, r_163__56_, r_163__55_, r_163__54_, r_163__53_, r_163__52_, r_163__51_, r_163__50_, r_163__49_, r_163__48_, r_163__47_, r_163__46_, r_163__45_, r_163__44_, r_163__43_, r_163__42_, r_163__41_, r_163__40_, r_163__39_, r_163__38_, r_163__37_, r_163__36_, r_163__35_, r_163__34_, r_163__33_, r_163__32_, r_163__31_, r_163__30_, r_163__29_, r_163__28_, r_163__27_, r_163__26_, r_163__25_, r_163__24_, r_163__23_, r_163__22_, r_163__21_, r_163__20_, r_163__19_, r_163__18_, r_163__17_, r_163__16_, r_163__15_, r_163__14_, r_163__13_, r_163__12_, r_163__11_, r_163__10_, r_163__9_, r_163__8_, r_163__7_, r_163__6_, r_163__5_, r_163__4_, r_163__3_, r_163__2_, r_163__1_, r_163__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N325)? data_i : 1'b0;
  assign N324 = sel_i[324];
  assign N325 = N1838;
  assign { r_n_163__63_, r_n_163__62_, r_n_163__61_, r_n_163__60_, r_n_163__59_, r_n_163__58_, r_n_163__57_, r_n_163__56_, r_n_163__55_, r_n_163__54_, r_n_163__53_, r_n_163__52_, r_n_163__51_, r_n_163__50_, r_n_163__49_, r_n_163__48_, r_n_163__47_, r_n_163__46_, r_n_163__45_, r_n_163__44_, r_n_163__43_, r_n_163__42_, r_n_163__41_, r_n_163__40_, r_n_163__39_, r_n_163__38_, r_n_163__37_, r_n_163__36_, r_n_163__35_, r_n_163__34_, r_n_163__33_, r_n_163__32_, r_n_163__31_, r_n_163__30_, r_n_163__29_, r_n_163__28_, r_n_163__27_, r_n_163__26_, r_n_163__25_, r_n_163__24_, r_n_163__23_, r_n_163__22_, r_n_163__21_, r_n_163__20_, r_n_163__19_, r_n_163__18_, r_n_163__17_, r_n_163__16_, r_n_163__15_, r_n_163__14_, r_n_163__13_, r_n_163__12_, r_n_163__11_, r_n_163__10_, r_n_163__9_, r_n_163__8_, r_n_163__7_, r_n_163__6_, r_n_163__5_, r_n_163__4_, r_n_163__3_, r_n_163__2_, r_n_163__1_, r_n_163__0_ } = (N326)? { r_164__63_, r_164__62_, r_164__61_, r_164__60_, r_164__59_, r_164__58_, r_164__57_, r_164__56_, r_164__55_, r_164__54_, r_164__53_, r_164__52_, r_164__51_, r_164__50_, r_164__49_, r_164__48_, r_164__47_, r_164__46_, r_164__45_, r_164__44_, r_164__43_, r_164__42_, r_164__41_, r_164__40_, r_164__39_, r_164__38_, r_164__37_, r_164__36_, r_164__35_, r_164__34_, r_164__33_, r_164__32_, r_164__31_, r_164__30_, r_164__29_, r_164__28_, r_164__27_, r_164__26_, r_164__25_, r_164__24_, r_164__23_, r_164__22_, r_164__21_, r_164__20_, r_164__19_, r_164__18_, r_164__17_, r_164__16_, r_164__15_, r_164__14_, r_164__13_, r_164__12_, r_164__11_, r_164__10_, r_164__9_, r_164__8_, r_164__7_, r_164__6_, r_164__5_, r_164__4_, r_164__3_, r_164__2_, r_164__1_, r_164__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N327)? data_i : 1'b0;
  assign N326 = sel_i[326];
  assign N327 = N1843;
  assign { r_n_164__63_, r_n_164__62_, r_n_164__61_, r_n_164__60_, r_n_164__59_, r_n_164__58_, r_n_164__57_, r_n_164__56_, r_n_164__55_, r_n_164__54_, r_n_164__53_, r_n_164__52_, r_n_164__51_, r_n_164__50_, r_n_164__49_, r_n_164__48_, r_n_164__47_, r_n_164__46_, r_n_164__45_, r_n_164__44_, r_n_164__43_, r_n_164__42_, r_n_164__41_, r_n_164__40_, r_n_164__39_, r_n_164__38_, r_n_164__37_, r_n_164__36_, r_n_164__35_, r_n_164__34_, r_n_164__33_, r_n_164__32_, r_n_164__31_, r_n_164__30_, r_n_164__29_, r_n_164__28_, r_n_164__27_, r_n_164__26_, r_n_164__25_, r_n_164__24_, r_n_164__23_, r_n_164__22_, r_n_164__21_, r_n_164__20_, r_n_164__19_, r_n_164__18_, r_n_164__17_, r_n_164__16_, r_n_164__15_, r_n_164__14_, r_n_164__13_, r_n_164__12_, r_n_164__11_, r_n_164__10_, r_n_164__9_, r_n_164__8_, r_n_164__7_, r_n_164__6_, r_n_164__5_, r_n_164__4_, r_n_164__3_, r_n_164__2_, r_n_164__1_, r_n_164__0_ } = (N328)? { r_165__63_, r_165__62_, r_165__61_, r_165__60_, r_165__59_, r_165__58_, r_165__57_, r_165__56_, r_165__55_, r_165__54_, r_165__53_, r_165__52_, r_165__51_, r_165__50_, r_165__49_, r_165__48_, r_165__47_, r_165__46_, r_165__45_, r_165__44_, r_165__43_, r_165__42_, r_165__41_, r_165__40_, r_165__39_, r_165__38_, r_165__37_, r_165__36_, r_165__35_, r_165__34_, r_165__33_, r_165__32_, r_165__31_, r_165__30_, r_165__29_, r_165__28_, r_165__27_, r_165__26_, r_165__25_, r_165__24_, r_165__23_, r_165__22_, r_165__21_, r_165__20_, r_165__19_, r_165__18_, r_165__17_, r_165__16_, r_165__15_, r_165__14_, r_165__13_, r_165__12_, r_165__11_, r_165__10_, r_165__9_, r_165__8_, r_165__7_, r_165__6_, r_165__5_, r_165__4_, r_165__3_, r_165__2_, r_165__1_, r_165__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N329)? data_i : 1'b0;
  assign N328 = sel_i[328];
  assign N329 = N1848;
  assign { r_n_165__63_, r_n_165__62_, r_n_165__61_, r_n_165__60_, r_n_165__59_, r_n_165__58_, r_n_165__57_, r_n_165__56_, r_n_165__55_, r_n_165__54_, r_n_165__53_, r_n_165__52_, r_n_165__51_, r_n_165__50_, r_n_165__49_, r_n_165__48_, r_n_165__47_, r_n_165__46_, r_n_165__45_, r_n_165__44_, r_n_165__43_, r_n_165__42_, r_n_165__41_, r_n_165__40_, r_n_165__39_, r_n_165__38_, r_n_165__37_, r_n_165__36_, r_n_165__35_, r_n_165__34_, r_n_165__33_, r_n_165__32_, r_n_165__31_, r_n_165__30_, r_n_165__29_, r_n_165__28_, r_n_165__27_, r_n_165__26_, r_n_165__25_, r_n_165__24_, r_n_165__23_, r_n_165__22_, r_n_165__21_, r_n_165__20_, r_n_165__19_, r_n_165__18_, r_n_165__17_, r_n_165__16_, r_n_165__15_, r_n_165__14_, r_n_165__13_, r_n_165__12_, r_n_165__11_, r_n_165__10_, r_n_165__9_, r_n_165__8_, r_n_165__7_, r_n_165__6_, r_n_165__5_, r_n_165__4_, r_n_165__3_, r_n_165__2_, r_n_165__1_, r_n_165__0_ } = (N330)? { r_166__63_, r_166__62_, r_166__61_, r_166__60_, r_166__59_, r_166__58_, r_166__57_, r_166__56_, r_166__55_, r_166__54_, r_166__53_, r_166__52_, r_166__51_, r_166__50_, r_166__49_, r_166__48_, r_166__47_, r_166__46_, r_166__45_, r_166__44_, r_166__43_, r_166__42_, r_166__41_, r_166__40_, r_166__39_, r_166__38_, r_166__37_, r_166__36_, r_166__35_, r_166__34_, r_166__33_, r_166__32_, r_166__31_, r_166__30_, r_166__29_, r_166__28_, r_166__27_, r_166__26_, r_166__25_, r_166__24_, r_166__23_, r_166__22_, r_166__21_, r_166__20_, r_166__19_, r_166__18_, r_166__17_, r_166__16_, r_166__15_, r_166__14_, r_166__13_, r_166__12_, r_166__11_, r_166__10_, r_166__9_, r_166__8_, r_166__7_, r_166__6_, r_166__5_, r_166__4_, r_166__3_, r_166__2_, r_166__1_, r_166__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N331)? data_i : 1'b0;
  assign N330 = sel_i[330];
  assign N331 = N1853;
  assign { r_n_166__63_, r_n_166__62_, r_n_166__61_, r_n_166__60_, r_n_166__59_, r_n_166__58_, r_n_166__57_, r_n_166__56_, r_n_166__55_, r_n_166__54_, r_n_166__53_, r_n_166__52_, r_n_166__51_, r_n_166__50_, r_n_166__49_, r_n_166__48_, r_n_166__47_, r_n_166__46_, r_n_166__45_, r_n_166__44_, r_n_166__43_, r_n_166__42_, r_n_166__41_, r_n_166__40_, r_n_166__39_, r_n_166__38_, r_n_166__37_, r_n_166__36_, r_n_166__35_, r_n_166__34_, r_n_166__33_, r_n_166__32_, r_n_166__31_, r_n_166__30_, r_n_166__29_, r_n_166__28_, r_n_166__27_, r_n_166__26_, r_n_166__25_, r_n_166__24_, r_n_166__23_, r_n_166__22_, r_n_166__21_, r_n_166__20_, r_n_166__19_, r_n_166__18_, r_n_166__17_, r_n_166__16_, r_n_166__15_, r_n_166__14_, r_n_166__13_, r_n_166__12_, r_n_166__11_, r_n_166__10_, r_n_166__9_, r_n_166__8_, r_n_166__7_, r_n_166__6_, r_n_166__5_, r_n_166__4_, r_n_166__3_, r_n_166__2_, r_n_166__1_, r_n_166__0_ } = (N332)? { r_167__63_, r_167__62_, r_167__61_, r_167__60_, r_167__59_, r_167__58_, r_167__57_, r_167__56_, r_167__55_, r_167__54_, r_167__53_, r_167__52_, r_167__51_, r_167__50_, r_167__49_, r_167__48_, r_167__47_, r_167__46_, r_167__45_, r_167__44_, r_167__43_, r_167__42_, r_167__41_, r_167__40_, r_167__39_, r_167__38_, r_167__37_, r_167__36_, r_167__35_, r_167__34_, r_167__33_, r_167__32_, r_167__31_, r_167__30_, r_167__29_, r_167__28_, r_167__27_, r_167__26_, r_167__25_, r_167__24_, r_167__23_, r_167__22_, r_167__21_, r_167__20_, r_167__19_, r_167__18_, r_167__17_, r_167__16_, r_167__15_, r_167__14_, r_167__13_, r_167__12_, r_167__11_, r_167__10_, r_167__9_, r_167__8_, r_167__7_, r_167__6_, r_167__5_, r_167__4_, r_167__3_, r_167__2_, r_167__1_, r_167__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N333)? data_i : 1'b0;
  assign N332 = sel_i[332];
  assign N333 = N1858;
  assign { r_n_167__63_, r_n_167__62_, r_n_167__61_, r_n_167__60_, r_n_167__59_, r_n_167__58_, r_n_167__57_, r_n_167__56_, r_n_167__55_, r_n_167__54_, r_n_167__53_, r_n_167__52_, r_n_167__51_, r_n_167__50_, r_n_167__49_, r_n_167__48_, r_n_167__47_, r_n_167__46_, r_n_167__45_, r_n_167__44_, r_n_167__43_, r_n_167__42_, r_n_167__41_, r_n_167__40_, r_n_167__39_, r_n_167__38_, r_n_167__37_, r_n_167__36_, r_n_167__35_, r_n_167__34_, r_n_167__33_, r_n_167__32_, r_n_167__31_, r_n_167__30_, r_n_167__29_, r_n_167__28_, r_n_167__27_, r_n_167__26_, r_n_167__25_, r_n_167__24_, r_n_167__23_, r_n_167__22_, r_n_167__21_, r_n_167__20_, r_n_167__19_, r_n_167__18_, r_n_167__17_, r_n_167__16_, r_n_167__15_, r_n_167__14_, r_n_167__13_, r_n_167__12_, r_n_167__11_, r_n_167__10_, r_n_167__9_, r_n_167__8_, r_n_167__7_, r_n_167__6_, r_n_167__5_, r_n_167__4_, r_n_167__3_, r_n_167__2_, r_n_167__1_, r_n_167__0_ } = (N334)? { r_168__63_, r_168__62_, r_168__61_, r_168__60_, r_168__59_, r_168__58_, r_168__57_, r_168__56_, r_168__55_, r_168__54_, r_168__53_, r_168__52_, r_168__51_, r_168__50_, r_168__49_, r_168__48_, r_168__47_, r_168__46_, r_168__45_, r_168__44_, r_168__43_, r_168__42_, r_168__41_, r_168__40_, r_168__39_, r_168__38_, r_168__37_, r_168__36_, r_168__35_, r_168__34_, r_168__33_, r_168__32_, r_168__31_, r_168__30_, r_168__29_, r_168__28_, r_168__27_, r_168__26_, r_168__25_, r_168__24_, r_168__23_, r_168__22_, r_168__21_, r_168__20_, r_168__19_, r_168__18_, r_168__17_, r_168__16_, r_168__15_, r_168__14_, r_168__13_, r_168__12_, r_168__11_, r_168__10_, r_168__9_, r_168__8_, r_168__7_, r_168__6_, r_168__5_, r_168__4_, r_168__3_, r_168__2_, r_168__1_, r_168__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N335)? data_i : 1'b0;
  assign N334 = sel_i[334];
  assign N335 = N1863;
  assign { r_n_168__63_, r_n_168__62_, r_n_168__61_, r_n_168__60_, r_n_168__59_, r_n_168__58_, r_n_168__57_, r_n_168__56_, r_n_168__55_, r_n_168__54_, r_n_168__53_, r_n_168__52_, r_n_168__51_, r_n_168__50_, r_n_168__49_, r_n_168__48_, r_n_168__47_, r_n_168__46_, r_n_168__45_, r_n_168__44_, r_n_168__43_, r_n_168__42_, r_n_168__41_, r_n_168__40_, r_n_168__39_, r_n_168__38_, r_n_168__37_, r_n_168__36_, r_n_168__35_, r_n_168__34_, r_n_168__33_, r_n_168__32_, r_n_168__31_, r_n_168__30_, r_n_168__29_, r_n_168__28_, r_n_168__27_, r_n_168__26_, r_n_168__25_, r_n_168__24_, r_n_168__23_, r_n_168__22_, r_n_168__21_, r_n_168__20_, r_n_168__19_, r_n_168__18_, r_n_168__17_, r_n_168__16_, r_n_168__15_, r_n_168__14_, r_n_168__13_, r_n_168__12_, r_n_168__11_, r_n_168__10_, r_n_168__9_, r_n_168__8_, r_n_168__7_, r_n_168__6_, r_n_168__5_, r_n_168__4_, r_n_168__3_, r_n_168__2_, r_n_168__1_, r_n_168__0_ } = (N336)? { r_169__63_, r_169__62_, r_169__61_, r_169__60_, r_169__59_, r_169__58_, r_169__57_, r_169__56_, r_169__55_, r_169__54_, r_169__53_, r_169__52_, r_169__51_, r_169__50_, r_169__49_, r_169__48_, r_169__47_, r_169__46_, r_169__45_, r_169__44_, r_169__43_, r_169__42_, r_169__41_, r_169__40_, r_169__39_, r_169__38_, r_169__37_, r_169__36_, r_169__35_, r_169__34_, r_169__33_, r_169__32_, r_169__31_, r_169__30_, r_169__29_, r_169__28_, r_169__27_, r_169__26_, r_169__25_, r_169__24_, r_169__23_, r_169__22_, r_169__21_, r_169__20_, r_169__19_, r_169__18_, r_169__17_, r_169__16_, r_169__15_, r_169__14_, r_169__13_, r_169__12_, r_169__11_, r_169__10_, r_169__9_, r_169__8_, r_169__7_, r_169__6_, r_169__5_, r_169__4_, r_169__3_, r_169__2_, r_169__1_, r_169__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N337)? data_i : 1'b0;
  assign N336 = sel_i[336];
  assign N337 = N1868;
  assign { r_n_169__63_, r_n_169__62_, r_n_169__61_, r_n_169__60_, r_n_169__59_, r_n_169__58_, r_n_169__57_, r_n_169__56_, r_n_169__55_, r_n_169__54_, r_n_169__53_, r_n_169__52_, r_n_169__51_, r_n_169__50_, r_n_169__49_, r_n_169__48_, r_n_169__47_, r_n_169__46_, r_n_169__45_, r_n_169__44_, r_n_169__43_, r_n_169__42_, r_n_169__41_, r_n_169__40_, r_n_169__39_, r_n_169__38_, r_n_169__37_, r_n_169__36_, r_n_169__35_, r_n_169__34_, r_n_169__33_, r_n_169__32_, r_n_169__31_, r_n_169__30_, r_n_169__29_, r_n_169__28_, r_n_169__27_, r_n_169__26_, r_n_169__25_, r_n_169__24_, r_n_169__23_, r_n_169__22_, r_n_169__21_, r_n_169__20_, r_n_169__19_, r_n_169__18_, r_n_169__17_, r_n_169__16_, r_n_169__15_, r_n_169__14_, r_n_169__13_, r_n_169__12_, r_n_169__11_, r_n_169__10_, r_n_169__9_, r_n_169__8_, r_n_169__7_, r_n_169__6_, r_n_169__5_, r_n_169__4_, r_n_169__3_, r_n_169__2_, r_n_169__1_, r_n_169__0_ } = (N338)? { r_170__63_, r_170__62_, r_170__61_, r_170__60_, r_170__59_, r_170__58_, r_170__57_, r_170__56_, r_170__55_, r_170__54_, r_170__53_, r_170__52_, r_170__51_, r_170__50_, r_170__49_, r_170__48_, r_170__47_, r_170__46_, r_170__45_, r_170__44_, r_170__43_, r_170__42_, r_170__41_, r_170__40_, r_170__39_, r_170__38_, r_170__37_, r_170__36_, r_170__35_, r_170__34_, r_170__33_, r_170__32_, r_170__31_, r_170__30_, r_170__29_, r_170__28_, r_170__27_, r_170__26_, r_170__25_, r_170__24_, r_170__23_, r_170__22_, r_170__21_, r_170__20_, r_170__19_, r_170__18_, r_170__17_, r_170__16_, r_170__15_, r_170__14_, r_170__13_, r_170__12_, r_170__11_, r_170__10_, r_170__9_, r_170__8_, r_170__7_, r_170__6_, r_170__5_, r_170__4_, r_170__3_, r_170__2_, r_170__1_, r_170__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N339)? data_i : 1'b0;
  assign N338 = sel_i[338];
  assign N339 = N1873;
  assign { r_n_170__63_, r_n_170__62_, r_n_170__61_, r_n_170__60_, r_n_170__59_, r_n_170__58_, r_n_170__57_, r_n_170__56_, r_n_170__55_, r_n_170__54_, r_n_170__53_, r_n_170__52_, r_n_170__51_, r_n_170__50_, r_n_170__49_, r_n_170__48_, r_n_170__47_, r_n_170__46_, r_n_170__45_, r_n_170__44_, r_n_170__43_, r_n_170__42_, r_n_170__41_, r_n_170__40_, r_n_170__39_, r_n_170__38_, r_n_170__37_, r_n_170__36_, r_n_170__35_, r_n_170__34_, r_n_170__33_, r_n_170__32_, r_n_170__31_, r_n_170__30_, r_n_170__29_, r_n_170__28_, r_n_170__27_, r_n_170__26_, r_n_170__25_, r_n_170__24_, r_n_170__23_, r_n_170__22_, r_n_170__21_, r_n_170__20_, r_n_170__19_, r_n_170__18_, r_n_170__17_, r_n_170__16_, r_n_170__15_, r_n_170__14_, r_n_170__13_, r_n_170__12_, r_n_170__11_, r_n_170__10_, r_n_170__9_, r_n_170__8_, r_n_170__7_, r_n_170__6_, r_n_170__5_, r_n_170__4_, r_n_170__3_, r_n_170__2_, r_n_170__1_, r_n_170__0_ } = (N340)? { r_171__63_, r_171__62_, r_171__61_, r_171__60_, r_171__59_, r_171__58_, r_171__57_, r_171__56_, r_171__55_, r_171__54_, r_171__53_, r_171__52_, r_171__51_, r_171__50_, r_171__49_, r_171__48_, r_171__47_, r_171__46_, r_171__45_, r_171__44_, r_171__43_, r_171__42_, r_171__41_, r_171__40_, r_171__39_, r_171__38_, r_171__37_, r_171__36_, r_171__35_, r_171__34_, r_171__33_, r_171__32_, r_171__31_, r_171__30_, r_171__29_, r_171__28_, r_171__27_, r_171__26_, r_171__25_, r_171__24_, r_171__23_, r_171__22_, r_171__21_, r_171__20_, r_171__19_, r_171__18_, r_171__17_, r_171__16_, r_171__15_, r_171__14_, r_171__13_, r_171__12_, r_171__11_, r_171__10_, r_171__9_, r_171__8_, r_171__7_, r_171__6_, r_171__5_, r_171__4_, r_171__3_, r_171__2_, r_171__1_, r_171__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N341)? data_i : 1'b0;
  assign N340 = sel_i[340];
  assign N341 = N1878;
  assign { r_n_171__63_, r_n_171__62_, r_n_171__61_, r_n_171__60_, r_n_171__59_, r_n_171__58_, r_n_171__57_, r_n_171__56_, r_n_171__55_, r_n_171__54_, r_n_171__53_, r_n_171__52_, r_n_171__51_, r_n_171__50_, r_n_171__49_, r_n_171__48_, r_n_171__47_, r_n_171__46_, r_n_171__45_, r_n_171__44_, r_n_171__43_, r_n_171__42_, r_n_171__41_, r_n_171__40_, r_n_171__39_, r_n_171__38_, r_n_171__37_, r_n_171__36_, r_n_171__35_, r_n_171__34_, r_n_171__33_, r_n_171__32_, r_n_171__31_, r_n_171__30_, r_n_171__29_, r_n_171__28_, r_n_171__27_, r_n_171__26_, r_n_171__25_, r_n_171__24_, r_n_171__23_, r_n_171__22_, r_n_171__21_, r_n_171__20_, r_n_171__19_, r_n_171__18_, r_n_171__17_, r_n_171__16_, r_n_171__15_, r_n_171__14_, r_n_171__13_, r_n_171__12_, r_n_171__11_, r_n_171__10_, r_n_171__9_, r_n_171__8_, r_n_171__7_, r_n_171__6_, r_n_171__5_, r_n_171__4_, r_n_171__3_, r_n_171__2_, r_n_171__1_, r_n_171__0_ } = (N342)? { r_172__63_, r_172__62_, r_172__61_, r_172__60_, r_172__59_, r_172__58_, r_172__57_, r_172__56_, r_172__55_, r_172__54_, r_172__53_, r_172__52_, r_172__51_, r_172__50_, r_172__49_, r_172__48_, r_172__47_, r_172__46_, r_172__45_, r_172__44_, r_172__43_, r_172__42_, r_172__41_, r_172__40_, r_172__39_, r_172__38_, r_172__37_, r_172__36_, r_172__35_, r_172__34_, r_172__33_, r_172__32_, r_172__31_, r_172__30_, r_172__29_, r_172__28_, r_172__27_, r_172__26_, r_172__25_, r_172__24_, r_172__23_, r_172__22_, r_172__21_, r_172__20_, r_172__19_, r_172__18_, r_172__17_, r_172__16_, r_172__15_, r_172__14_, r_172__13_, r_172__12_, r_172__11_, r_172__10_, r_172__9_, r_172__8_, r_172__7_, r_172__6_, r_172__5_, r_172__4_, r_172__3_, r_172__2_, r_172__1_, r_172__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N343)? data_i : 1'b0;
  assign N342 = sel_i[342];
  assign N343 = N1883;
  assign { r_n_172__63_, r_n_172__62_, r_n_172__61_, r_n_172__60_, r_n_172__59_, r_n_172__58_, r_n_172__57_, r_n_172__56_, r_n_172__55_, r_n_172__54_, r_n_172__53_, r_n_172__52_, r_n_172__51_, r_n_172__50_, r_n_172__49_, r_n_172__48_, r_n_172__47_, r_n_172__46_, r_n_172__45_, r_n_172__44_, r_n_172__43_, r_n_172__42_, r_n_172__41_, r_n_172__40_, r_n_172__39_, r_n_172__38_, r_n_172__37_, r_n_172__36_, r_n_172__35_, r_n_172__34_, r_n_172__33_, r_n_172__32_, r_n_172__31_, r_n_172__30_, r_n_172__29_, r_n_172__28_, r_n_172__27_, r_n_172__26_, r_n_172__25_, r_n_172__24_, r_n_172__23_, r_n_172__22_, r_n_172__21_, r_n_172__20_, r_n_172__19_, r_n_172__18_, r_n_172__17_, r_n_172__16_, r_n_172__15_, r_n_172__14_, r_n_172__13_, r_n_172__12_, r_n_172__11_, r_n_172__10_, r_n_172__9_, r_n_172__8_, r_n_172__7_, r_n_172__6_, r_n_172__5_, r_n_172__4_, r_n_172__3_, r_n_172__2_, r_n_172__1_, r_n_172__0_ } = (N344)? { r_173__63_, r_173__62_, r_173__61_, r_173__60_, r_173__59_, r_173__58_, r_173__57_, r_173__56_, r_173__55_, r_173__54_, r_173__53_, r_173__52_, r_173__51_, r_173__50_, r_173__49_, r_173__48_, r_173__47_, r_173__46_, r_173__45_, r_173__44_, r_173__43_, r_173__42_, r_173__41_, r_173__40_, r_173__39_, r_173__38_, r_173__37_, r_173__36_, r_173__35_, r_173__34_, r_173__33_, r_173__32_, r_173__31_, r_173__30_, r_173__29_, r_173__28_, r_173__27_, r_173__26_, r_173__25_, r_173__24_, r_173__23_, r_173__22_, r_173__21_, r_173__20_, r_173__19_, r_173__18_, r_173__17_, r_173__16_, r_173__15_, r_173__14_, r_173__13_, r_173__12_, r_173__11_, r_173__10_, r_173__9_, r_173__8_, r_173__7_, r_173__6_, r_173__5_, r_173__4_, r_173__3_, r_173__2_, r_173__1_, r_173__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N345)? data_i : 1'b0;
  assign N344 = sel_i[344];
  assign N345 = N1888;
  assign { r_n_173__63_, r_n_173__62_, r_n_173__61_, r_n_173__60_, r_n_173__59_, r_n_173__58_, r_n_173__57_, r_n_173__56_, r_n_173__55_, r_n_173__54_, r_n_173__53_, r_n_173__52_, r_n_173__51_, r_n_173__50_, r_n_173__49_, r_n_173__48_, r_n_173__47_, r_n_173__46_, r_n_173__45_, r_n_173__44_, r_n_173__43_, r_n_173__42_, r_n_173__41_, r_n_173__40_, r_n_173__39_, r_n_173__38_, r_n_173__37_, r_n_173__36_, r_n_173__35_, r_n_173__34_, r_n_173__33_, r_n_173__32_, r_n_173__31_, r_n_173__30_, r_n_173__29_, r_n_173__28_, r_n_173__27_, r_n_173__26_, r_n_173__25_, r_n_173__24_, r_n_173__23_, r_n_173__22_, r_n_173__21_, r_n_173__20_, r_n_173__19_, r_n_173__18_, r_n_173__17_, r_n_173__16_, r_n_173__15_, r_n_173__14_, r_n_173__13_, r_n_173__12_, r_n_173__11_, r_n_173__10_, r_n_173__9_, r_n_173__8_, r_n_173__7_, r_n_173__6_, r_n_173__5_, r_n_173__4_, r_n_173__3_, r_n_173__2_, r_n_173__1_, r_n_173__0_ } = (N346)? { r_174__63_, r_174__62_, r_174__61_, r_174__60_, r_174__59_, r_174__58_, r_174__57_, r_174__56_, r_174__55_, r_174__54_, r_174__53_, r_174__52_, r_174__51_, r_174__50_, r_174__49_, r_174__48_, r_174__47_, r_174__46_, r_174__45_, r_174__44_, r_174__43_, r_174__42_, r_174__41_, r_174__40_, r_174__39_, r_174__38_, r_174__37_, r_174__36_, r_174__35_, r_174__34_, r_174__33_, r_174__32_, r_174__31_, r_174__30_, r_174__29_, r_174__28_, r_174__27_, r_174__26_, r_174__25_, r_174__24_, r_174__23_, r_174__22_, r_174__21_, r_174__20_, r_174__19_, r_174__18_, r_174__17_, r_174__16_, r_174__15_, r_174__14_, r_174__13_, r_174__12_, r_174__11_, r_174__10_, r_174__9_, r_174__8_, r_174__7_, r_174__6_, r_174__5_, r_174__4_, r_174__3_, r_174__2_, r_174__1_, r_174__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N347)? data_i : 1'b0;
  assign N346 = sel_i[346];
  assign N347 = N1893;
  assign { r_n_174__63_, r_n_174__62_, r_n_174__61_, r_n_174__60_, r_n_174__59_, r_n_174__58_, r_n_174__57_, r_n_174__56_, r_n_174__55_, r_n_174__54_, r_n_174__53_, r_n_174__52_, r_n_174__51_, r_n_174__50_, r_n_174__49_, r_n_174__48_, r_n_174__47_, r_n_174__46_, r_n_174__45_, r_n_174__44_, r_n_174__43_, r_n_174__42_, r_n_174__41_, r_n_174__40_, r_n_174__39_, r_n_174__38_, r_n_174__37_, r_n_174__36_, r_n_174__35_, r_n_174__34_, r_n_174__33_, r_n_174__32_, r_n_174__31_, r_n_174__30_, r_n_174__29_, r_n_174__28_, r_n_174__27_, r_n_174__26_, r_n_174__25_, r_n_174__24_, r_n_174__23_, r_n_174__22_, r_n_174__21_, r_n_174__20_, r_n_174__19_, r_n_174__18_, r_n_174__17_, r_n_174__16_, r_n_174__15_, r_n_174__14_, r_n_174__13_, r_n_174__12_, r_n_174__11_, r_n_174__10_, r_n_174__9_, r_n_174__8_, r_n_174__7_, r_n_174__6_, r_n_174__5_, r_n_174__4_, r_n_174__3_, r_n_174__2_, r_n_174__1_, r_n_174__0_ } = (N348)? { r_175__63_, r_175__62_, r_175__61_, r_175__60_, r_175__59_, r_175__58_, r_175__57_, r_175__56_, r_175__55_, r_175__54_, r_175__53_, r_175__52_, r_175__51_, r_175__50_, r_175__49_, r_175__48_, r_175__47_, r_175__46_, r_175__45_, r_175__44_, r_175__43_, r_175__42_, r_175__41_, r_175__40_, r_175__39_, r_175__38_, r_175__37_, r_175__36_, r_175__35_, r_175__34_, r_175__33_, r_175__32_, r_175__31_, r_175__30_, r_175__29_, r_175__28_, r_175__27_, r_175__26_, r_175__25_, r_175__24_, r_175__23_, r_175__22_, r_175__21_, r_175__20_, r_175__19_, r_175__18_, r_175__17_, r_175__16_, r_175__15_, r_175__14_, r_175__13_, r_175__12_, r_175__11_, r_175__10_, r_175__9_, r_175__8_, r_175__7_, r_175__6_, r_175__5_, r_175__4_, r_175__3_, r_175__2_, r_175__1_, r_175__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N349)? data_i : 1'b0;
  assign N348 = sel_i[348];
  assign N349 = N1898;
  assign { r_n_175__63_, r_n_175__62_, r_n_175__61_, r_n_175__60_, r_n_175__59_, r_n_175__58_, r_n_175__57_, r_n_175__56_, r_n_175__55_, r_n_175__54_, r_n_175__53_, r_n_175__52_, r_n_175__51_, r_n_175__50_, r_n_175__49_, r_n_175__48_, r_n_175__47_, r_n_175__46_, r_n_175__45_, r_n_175__44_, r_n_175__43_, r_n_175__42_, r_n_175__41_, r_n_175__40_, r_n_175__39_, r_n_175__38_, r_n_175__37_, r_n_175__36_, r_n_175__35_, r_n_175__34_, r_n_175__33_, r_n_175__32_, r_n_175__31_, r_n_175__30_, r_n_175__29_, r_n_175__28_, r_n_175__27_, r_n_175__26_, r_n_175__25_, r_n_175__24_, r_n_175__23_, r_n_175__22_, r_n_175__21_, r_n_175__20_, r_n_175__19_, r_n_175__18_, r_n_175__17_, r_n_175__16_, r_n_175__15_, r_n_175__14_, r_n_175__13_, r_n_175__12_, r_n_175__11_, r_n_175__10_, r_n_175__9_, r_n_175__8_, r_n_175__7_, r_n_175__6_, r_n_175__5_, r_n_175__4_, r_n_175__3_, r_n_175__2_, r_n_175__1_, r_n_175__0_ } = (N350)? { r_176__63_, r_176__62_, r_176__61_, r_176__60_, r_176__59_, r_176__58_, r_176__57_, r_176__56_, r_176__55_, r_176__54_, r_176__53_, r_176__52_, r_176__51_, r_176__50_, r_176__49_, r_176__48_, r_176__47_, r_176__46_, r_176__45_, r_176__44_, r_176__43_, r_176__42_, r_176__41_, r_176__40_, r_176__39_, r_176__38_, r_176__37_, r_176__36_, r_176__35_, r_176__34_, r_176__33_, r_176__32_, r_176__31_, r_176__30_, r_176__29_, r_176__28_, r_176__27_, r_176__26_, r_176__25_, r_176__24_, r_176__23_, r_176__22_, r_176__21_, r_176__20_, r_176__19_, r_176__18_, r_176__17_, r_176__16_, r_176__15_, r_176__14_, r_176__13_, r_176__12_, r_176__11_, r_176__10_, r_176__9_, r_176__8_, r_176__7_, r_176__6_, r_176__5_, r_176__4_, r_176__3_, r_176__2_, r_176__1_, r_176__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N351)? data_i : 1'b0;
  assign N350 = sel_i[350];
  assign N351 = N1903;
  assign { r_n_176__63_, r_n_176__62_, r_n_176__61_, r_n_176__60_, r_n_176__59_, r_n_176__58_, r_n_176__57_, r_n_176__56_, r_n_176__55_, r_n_176__54_, r_n_176__53_, r_n_176__52_, r_n_176__51_, r_n_176__50_, r_n_176__49_, r_n_176__48_, r_n_176__47_, r_n_176__46_, r_n_176__45_, r_n_176__44_, r_n_176__43_, r_n_176__42_, r_n_176__41_, r_n_176__40_, r_n_176__39_, r_n_176__38_, r_n_176__37_, r_n_176__36_, r_n_176__35_, r_n_176__34_, r_n_176__33_, r_n_176__32_, r_n_176__31_, r_n_176__30_, r_n_176__29_, r_n_176__28_, r_n_176__27_, r_n_176__26_, r_n_176__25_, r_n_176__24_, r_n_176__23_, r_n_176__22_, r_n_176__21_, r_n_176__20_, r_n_176__19_, r_n_176__18_, r_n_176__17_, r_n_176__16_, r_n_176__15_, r_n_176__14_, r_n_176__13_, r_n_176__12_, r_n_176__11_, r_n_176__10_, r_n_176__9_, r_n_176__8_, r_n_176__7_, r_n_176__6_, r_n_176__5_, r_n_176__4_, r_n_176__3_, r_n_176__2_, r_n_176__1_, r_n_176__0_ } = (N352)? { r_177__63_, r_177__62_, r_177__61_, r_177__60_, r_177__59_, r_177__58_, r_177__57_, r_177__56_, r_177__55_, r_177__54_, r_177__53_, r_177__52_, r_177__51_, r_177__50_, r_177__49_, r_177__48_, r_177__47_, r_177__46_, r_177__45_, r_177__44_, r_177__43_, r_177__42_, r_177__41_, r_177__40_, r_177__39_, r_177__38_, r_177__37_, r_177__36_, r_177__35_, r_177__34_, r_177__33_, r_177__32_, r_177__31_, r_177__30_, r_177__29_, r_177__28_, r_177__27_, r_177__26_, r_177__25_, r_177__24_, r_177__23_, r_177__22_, r_177__21_, r_177__20_, r_177__19_, r_177__18_, r_177__17_, r_177__16_, r_177__15_, r_177__14_, r_177__13_, r_177__12_, r_177__11_, r_177__10_, r_177__9_, r_177__8_, r_177__7_, r_177__6_, r_177__5_, r_177__4_, r_177__3_, r_177__2_, r_177__1_, r_177__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N353)? data_i : 1'b0;
  assign N352 = sel_i[352];
  assign N353 = N1908;
  assign { r_n_177__63_, r_n_177__62_, r_n_177__61_, r_n_177__60_, r_n_177__59_, r_n_177__58_, r_n_177__57_, r_n_177__56_, r_n_177__55_, r_n_177__54_, r_n_177__53_, r_n_177__52_, r_n_177__51_, r_n_177__50_, r_n_177__49_, r_n_177__48_, r_n_177__47_, r_n_177__46_, r_n_177__45_, r_n_177__44_, r_n_177__43_, r_n_177__42_, r_n_177__41_, r_n_177__40_, r_n_177__39_, r_n_177__38_, r_n_177__37_, r_n_177__36_, r_n_177__35_, r_n_177__34_, r_n_177__33_, r_n_177__32_, r_n_177__31_, r_n_177__30_, r_n_177__29_, r_n_177__28_, r_n_177__27_, r_n_177__26_, r_n_177__25_, r_n_177__24_, r_n_177__23_, r_n_177__22_, r_n_177__21_, r_n_177__20_, r_n_177__19_, r_n_177__18_, r_n_177__17_, r_n_177__16_, r_n_177__15_, r_n_177__14_, r_n_177__13_, r_n_177__12_, r_n_177__11_, r_n_177__10_, r_n_177__9_, r_n_177__8_, r_n_177__7_, r_n_177__6_, r_n_177__5_, r_n_177__4_, r_n_177__3_, r_n_177__2_, r_n_177__1_, r_n_177__0_ } = (N354)? { r_178__63_, r_178__62_, r_178__61_, r_178__60_, r_178__59_, r_178__58_, r_178__57_, r_178__56_, r_178__55_, r_178__54_, r_178__53_, r_178__52_, r_178__51_, r_178__50_, r_178__49_, r_178__48_, r_178__47_, r_178__46_, r_178__45_, r_178__44_, r_178__43_, r_178__42_, r_178__41_, r_178__40_, r_178__39_, r_178__38_, r_178__37_, r_178__36_, r_178__35_, r_178__34_, r_178__33_, r_178__32_, r_178__31_, r_178__30_, r_178__29_, r_178__28_, r_178__27_, r_178__26_, r_178__25_, r_178__24_, r_178__23_, r_178__22_, r_178__21_, r_178__20_, r_178__19_, r_178__18_, r_178__17_, r_178__16_, r_178__15_, r_178__14_, r_178__13_, r_178__12_, r_178__11_, r_178__10_, r_178__9_, r_178__8_, r_178__7_, r_178__6_, r_178__5_, r_178__4_, r_178__3_, r_178__2_, r_178__1_, r_178__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N355)? data_i : 1'b0;
  assign N354 = sel_i[354];
  assign N355 = N1913;
  assign { r_n_178__63_, r_n_178__62_, r_n_178__61_, r_n_178__60_, r_n_178__59_, r_n_178__58_, r_n_178__57_, r_n_178__56_, r_n_178__55_, r_n_178__54_, r_n_178__53_, r_n_178__52_, r_n_178__51_, r_n_178__50_, r_n_178__49_, r_n_178__48_, r_n_178__47_, r_n_178__46_, r_n_178__45_, r_n_178__44_, r_n_178__43_, r_n_178__42_, r_n_178__41_, r_n_178__40_, r_n_178__39_, r_n_178__38_, r_n_178__37_, r_n_178__36_, r_n_178__35_, r_n_178__34_, r_n_178__33_, r_n_178__32_, r_n_178__31_, r_n_178__30_, r_n_178__29_, r_n_178__28_, r_n_178__27_, r_n_178__26_, r_n_178__25_, r_n_178__24_, r_n_178__23_, r_n_178__22_, r_n_178__21_, r_n_178__20_, r_n_178__19_, r_n_178__18_, r_n_178__17_, r_n_178__16_, r_n_178__15_, r_n_178__14_, r_n_178__13_, r_n_178__12_, r_n_178__11_, r_n_178__10_, r_n_178__9_, r_n_178__8_, r_n_178__7_, r_n_178__6_, r_n_178__5_, r_n_178__4_, r_n_178__3_, r_n_178__2_, r_n_178__1_, r_n_178__0_ } = (N356)? { r_179__63_, r_179__62_, r_179__61_, r_179__60_, r_179__59_, r_179__58_, r_179__57_, r_179__56_, r_179__55_, r_179__54_, r_179__53_, r_179__52_, r_179__51_, r_179__50_, r_179__49_, r_179__48_, r_179__47_, r_179__46_, r_179__45_, r_179__44_, r_179__43_, r_179__42_, r_179__41_, r_179__40_, r_179__39_, r_179__38_, r_179__37_, r_179__36_, r_179__35_, r_179__34_, r_179__33_, r_179__32_, r_179__31_, r_179__30_, r_179__29_, r_179__28_, r_179__27_, r_179__26_, r_179__25_, r_179__24_, r_179__23_, r_179__22_, r_179__21_, r_179__20_, r_179__19_, r_179__18_, r_179__17_, r_179__16_, r_179__15_, r_179__14_, r_179__13_, r_179__12_, r_179__11_, r_179__10_, r_179__9_, r_179__8_, r_179__7_, r_179__6_, r_179__5_, r_179__4_, r_179__3_, r_179__2_, r_179__1_, r_179__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N357)? data_i : 1'b0;
  assign N356 = sel_i[356];
  assign N357 = N1918;
  assign { r_n_179__63_, r_n_179__62_, r_n_179__61_, r_n_179__60_, r_n_179__59_, r_n_179__58_, r_n_179__57_, r_n_179__56_, r_n_179__55_, r_n_179__54_, r_n_179__53_, r_n_179__52_, r_n_179__51_, r_n_179__50_, r_n_179__49_, r_n_179__48_, r_n_179__47_, r_n_179__46_, r_n_179__45_, r_n_179__44_, r_n_179__43_, r_n_179__42_, r_n_179__41_, r_n_179__40_, r_n_179__39_, r_n_179__38_, r_n_179__37_, r_n_179__36_, r_n_179__35_, r_n_179__34_, r_n_179__33_, r_n_179__32_, r_n_179__31_, r_n_179__30_, r_n_179__29_, r_n_179__28_, r_n_179__27_, r_n_179__26_, r_n_179__25_, r_n_179__24_, r_n_179__23_, r_n_179__22_, r_n_179__21_, r_n_179__20_, r_n_179__19_, r_n_179__18_, r_n_179__17_, r_n_179__16_, r_n_179__15_, r_n_179__14_, r_n_179__13_, r_n_179__12_, r_n_179__11_, r_n_179__10_, r_n_179__9_, r_n_179__8_, r_n_179__7_, r_n_179__6_, r_n_179__5_, r_n_179__4_, r_n_179__3_, r_n_179__2_, r_n_179__1_, r_n_179__0_ } = (N358)? { r_180__63_, r_180__62_, r_180__61_, r_180__60_, r_180__59_, r_180__58_, r_180__57_, r_180__56_, r_180__55_, r_180__54_, r_180__53_, r_180__52_, r_180__51_, r_180__50_, r_180__49_, r_180__48_, r_180__47_, r_180__46_, r_180__45_, r_180__44_, r_180__43_, r_180__42_, r_180__41_, r_180__40_, r_180__39_, r_180__38_, r_180__37_, r_180__36_, r_180__35_, r_180__34_, r_180__33_, r_180__32_, r_180__31_, r_180__30_, r_180__29_, r_180__28_, r_180__27_, r_180__26_, r_180__25_, r_180__24_, r_180__23_, r_180__22_, r_180__21_, r_180__20_, r_180__19_, r_180__18_, r_180__17_, r_180__16_, r_180__15_, r_180__14_, r_180__13_, r_180__12_, r_180__11_, r_180__10_, r_180__9_, r_180__8_, r_180__7_, r_180__6_, r_180__5_, r_180__4_, r_180__3_, r_180__2_, r_180__1_, r_180__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N359)? data_i : 1'b0;
  assign N358 = sel_i[358];
  assign N359 = N1923;
  assign { r_n_180__63_, r_n_180__62_, r_n_180__61_, r_n_180__60_, r_n_180__59_, r_n_180__58_, r_n_180__57_, r_n_180__56_, r_n_180__55_, r_n_180__54_, r_n_180__53_, r_n_180__52_, r_n_180__51_, r_n_180__50_, r_n_180__49_, r_n_180__48_, r_n_180__47_, r_n_180__46_, r_n_180__45_, r_n_180__44_, r_n_180__43_, r_n_180__42_, r_n_180__41_, r_n_180__40_, r_n_180__39_, r_n_180__38_, r_n_180__37_, r_n_180__36_, r_n_180__35_, r_n_180__34_, r_n_180__33_, r_n_180__32_, r_n_180__31_, r_n_180__30_, r_n_180__29_, r_n_180__28_, r_n_180__27_, r_n_180__26_, r_n_180__25_, r_n_180__24_, r_n_180__23_, r_n_180__22_, r_n_180__21_, r_n_180__20_, r_n_180__19_, r_n_180__18_, r_n_180__17_, r_n_180__16_, r_n_180__15_, r_n_180__14_, r_n_180__13_, r_n_180__12_, r_n_180__11_, r_n_180__10_, r_n_180__9_, r_n_180__8_, r_n_180__7_, r_n_180__6_, r_n_180__5_, r_n_180__4_, r_n_180__3_, r_n_180__2_, r_n_180__1_, r_n_180__0_ } = (N360)? { r_181__63_, r_181__62_, r_181__61_, r_181__60_, r_181__59_, r_181__58_, r_181__57_, r_181__56_, r_181__55_, r_181__54_, r_181__53_, r_181__52_, r_181__51_, r_181__50_, r_181__49_, r_181__48_, r_181__47_, r_181__46_, r_181__45_, r_181__44_, r_181__43_, r_181__42_, r_181__41_, r_181__40_, r_181__39_, r_181__38_, r_181__37_, r_181__36_, r_181__35_, r_181__34_, r_181__33_, r_181__32_, r_181__31_, r_181__30_, r_181__29_, r_181__28_, r_181__27_, r_181__26_, r_181__25_, r_181__24_, r_181__23_, r_181__22_, r_181__21_, r_181__20_, r_181__19_, r_181__18_, r_181__17_, r_181__16_, r_181__15_, r_181__14_, r_181__13_, r_181__12_, r_181__11_, r_181__10_, r_181__9_, r_181__8_, r_181__7_, r_181__6_, r_181__5_, r_181__4_, r_181__3_, r_181__2_, r_181__1_, r_181__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N361)? data_i : 1'b0;
  assign N360 = sel_i[360];
  assign N361 = N1928;
  assign { r_n_181__63_, r_n_181__62_, r_n_181__61_, r_n_181__60_, r_n_181__59_, r_n_181__58_, r_n_181__57_, r_n_181__56_, r_n_181__55_, r_n_181__54_, r_n_181__53_, r_n_181__52_, r_n_181__51_, r_n_181__50_, r_n_181__49_, r_n_181__48_, r_n_181__47_, r_n_181__46_, r_n_181__45_, r_n_181__44_, r_n_181__43_, r_n_181__42_, r_n_181__41_, r_n_181__40_, r_n_181__39_, r_n_181__38_, r_n_181__37_, r_n_181__36_, r_n_181__35_, r_n_181__34_, r_n_181__33_, r_n_181__32_, r_n_181__31_, r_n_181__30_, r_n_181__29_, r_n_181__28_, r_n_181__27_, r_n_181__26_, r_n_181__25_, r_n_181__24_, r_n_181__23_, r_n_181__22_, r_n_181__21_, r_n_181__20_, r_n_181__19_, r_n_181__18_, r_n_181__17_, r_n_181__16_, r_n_181__15_, r_n_181__14_, r_n_181__13_, r_n_181__12_, r_n_181__11_, r_n_181__10_, r_n_181__9_, r_n_181__8_, r_n_181__7_, r_n_181__6_, r_n_181__5_, r_n_181__4_, r_n_181__3_, r_n_181__2_, r_n_181__1_, r_n_181__0_ } = (N362)? { r_182__63_, r_182__62_, r_182__61_, r_182__60_, r_182__59_, r_182__58_, r_182__57_, r_182__56_, r_182__55_, r_182__54_, r_182__53_, r_182__52_, r_182__51_, r_182__50_, r_182__49_, r_182__48_, r_182__47_, r_182__46_, r_182__45_, r_182__44_, r_182__43_, r_182__42_, r_182__41_, r_182__40_, r_182__39_, r_182__38_, r_182__37_, r_182__36_, r_182__35_, r_182__34_, r_182__33_, r_182__32_, r_182__31_, r_182__30_, r_182__29_, r_182__28_, r_182__27_, r_182__26_, r_182__25_, r_182__24_, r_182__23_, r_182__22_, r_182__21_, r_182__20_, r_182__19_, r_182__18_, r_182__17_, r_182__16_, r_182__15_, r_182__14_, r_182__13_, r_182__12_, r_182__11_, r_182__10_, r_182__9_, r_182__8_, r_182__7_, r_182__6_, r_182__5_, r_182__4_, r_182__3_, r_182__2_, r_182__1_, r_182__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N363)? data_i : 1'b0;
  assign N362 = sel_i[362];
  assign N363 = N1933;
  assign { r_n_182__63_, r_n_182__62_, r_n_182__61_, r_n_182__60_, r_n_182__59_, r_n_182__58_, r_n_182__57_, r_n_182__56_, r_n_182__55_, r_n_182__54_, r_n_182__53_, r_n_182__52_, r_n_182__51_, r_n_182__50_, r_n_182__49_, r_n_182__48_, r_n_182__47_, r_n_182__46_, r_n_182__45_, r_n_182__44_, r_n_182__43_, r_n_182__42_, r_n_182__41_, r_n_182__40_, r_n_182__39_, r_n_182__38_, r_n_182__37_, r_n_182__36_, r_n_182__35_, r_n_182__34_, r_n_182__33_, r_n_182__32_, r_n_182__31_, r_n_182__30_, r_n_182__29_, r_n_182__28_, r_n_182__27_, r_n_182__26_, r_n_182__25_, r_n_182__24_, r_n_182__23_, r_n_182__22_, r_n_182__21_, r_n_182__20_, r_n_182__19_, r_n_182__18_, r_n_182__17_, r_n_182__16_, r_n_182__15_, r_n_182__14_, r_n_182__13_, r_n_182__12_, r_n_182__11_, r_n_182__10_, r_n_182__9_, r_n_182__8_, r_n_182__7_, r_n_182__6_, r_n_182__5_, r_n_182__4_, r_n_182__3_, r_n_182__2_, r_n_182__1_, r_n_182__0_ } = (N364)? { r_183__63_, r_183__62_, r_183__61_, r_183__60_, r_183__59_, r_183__58_, r_183__57_, r_183__56_, r_183__55_, r_183__54_, r_183__53_, r_183__52_, r_183__51_, r_183__50_, r_183__49_, r_183__48_, r_183__47_, r_183__46_, r_183__45_, r_183__44_, r_183__43_, r_183__42_, r_183__41_, r_183__40_, r_183__39_, r_183__38_, r_183__37_, r_183__36_, r_183__35_, r_183__34_, r_183__33_, r_183__32_, r_183__31_, r_183__30_, r_183__29_, r_183__28_, r_183__27_, r_183__26_, r_183__25_, r_183__24_, r_183__23_, r_183__22_, r_183__21_, r_183__20_, r_183__19_, r_183__18_, r_183__17_, r_183__16_, r_183__15_, r_183__14_, r_183__13_, r_183__12_, r_183__11_, r_183__10_, r_183__9_, r_183__8_, r_183__7_, r_183__6_, r_183__5_, r_183__4_, r_183__3_, r_183__2_, r_183__1_, r_183__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N365)? data_i : 1'b0;
  assign N364 = sel_i[364];
  assign N365 = N1938;
  assign { r_n_183__63_, r_n_183__62_, r_n_183__61_, r_n_183__60_, r_n_183__59_, r_n_183__58_, r_n_183__57_, r_n_183__56_, r_n_183__55_, r_n_183__54_, r_n_183__53_, r_n_183__52_, r_n_183__51_, r_n_183__50_, r_n_183__49_, r_n_183__48_, r_n_183__47_, r_n_183__46_, r_n_183__45_, r_n_183__44_, r_n_183__43_, r_n_183__42_, r_n_183__41_, r_n_183__40_, r_n_183__39_, r_n_183__38_, r_n_183__37_, r_n_183__36_, r_n_183__35_, r_n_183__34_, r_n_183__33_, r_n_183__32_, r_n_183__31_, r_n_183__30_, r_n_183__29_, r_n_183__28_, r_n_183__27_, r_n_183__26_, r_n_183__25_, r_n_183__24_, r_n_183__23_, r_n_183__22_, r_n_183__21_, r_n_183__20_, r_n_183__19_, r_n_183__18_, r_n_183__17_, r_n_183__16_, r_n_183__15_, r_n_183__14_, r_n_183__13_, r_n_183__12_, r_n_183__11_, r_n_183__10_, r_n_183__9_, r_n_183__8_, r_n_183__7_, r_n_183__6_, r_n_183__5_, r_n_183__4_, r_n_183__3_, r_n_183__2_, r_n_183__1_, r_n_183__0_ } = (N366)? { r_184__63_, r_184__62_, r_184__61_, r_184__60_, r_184__59_, r_184__58_, r_184__57_, r_184__56_, r_184__55_, r_184__54_, r_184__53_, r_184__52_, r_184__51_, r_184__50_, r_184__49_, r_184__48_, r_184__47_, r_184__46_, r_184__45_, r_184__44_, r_184__43_, r_184__42_, r_184__41_, r_184__40_, r_184__39_, r_184__38_, r_184__37_, r_184__36_, r_184__35_, r_184__34_, r_184__33_, r_184__32_, r_184__31_, r_184__30_, r_184__29_, r_184__28_, r_184__27_, r_184__26_, r_184__25_, r_184__24_, r_184__23_, r_184__22_, r_184__21_, r_184__20_, r_184__19_, r_184__18_, r_184__17_, r_184__16_, r_184__15_, r_184__14_, r_184__13_, r_184__12_, r_184__11_, r_184__10_, r_184__9_, r_184__8_, r_184__7_, r_184__6_, r_184__5_, r_184__4_, r_184__3_, r_184__2_, r_184__1_, r_184__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N367)? data_i : 1'b0;
  assign N366 = sel_i[366];
  assign N367 = N1943;
  assign { r_n_184__63_, r_n_184__62_, r_n_184__61_, r_n_184__60_, r_n_184__59_, r_n_184__58_, r_n_184__57_, r_n_184__56_, r_n_184__55_, r_n_184__54_, r_n_184__53_, r_n_184__52_, r_n_184__51_, r_n_184__50_, r_n_184__49_, r_n_184__48_, r_n_184__47_, r_n_184__46_, r_n_184__45_, r_n_184__44_, r_n_184__43_, r_n_184__42_, r_n_184__41_, r_n_184__40_, r_n_184__39_, r_n_184__38_, r_n_184__37_, r_n_184__36_, r_n_184__35_, r_n_184__34_, r_n_184__33_, r_n_184__32_, r_n_184__31_, r_n_184__30_, r_n_184__29_, r_n_184__28_, r_n_184__27_, r_n_184__26_, r_n_184__25_, r_n_184__24_, r_n_184__23_, r_n_184__22_, r_n_184__21_, r_n_184__20_, r_n_184__19_, r_n_184__18_, r_n_184__17_, r_n_184__16_, r_n_184__15_, r_n_184__14_, r_n_184__13_, r_n_184__12_, r_n_184__11_, r_n_184__10_, r_n_184__9_, r_n_184__8_, r_n_184__7_, r_n_184__6_, r_n_184__5_, r_n_184__4_, r_n_184__3_, r_n_184__2_, r_n_184__1_, r_n_184__0_ } = (N368)? { r_185__63_, r_185__62_, r_185__61_, r_185__60_, r_185__59_, r_185__58_, r_185__57_, r_185__56_, r_185__55_, r_185__54_, r_185__53_, r_185__52_, r_185__51_, r_185__50_, r_185__49_, r_185__48_, r_185__47_, r_185__46_, r_185__45_, r_185__44_, r_185__43_, r_185__42_, r_185__41_, r_185__40_, r_185__39_, r_185__38_, r_185__37_, r_185__36_, r_185__35_, r_185__34_, r_185__33_, r_185__32_, r_185__31_, r_185__30_, r_185__29_, r_185__28_, r_185__27_, r_185__26_, r_185__25_, r_185__24_, r_185__23_, r_185__22_, r_185__21_, r_185__20_, r_185__19_, r_185__18_, r_185__17_, r_185__16_, r_185__15_, r_185__14_, r_185__13_, r_185__12_, r_185__11_, r_185__10_, r_185__9_, r_185__8_, r_185__7_, r_185__6_, r_185__5_, r_185__4_, r_185__3_, r_185__2_, r_185__1_, r_185__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N369)? data_i : 1'b0;
  assign N368 = sel_i[368];
  assign N369 = N1948;
  assign { r_n_185__63_, r_n_185__62_, r_n_185__61_, r_n_185__60_, r_n_185__59_, r_n_185__58_, r_n_185__57_, r_n_185__56_, r_n_185__55_, r_n_185__54_, r_n_185__53_, r_n_185__52_, r_n_185__51_, r_n_185__50_, r_n_185__49_, r_n_185__48_, r_n_185__47_, r_n_185__46_, r_n_185__45_, r_n_185__44_, r_n_185__43_, r_n_185__42_, r_n_185__41_, r_n_185__40_, r_n_185__39_, r_n_185__38_, r_n_185__37_, r_n_185__36_, r_n_185__35_, r_n_185__34_, r_n_185__33_, r_n_185__32_, r_n_185__31_, r_n_185__30_, r_n_185__29_, r_n_185__28_, r_n_185__27_, r_n_185__26_, r_n_185__25_, r_n_185__24_, r_n_185__23_, r_n_185__22_, r_n_185__21_, r_n_185__20_, r_n_185__19_, r_n_185__18_, r_n_185__17_, r_n_185__16_, r_n_185__15_, r_n_185__14_, r_n_185__13_, r_n_185__12_, r_n_185__11_, r_n_185__10_, r_n_185__9_, r_n_185__8_, r_n_185__7_, r_n_185__6_, r_n_185__5_, r_n_185__4_, r_n_185__3_, r_n_185__2_, r_n_185__1_, r_n_185__0_ } = (N370)? { r_186__63_, r_186__62_, r_186__61_, r_186__60_, r_186__59_, r_186__58_, r_186__57_, r_186__56_, r_186__55_, r_186__54_, r_186__53_, r_186__52_, r_186__51_, r_186__50_, r_186__49_, r_186__48_, r_186__47_, r_186__46_, r_186__45_, r_186__44_, r_186__43_, r_186__42_, r_186__41_, r_186__40_, r_186__39_, r_186__38_, r_186__37_, r_186__36_, r_186__35_, r_186__34_, r_186__33_, r_186__32_, r_186__31_, r_186__30_, r_186__29_, r_186__28_, r_186__27_, r_186__26_, r_186__25_, r_186__24_, r_186__23_, r_186__22_, r_186__21_, r_186__20_, r_186__19_, r_186__18_, r_186__17_, r_186__16_, r_186__15_, r_186__14_, r_186__13_, r_186__12_, r_186__11_, r_186__10_, r_186__9_, r_186__8_, r_186__7_, r_186__6_, r_186__5_, r_186__4_, r_186__3_, r_186__2_, r_186__1_, r_186__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N371)? data_i : 1'b0;
  assign N370 = sel_i[370];
  assign N371 = N1953;
  assign { r_n_186__63_, r_n_186__62_, r_n_186__61_, r_n_186__60_, r_n_186__59_, r_n_186__58_, r_n_186__57_, r_n_186__56_, r_n_186__55_, r_n_186__54_, r_n_186__53_, r_n_186__52_, r_n_186__51_, r_n_186__50_, r_n_186__49_, r_n_186__48_, r_n_186__47_, r_n_186__46_, r_n_186__45_, r_n_186__44_, r_n_186__43_, r_n_186__42_, r_n_186__41_, r_n_186__40_, r_n_186__39_, r_n_186__38_, r_n_186__37_, r_n_186__36_, r_n_186__35_, r_n_186__34_, r_n_186__33_, r_n_186__32_, r_n_186__31_, r_n_186__30_, r_n_186__29_, r_n_186__28_, r_n_186__27_, r_n_186__26_, r_n_186__25_, r_n_186__24_, r_n_186__23_, r_n_186__22_, r_n_186__21_, r_n_186__20_, r_n_186__19_, r_n_186__18_, r_n_186__17_, r_n_186__16_, r_n_186__15_, r_n_186__14_, r_n_186__13_, r_n_186__12_, r_n_186__11_, r_n_186__10_, r_n_186__9_, r_n_186__8_, r_n_186__7_, r_n_186__6_, r_n_186__5_, r_n_186__4_, r_n_186__3_, r_n_186__2_, r_n_186__1_, r_n_186__0_ } = (N372)? { r_187__63_, r_187__62_, r_187__61_, r_187__60_, r_187__59_, r_187__58_, r_187__57_, r_187__56_, r_187__55_, r_187__54_, r_187__53_, r_187__52_, r_187__51_, r_187__50_, r_187__49_, r_187__48_, r_187__47_, r_187__46_, r_187__45_, r_187__44_, r_187__43_, r_187__42_, r_187__41_, r_187__40_, r_187__39_, r_187__38_, r_187__37_, r_187__36_, r_187__35_, r_187__34_, r_187__33_, r_187__32_, r_187__31_, r_187__30_, r_187__29_, r_187__28_, r_187__27_, r_187__26_, r_187__25_, r_187__24_, r_187__23_, r_187__22_, r_187__21_, r_187__20_, r_187__19_, r_187__18_, r_187__17_, r_187__16_, r_187__15_, r_187__14_, r_187__13_, r_187__12_, r_187__11_, r_187__10_, r_187__9_, r_187__8_, r_187__7_, r_187__6_, r_187__5_, r_187__4_, r_187__3_, r_187__2_, r_187__1_, r_187__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N373)? data_i : 1'b0;
  assign N372 = sel_i[372];
  assign N373 = N1958;
  assign { r_n_187__63_, r_n_187__62_, r_n_187__61_, r_n_187__60_, r_n_187__59_, r_n_187__58_, r_n_187__57_, r_n_187__56_, r_n_187__55_, r_n_187__54_, r_n_187__53_, r_n_187__52_, r_n_187__51_, r_n_187__50_, r_n_187__49_, r_n_187__48_, r_n_187__47_, r_n_187__46_, r_n_187__45_, r_n_187__44_, r_n_187__43_, r_n_187__42_, r_n_187__41_, r_n_187__40_, r_n_187__39_, r_n_187__38_, r_n_187__37_, r_n_187__36_, r_n_187__35_, r_n_187__34_, r_n_187__33_, r_n_187__32_, r_n_187__31_, r_n_187__30_, r_n_187__29_, r_n_187__28_, r_n_187__27_, r_n_187__26_, r_n_187__25_, r_n_187__24_, r_n_187__23_, r_n_187__22_, r_n_187__21_, r_n_187__20_, r_n_187__19_, r_n_187__18_, r_n_187__17_, r_n_187__16_, r_n_187__15_, r_n_187__14_, r_n_187__13_, r_n_187__12_, r_n_187__11_, r_n_187__10_, r_n_187__9_, r_n_187__8_, r_n_187__7_, r_n_187__6_, r_n_187__5_, r_n_187__4_, r_n_187__3_, r_n_187__2_, r_n_187__1_, r_n_187__0_ } = (N374)? { r_188__63_, r_188__62_, r_188__61_, r_188__60_, r_188__59_, r_188__58_, r_188__57_, r_188__56_, r_188__55_, r_188__54_, r_188__53_, r_188__52_, r_188__51_, r_188__50_, r_188__49_, r_188__48_, r_188__47_, r_188__46_, r_188__45_, r_188__44_, r_188__43_, r_188__42_, r_188__41_, r_188__40_, r_188__39_, r_188__38_, r_188__37_, r_188__36_, r_188__35_, r_188__34_, r_188__33_, r_188__32_, r_188__31_, r_188__30_, r_188__29_, r_188__28_, r_188__27_, r_188__26_, r_188__25_, r_188__24_, r_188__23_, r_188__22_, r_188__21_, r_188__20_, r_188__19_, r_188__18_, r_188__17_, r_188__16_, r_188__15_, r_188__14_, r_188__13_, r_188__12_, r_188__11_, r_188__10_, r_188__9_, r_188__8_, r_188__7_, r_188__6_, r_188__5_, r_188__4_, r_188__3_, r_188__2_, r_188__1_, r_188__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N375)? data_i : 1'b0;
  assign N374 = sel_i[374];
  assign N375 = N1963;
  assign { r_n_188__63_, r_n_188__62_, r_n_188__61_, r_n_188__60_, r_n_188__59_, r_n_188__58_, r_n_188__57_, r_n_188__56_, r_n_188__55_, r_n_188__54_, r_n_188__53_, r_n_188__52_, r_n_188__51_, r_n_188__50_, r_n_188__49_, r_n_188__48_, r_n_188__47_, r_n_188__46_, r_n_188__45_, r_n_188__44_, r_n_188__43_, r_n_188__42_, r_n_188__41_, r_n_188__40_, r_n_188__39_, r_n_188__38_, r_n_188__37_, r_n_188__36_, r_n_188__35_, r_n_188__34_, r_n_188__33_, r_n_188__32_, r_n_188__31_, r_n_188__30_, r_n_188__29_, r_n_188__28_, r_n_188__27_, r_n_188__26_, r_n_188__25_, r_n_188__24_, r_n_188__23_, r_n_188__22_, r_n_188__21_, r_n_188__20_, r_n_188__19_, r_n_188__18_, r_n_188__17_, r_n_188__16_, r_n_188__15_, r_n_188__14_, r_n_188__13_, r_n_188__12_, r_n_188__11_, r_n_188__10_, r_n_188__9_, r_n_188__8_, r_n_188__7_, r_n_188__6_, r_n_188__5_, r_n_188__4_, r_n_188__3_, r_n_188__2_, r_n_188__1_, r_n_188__0_ } = (N376)? { r_189__63_, r_189__62_, r_189__61_, r_189__60_, r_189__59_, r_189__58_, r_189__57_, r_189__56_, r_189__55_, r_189__54_, r_189__53_, r_189__52_, r_189__51_, r_189__50_, r_189__49_, r_189__48_, r_189__47_, r_189__46_, r_189__45_, r_189__44_, r_189__43_, r_189__42_, r_189__41_, r_189__40_, r_189__39_, r_189__38_, r_189__37_, r_189__36_, r_189__35_, r_189__34_, r_189__33_, r_189__32_, r_189__31_, r_189__30_, r_189__29_, r_189__28_, r_189__27_, r_189__26_, r_189__25_, r_189__24_, r_189__23_, r_189__22_, r_189__21_, r_189__20_, r_189__19_, r_189__18_, r_189__17_, r_189__16_, r_189__15_, r_189__14_, r_189__13_, r_189__12_, r_189__11_, r_189__10_, r_189__9_, r_189__8_, r_189__7_, r_189__6_, r_189__5_, r_189__4_, r_189__3_, r_189__2_, r_189__1_, r_189__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N377)? data_i : 1'b0;
  assign N376 = sel_i[376];
  assign N377 = N1968;
  assign { r_n_189__63_, r_n_189__62_, r_n_189__61_, r_n_189__60_, r_n_189__59_, r_n_189__58_, r_n_189__57_, r_n_189__56_, r_n_189__55_, r_n_189__54_, r_n_189__53_, r_n_189__52_, r_n_189__51_, r_n_189__50_, r_n_189__49_, r_n_189__48_, r_n_189__47_, r_n_189__46_, r_n_189__45_, r_n_189__44_, r_n_189__43_, r_n_189__42_, r_n_189__41_, r_n_189__40_, r_n_189__39_, r_n_189__38_, r_n_189__37_, r_n_189__36_, r_n_189__35_, r_n_189__34_, r_n_189__33_, r_n_189__32_, r_n_189__31_, r_n_189__30_, r_n_189__29_, r_n_189__28_, r_n_189__27_, r_n_189__26_, r_n_189__25_, r_n_189__24_, r_n_189__23_, r_n_189__22_, r_n_189__21_, r_n_189__20_, r_n_189__19_, r_n_189__18_, r_n_189__17_, r_n_189__16_, r_n_189__15_, r_n_189__14_, r_n_189__13_, r_n_189__12_, r_n_189__11_, r_n_189__10_, r_n_189__9_, r_n_189__8_, r_n_189__7_, r_n_189__6_, r_n_189__5_, r_n_189__4_, r_n_189__3_, r_n_189__2_, r_n_189__1_, r_n_189__0_ } = (N378)? { r_190__63_, r_190__62_, r_190__61_, r_190__60_, r_190__59_, r_190__58_, r_190__57_, r_190__56_, r_190__55_, r_190__54_, r_190__53_, r_190__52_, r_190__51_, r_190__50_, r_190__49_, r_190__48_, r_190__47_, r_190__46_, r_190__45_, r_190__44_, r_190__43_, r_190__42_, r_190__41_, r_190__40_, r_190__39_, r_190__38_, r_190__37_, r_190__36_, r_190__35_, r_190__34_, r_190__33_, r_190__32_, r_190__31_, r_190__30_, r_190__29_, r_190__28_, r_190__27_, r_190__26_, r_190__25_, r_190__24_, r_190__23_, r_190__22_, r_190__21_, r_190__20_, r_190__19_, r_190__18_, r_190__17_, r_190__16_, r_190__15_, r_190__14_, r_190__13_, r_190__12_, r_190__11_, r_190__10_, r_190__9_, r_190__8_, r_190__7_, r_190__6_, r_190__5_, r_190__4_, r_190__3_, r_190__2_, r_190__1_, r_190__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N379)? data_i : 1'b0;
  assign N378 = sel_i[378];
  assign N379 = N1973;
  assign { r_n_190__63_, r_n_190__62_, r_n_190__61_, r_n_190__60_, r_n_190__59_, r_n_190__58_, r_n_190__57_, r_n_190__56_, r_n_190__55_, r_n_190__54_, r_n_190__53_, r_n_190__52_, r_n_190__51_, r_n_190__50_, r_n_190__49_, r_n_190__48_, r_n_190__47_, r_n_190__46_, r_n_190__45_, r_n_190__44_, r_n_190__43_, r_n_190__42_, r_n_190__41_, r_n_190__40_, r_n_190__39_, r_n_190__38_, r_n_190__37_, r_n_190__36_, r_n_190__35_, r_n_190__34_, r_n_190__33_, r_n_190__32_, r_n_190__31_, r_n_190__30_, r_n_190__29_, r_n_190__28_, r_n_190__27_, r_n_190__26_, r_n_190__25_, r_n_190__24_, r_n_190__23_, r_n_190__22_, r_n_190__21_, r_n_190__20_, r_n_190__19_, r_n_190__18_, r_n_190__17_, r_n_190__16_, r_n_190__15_, r_n_190__14_, r_n_190__13_, r_n_190__12_, r_n_190__11_, r_n_190__10_, r_n_190__9_, r_n_190__8_, r_n_190__7_, r_n_190__6_, r_n_190__5_, r_n_190__4_, r_n_190__3_, r_n_190__2_, r_n_190__1_, r_n_190__0_ } = (N380)? { r_191__63_, r_191__62_, r_191__61_, r_191__60_, r_191__59_, r_191__58_, r_191__57_, r_191__56_, r_191__55_, r_191__54_, r_191__53_, r_191__52_, r_191__51_, r_191__50_, r_191__49_, r_191__48_, r_191__47_, r_191__46_, r_191__45_, r_191__44_, r_191__43_, r_191__42_, r_191__41_, r_191__40_, r_191__39_, r_191__38_, r_191__37_, r_191__36_, r_191__35_, r_191__34_, r_191__33_, r_191__32_, r_191__31_, r_191__30_, r_191__29_, r_191__28_, r_191__27_, r_191__26_, r_191__25_, r_191__24_, r_191__23_, r_191__22_, r_191__21_, r_191__20_, r_191__19_, r_191__18_, r_191__17_, r_191__16_, r_191__15_, r_191__14_, r_191__13_, r_191__12_, r_191__11_, r_191__10_, r_191__9_, r_191__8_, r_191__7_, r_191__6_, r_191__5_, r_191__4_, r_191__3_, r_191__2_, r_191__1_, r_191__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N381)? data_i : 1'b0;
  assign N380 = sel_i[380];
  assign N381 = N1978;
  assign { r_n_191__63_, r_n_191__62_, r_n_191__61_, r_n_191__60_, r_n_191__59_, r_n_191__58_, r_n_191__57_, r_n_191__56_, r_n_191__55_, r_n_191__54_, r_n_191__53_, r_n_191__52_, r_n_191__51_, r_n_191__50_, r_n_191__49_, r_n_191__48_, r_n_191__47_, r_n_191__46_, r_n_191__45_, r_n_191__44_, r_n_191__43_, r_n_191__42_, r_n_191__41_, r_n_191__40_, r_n_191__39_, r_n_191__38_, r_n_191__37_, r_n_191__36_, r_n_191__35_, r_n_191__34_, r_n_191__33_, r_n_191__32_, r_n_191__31_, r_n_191__30_, r_n_191__29_, r_n_191__28_, r_n_191__27_, r_n_191__26_, r_n_191__25_, r_n_191__24_, r_n_191__23_, r_n_191__22_, r_n_191__21_, r_n_191__20_, r_n_191__19_, r_n_191__18_, r_n_191__17_, r_n_191__16_, r_n_191__15_, r_n_191__14_, r_n_191__13_, r_n_191__12_, r_n_191__11_, r_n_191__10_, r_n_191__9_, r_n_191__8_, r_n_191__7_, r_n_191__6_, r_n_191__5_, r_n_191__4_, r_n_191__3_, r_n_191__2_, r_n_191__1_, r_n_191__0_ } = (N382)? { r_192__63_, r_192__62_, r_192__61_, r_192__60_, r_192__59_, r_192__58_, r_192__57_, r_192__56_, r_192__55_, r_192__54_, r_192__53_, r_192__52_, r_192__51_, r_192__50_, r_192__49_, r_192__48_, r_192__47_, r_192__46_, r_192__45_, r_192__44_, r_192__43_, r_192__42_, r_192__41_, r_192__40_, r_192__39_, r_192__38_, r_192__37_, r_192__36_, r_192__35_, r_192__34_, r_192__33_, r_192__32_, r_192__31_, r_192__30_, r_192__29_, r_192__28_, r_192__27_, r_192__26_, r_192__25_, r_192__24_, r_192__23_, r_192__22_, r_192__21_, r_192__20_, r_192__19_, r_192__18_, r_192__17_, r_192__16_, r_192__15_, r_192__14_, r_192__13_, r_192__12_, r_192__11_, r_192__10_, r_192__9_, r_192__8_, r_192__7_, r_192__6_, r_192__5_, r_192__4_, r_192__3_, r_192__2_, r_192__1_, r_192__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N383)? data_i : 1'b0;
  assign N382 = sel_i[382];
  assign N383 = N1983;
  assign { r_n_192__63_, r_n_192__62_, r_n_192__61_, r_n_192__60_, r_n_192__59_, r_n_192__58_, r_n_192__57_, r_n_192__56_, r_n_192__55_, r_n_192__54_, r_n_192__53_, r_n_192__52_, r_n_192__51_, r_n_192__50_, r_n_192__49_, r_n_192__48_, r_n_192__47_, r_n_192__46_, r_n_192__45_, r_n_192__44_, r_n_192__43_, r_n_192__42_, r_n_192__41_, r_n_192__40_, r_n_192__39_, r_n_192__38_, r_n_192__37_, r_n_192__36_, r_n_192__35_, r_n_192__34_, r_n_192__33_, r_n_192__32_, r_n_192__31_, r_n_192__30_, r_n_192__29_, r_n_192__28_, r_n_192__27_, r_n_192__26_, r_n_192__25_, r_n_192__24_, r_n_192__23_, r_n_192__22_, r_n_192__21_, r_n_192__20_, r_n_192__19_, r_n_192__18_, r_n_192__17_, r_n_192__16_, r_n_192__15_, r_n_192__14_, r_n_192__13_, r_n_192__12_, r_n_192__11_, r_n_192__10_, r_n_192__9_, r_n_192__8_, r_n_192__7_, r_n_192__6_, r_n_192__5_, r_n_192__4_, r_n_192__3_, r_n_192__2_, r_n_192__1_, r_n_192__0_ } = (N384)? { r_193__63_, r_193__62_, r_193__61_, r_193__60_, r_193__59_, r_193__58_, r_193__57_, r_193__56_, r_193__55_, r_193__54_, r_193__53_, r_193__52_, r_193__51_, r_193__50_, r_193__49_, r_193__48_, r_193__47_, r_193__46_, r_193__45_, r_193__44_, r_193__43_, r_193__42_, r_193__41_, r_193__40_, r_193__39_, r_193__38_, r_193__37_, r_193__36_, r_193__35_, r_193__34_, r_193__33_, r_193__32_, r_193__31_, r_193__30_, r_193__29_, r_193__28_, r_193__27_, r_193__26_, r_193__25_, r_193__24_, r_193__23_, r_193__22_, r_193__21_, r_193__20_, r_193__19_, r_193__18_, r_193__17_, r_193__16_, r_193__15_, r_193__14_, r_193__13_, r_193__12_, r_193__11_, r_193__10_, r_193__9_, r_193__8_, r_193__7_, r_193__6_, r_193__5_, r_193__4_, r_193__3_, r_193__2_, r_193__1_, r_193__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N385)? data_i : 1'b0;
  assign N384 = sel_i[384];
  assign N385 = N1988;
  assign { r_n_193__63_, r_n_193__62_, r_n_193__61_, r_n_193__60_, r_n_193__59_, r_n_193__58_, r_n_193__57_, r_n_193__56_, r_n_193__55_, r_n_193__54_, r_n_193__53_, r_n_193__52_, r_n_193__51_, r_n_193__50_, r_n_193__49_, r_n_193__48_, r_n_193__47_, r_n_193__46_, r_n_193__45_, r_n_193__44_, r_n_193__43_, r_n_193__42_, r_n_193__41_, r_n_193__40_, r_n_193__39_, r_n_193__38_, r_n_193__37_, r_n_193__36_, r_n_193__35_, r_n_193__34_, r_n_193__33_, r_n_193__32_, r_n_193__31_, r_n_193__30_, r_n_193__29_, r_n_193__28_, r_n_193__27_, r_n_193__26_, r_n_193__25_, r_n_193__24_, r_n_193__23_, r_n_193__22_, r_n_193__21_, r_n_193__20_, r_n_193__19_, r_n_193__18_, r_n_193__17_, r_n_193__16_, r_n_193__15_, r_n_193__14_, r_n_193__13_, r_n_193__12_, r_n_193__11_, r_n_193__10_, r_n_193__9_, r_n_193__8_, r_n_193__7_, r_n_193__6_, r_n_193__5_, r_n_193__4_, r_n_193__3_, r_n_193__2_, r_n_193__1_, r_n_193__0_ } = (N386)? { r_194__63_, r_194__62_, r_194__61_, r_194__60_, r_194__59_, r_194__58_, r_194__57_, r_194__56_, r_194__55_, r_194__54_, r_194__53_, r_194__52_, r_194__51_, r_194__50_, r_194__49_, r_194__48_, r_194__47_, r_194__46_, r_194__45_, r_194__44_, r_194__43_, r_194__42_, r_194__41_, r_194__40_, r_194__39_, r_194__38_, r_194__37_, r_194__36_, r_194__35_, r_194__34_, r_194__33_, r_194__32_, r_194__31_, r_194__30_, r_194__29_, r_194__28_, r_194__27_, r_194__26_, r_194__25_, r_194__24_, r_194__23_, r_194__22_, r_194__21_, r_194__20_, r_194__19_, r_194__18_, r_194__17_, r_194__16_, r_194__15_, r_194__14_, r_194__13_, r_194__12_, r_194__11_, r_194__10_, r_194__9_, r_194__8_, r_194__7_, r_194__6_, r_194__5_, r_194__4_, r_194__3_, r_194__2_, r_194__1_, r_194__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N387)? data_i : 1'b0;
  assign N386 = sel_i[386];
  assign N387 = N1993;
  assign { r_n_194__63_, r_n_194__62_, r_n_194__61_, r_n_194__60_, r_n_194__59_, r_n_194__58_, r_n_194__57_, r_n_194__56_, r_n_194__55_, r_n_194__54_, r_n_194__53_, r_n_194__52_, r_n_194__51_, r_n_194__50_, r_n_194__49_, r_n_194__48_, r_n_194__47_, r_n_194__46_, r_n_194__45_, r_n_194__44_, r_n_194__43_, r_n_194__42_, r_n_194__41_, r_n_194__40_, r_n_194__39_, r_n_194__38_, r_n_194__37_, r_n_194__36_, r_n_194__35_, r_n_194__34_, r_n_194__33_, r_n_194__32_, r_n_194__31_, r_n_194__30_, r_n_194__29_, r_n_194__28_, r_n_194__27_, r_n_194__26_, r_n_194__25_, r_n_194__24_, r_n_194__23_, r_n_194__22_, r_n_194__21_, r_n_194__20_, r_n_194__19_, r_n_194__18_, r_n_194__17_, r_n_194__16_, r_n_194__15_, r_n_194__14_, r_n_194__13_, r_n_194__12_, r_n_194__11_, r_n_194__10_, r_n_194__9_, r_n_194__8_, r_n_194__7_, r_n_194__6_, r_n_194__5_, r_n_194__4_, r_n_194__3_, r_n_194__2_, r_n_194__1_, r_n_194__0_ } = (N388)? { r_195__63_, r_195__62_, r_195__61_, r_195__60_, r_195__59_, r_195__58_, r_195__57_, r_195__56_, r_195__55_, r_195__54_, r_195__53_, r_195__52_, r_195__51_, r_195__50_, r_195__49_, r_195__48_, r_195__47_, r_195__46_, r_195__45_, r_195__44_, r_195__43_, r_195__42_, r_195__41_, r_195__40_, r_195__39_, r_195__38_, r_195__37_, r_195__36_, r_195__35_, r_195__34_, r_195__33_, r_195__32_, r_195__31_, r_195__30_, r_195__29_, r_195__28_, r_195__27_, r_195__26_, r_195__25_, r_195__24_, r_195__23_, r_195__22_, r_195__21_, r_195__20_, r_195__19_, r_195__18_, r_195__17_, r_195__16_, r_195__15_, r_195__14_, r_195__13_, r_195__12_, r_195__11_, r_195__10_, r_195__9_, r_195__8_, r_195__7_, r_195__6_, r_195__5_, r_195__4_, r_195__3_, r_195__2_, r_195__1_, r_195__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N389)? data_i : 1'b0;
  assign N388 = sel_i[388];
  assign N389 = N1998;
  assign { r_n_195__63_, r_n_195__62_, r_n_195__61_, r_n_195__60_, r_n_195__59_, r_n_195__58_, r_n_195__57_, r_n_195__56_, r_n_195__55_, r_n_195__54_, r_n_195__53_, r_n_195__52_, r_n_195__51_, r_n_195__50_, r_n_195__49_, r_n_195__48_, r_n_195__47_, r_n_195__46_, r_n_195__45_, r_n_195__44_, r_n_195__43_, r_n_195__42_, r_n_195__41_, r_n_195__40_, r_n_195__39_, r_n_195__38_, r_n_195__37_, r_n_195__36_, r_n_195__35_, r_n_195__34_, r_n_195__33_, r_n_195__32_, r_n_195__31_, r_n_195__30_, r_n_195__29_, r_n_195__28_, r_n_195__27_, r_n_195__26_, r_n_195__25_, r_n_195__24_, r_n_195__23_, r_n_195__22_, r_n_195__21_, r_n_195__20_, r_n_195__19_, r_n_195__18_, r_n_195__17_, r_n_195__16_, r_n_195__15_, r_n_195__14_, r_n_195__13_, r_n_195__12_, r_n_195__11_, r_n_195__10_, r_n_195__9_, r_n_195__8_, r_n_195__7_, r_n_195__6_, r_n_195__5_, r_n_195__4_, r_n_195__3_, r_n_195__2_, r_n_195__1_, r_n_195__0_ } = (N390)? { r_196__63_, r_196__62_, r_196__61_, r_196__60_, r_196__59_, r_196__58_, r_196__57_, r_196__56_, r_196__55_, r_196__54_, r_196__53_, r_196__52_, r_196__51_, r_196__50_, r_196__49_, r_196__48_, r_196__47_, r_196__46_, r_196__45_, r_196__44_, r_196__43_, r_196__42_, r_196__41_, r_196__40_, r_196__39_, r_196__38_, r_196__37_, r_196__36_, r_196__35_, r_196__34_, r_196__33_, r_196__32_, r_196__31_, r_196__30_, r_196__29_, r_196__28_, r_196__27_, r_196__26_, r_196__25_, r_196__24_, r_196__23_, r_196__22_, r_196__21_, r_196__20_, r_196__19_, r_196__18_, r_196__17_, r_196__16_, r_196__15_, r_196__14_, r_196__13_, r_196__12_, r_196__11_, r_196__10_, r_196__9_, r_196__8_, r_196__7_, r_196__6_, r_196__5_, r_196__4_, r_196__3_, r_196__2_, r_196__1_, r_196__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N391)? data_i : 1'b0;
  assign N390 = sel_i[390];
  assign N391 = N2003;
  assign { r_n_196__63_, r_n_196__62_, r_n_196__61_, r_n_196__60_, r_n_196__59_, r_n_196__58_, r_n_196__57_, r_n_196__56_, r_n_196__55_, r_n_196__54_, r_n_196__53_, r_n_196__52_, r_n_196__51_, r_n_196__50_, r_n_196__49_, r_n_196__48_, r_n_196__47_, r_n_196__46_, r_n_196__45_, r_n_196__44_, r_n_196__43_, r_n_196__42_, r_n_196__41_, r_n_196__40_, r_n_196__39_, r_n_196__38_, r_n_196__37_, r_n_196__36_, r_n_196__35_, r_n_196__34_, r_n_196__33_, r_n_196__32_, r_n_196__31_, r_n_196__30_, r_n_196__29_, r_n_196__28_, r_n_196__27_, r_n_196__26_, r_n_196__25_, r_n_196__24_, r_n_196__23_, r_n_196__22_, r_n_196__21_, r_n_196__20_, r_n_196__19_, r_n_196__18_, r_n_196__17_, r_n_196__16_, r_n_196__15_, r_n_196__14_, r_n_196__13_, r_n_196__12_, r_n_196__11_, r_n_196__10_, r_n_196__9_, r_n_196__8_, r_n_196__7_, r_n_196__6_, r_n_196__5_, r_n_196__4_, r_n_196__3_, r_n_196__2_, r_n_196__1_, r_n_196__0_ } = (N392)? { r_197__63_, r_197__62_, r_197__61_, r_197__60_, r_197__59_, r_197__58_, r_197__57_, r_197__56_, r_197__55_, r_197__54_, r_197__53_, r_197__52_, r_197__51_, r_197__50_, r_197__49_, r_197__48_, r_197__47_, r_197__46_, r_197__45_, r_197__44_, r_197__43_, r_197__42_, r_197__41_, r_197__40_, r_197__39_, r_197__38_, r_197__37_, r_197__36_, r_197__35_, r_197__34_, r_197__33_, r_197__32_, r_197__31_, r_197__30_, r_197__29_, r_197__28_, r_197__27_, r_197__26_, r_197__25_, r_197__24_, r_197__23_, r_197__22_, r_197__21_, r_197__20_, r_197__19_, r_197__18_, r_197__17_, r_197__16_, r_197__15_, r_197__14_, r_197__13_, r_197__12_, r_197__11_, r_197__10_, r_197__9_, r_197__8_, r_197__7_, r_197__6_, r_197__5_, r_197__4_, r_197__3_, r_197__2_, r_197__1_, r_197__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N393)? data_i : 1'b0;
  assign N392 = sel_i[392];
  assign N393 = N2008;
  assign { r_n_197__63_, r_n_197__62_, r_n_197__61_, r_n_197__60_, r_n_197__59_, r_n_197__58_, r_n_197__57_, r_n_197__56_, r_n_197__55_, r_n_197__54_, r_n_197__53_, r_n_197__52_, r_n_197__51_, r_n_197__50_, r_n_197__49_, r_n_197__48_, r_n_197__47_, r_n_197__46_, r_n_197__45_, r_n_197__44_, r_n_197__43_, r_n_197__42_, r_n_197__41_, r_n_197__40_, r_n_197__39_, r_n_197__38_, r_n_197__37_, r_n_197__36_, r_n_197__35_, r_n_197__34_, r_n_197__33_, r_n_197__32_, r_n_197__31_, r_n_197__30_, r_n_197__29_, r_n_197__28_, r_n_197__27_, r_n_197__26_, r_n_197__25_, r_n_197__24_, r_n_197__23_, r_n_197__22_, r_n_197__21_, r_n_197__20_, r_n_197__19_, r_n_197__18_, r_n_197__17_, r_n_197__16_, r_n_197__15_, r_n_197__14_, r_n_197__13_, r_n_197__12_, r_n_197__11_, r_n_197__10_, r_n_197__9_, r_n_197__8_, r_n_197__7_, r_n_197__6_, r_n_197__5_, r_n_197__4_, r_n_197__3_, r_n_197__2_, r_n_197__1_, r_n_197__0_ } = (N394)? { r_198__63_, r_198__62_, r_198__61_, r_198__60_, r_198__59_, r_198__58_, r_198__57_, r_198__56_, r_198__55_, r_198__54_, r_198__53_, r_198__52_, r_198__51_, r_198__50_, r_198__49_, r_198__48_, r_198__47_, r_198__46_, r_198__45_, r_198__44_, r_198__43_, r_198__42_, r_198__41_, r_198__40_, r_198__39_, r_198__38_, r_198__37_, r_198__36_, r_198__35_, r_198__34_, r_198__33_, r_198__32_, r_198__31_, r_198__30_, r_198__29_, r_198__28_, r_198__27_, r_198__26_, r_198__25_, r_198__24_, r_198__23_, r_198__22_, r_198__21_, r_198__20_, r_198__19_, r_198__18_, r_198__17_, r_198__16_, r_198__15_, r_198__14_, r_198__13_, r_198__12_, r_198__11_, r_198__10_, r_198__9_, r_198__8_, r_198__7_, r_198__6_, r_198__5_, r_198__4_, r_198__3_, r_198__2_, r_198__1_, r_198__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N395)? data_i : 1'b0;
  assign N394 = sel_i[394];
  assign N395 = N2013;
  assign { r_n_198__63_, r_n_198__62_, r_n_198__61_, r_n_198__60_, r_n_198__59_, r_n_198__58_, r_n_198__57_, r_n_198__56_, r_n_198__55_, r_n_198__54_, r_n_198__53_, r_n_198__52_, r_n_198__51_, r_n_198__50_, r_n_198__49_, r_n_198__48_, r_n_198__47_, r_n_198__46_, r_n_198__45_, r_n_198__44_, r_n_198__43_, r_n_198__42_, r_n_198__41_, r_n_198__40_, r_n_198__39_, r_n_198__38_, r_n_198__37_, r_n_198__36_, r_n_198__35_, r_n_198__34_, r_n_198__33_, r_n_198__32_, r_n_198__31_, r_n_198__30_, r_n_198__29_, r_n_198__28_, r_n_198__27_, r_n_198__26_, r_n_198__25_, r_n_198__24_, r_n_198__23_, r_n_198__22_, r_n_198__21_, r_n_198__20_, r_n_198__19_, r_n_198__18_, r_n_198__17_, r_n_198__16_, r_n_198__15_, r_n_198__14_, r_n_198__13_, r_n_198__12_, r_n_198__11_, r_n_198__10_, r_n_198__9_, r_n_198__8_, r_n_198__7_, r_n_198__6_, r_n_198__5_, r_n_198__4_, r_n_198__3_, r_n_198__2_, r_n_198__1_, r_n_198__0_ } = (N396)? { r_199__63_, r_199__62_, r_199__61_, r_199__60_, r_199__59_, r_199__58_, r_199__57_, r_199__56_, r_199__55_, r_199__54_, r_199__53_, r_199__52_, r_199__51_, r_199__50_, r_199__49_, r_199__48_, r_199__47_, r_199__46_, r_199__45_, r_199__44_, r_199__43_, r_199__42_, r_199__41_, r_199__40_, r_199__39_, r_199__38_, r_199__37_, r_199__36_, r_199__35_, r_199__34_, r_199__33_, r_199__32_, r_199__31_, r_199__30_, r_199__29_, r_199__28_, r_199__27_, r_199__26_, r_199__25_, r_199__24_, r_199__23_, r_199__22_, r_199__21_, r_199__20_, r_199__19_, r_199__18_, r_199__17_, r_199__16_, r_199__15_, r_199__14_, r_199__13_, r_199__12_, r_199__11_, r_199__10_, r_199__9_, r_199__8_, r_199__7_, r_199__6_, r_199__5_, r_199__4_, r_199__3_, r_199__2_, r_199__1_, r_199__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N397)? data_i : 1'b0;
  assign N396 = sel_i[396];
  assign N397 = N2018;
  assign { r_n_199__63_, r_n_199__62_, r_n_199__61_, r_n_199__60_, r_n_199__59_, r_n_199__58_, r_n_199__57_, r_n_199__56_, r_n_199__55_, r_n_199__54_, r_n_199__53_, r_n_199__52_, r_n_199__51_, r_n_199__50_, r_n_199__49_, r_n_199__48_, r_n_199__47_, r_n_199__46_, r_n_199__45_, r_n_199__44_, r_n_199__43_, r_n_199__42_, r_n_199__41_, r_n_199__40_, r_n_199__39_, r_n_199__38_, r_n_199__37_, r_n_199__36_, r_n_199__35_, r_n_199__34_, r_n_199__33_, r_n_199__32_, r_n_199__31_, r_n_199__30_, r_n_199__29_, r_n_199__28_, r_n_199__27_, r_n_199__26_, r_n_199__25_, r_n_199__24_, r_n_199__23_, r_n_199__22_, r_n_199__21_, r_n_199__20_, r_n_199__19_, r_n_199__18_, r_n_199__17_, r_n_199__16_, r_n_199__15_, r_n_199__14_, r_n_199__13_, r_n_199__12_, r_n_199__11_, r_n_199__10_, r_n_199__9_, r_n_199__8_, r_n_199__7_, r_n_199__6_, r_n_199__5_, r_n_199__4_, r_n_199__3_, r_n_199__2_, r_n_199__1_, r_n_199__0_ } = (N398)? { r_200__63_, r_200__62_, r_200__61_, r_200__60_, r_200__59_, r_200__58_, r_200__57_, r_200__56_, r_200__55_, r_200__54_, r_200__53_, r_200__52_, r_200__51_, r_200__50_, r_200__49_, r_200__48_, r_200__47_, r_200__46_, r_200__45_, r_200__44_, r_200__43_, r_200__42_, r_200__41_, r_200__40_, r_200__39_, r_200__38_, r_200__37_, r_200__36_, r_200__35_, r_200__34_, r_200__33_, r_200__32_, r_200__31_, r_200__30_, r_200__29_, r_200__28_, r_200__27_, r_200__26_, r_200__25_, r_200__24_, r_200__23_, r_200__22_, r_200__21_, r_200__20_, r_200__19_, r_200__18_, r_200__17_, r_200__16_, r_200__15_, r_200__14_, r_200__13_, r_200__12_, r_200__11_, r_200__10_, r_200__9_, r_200__8_, r_200__7_, r_200__6_, r_200__5_, r_200__4_, r_200__3_, r_200__2_, r_200__1_, r_200__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N399)? data_i : 1'b0;
  assign N398 = sel_i[398];
  assign N399 = N2023;
  assign { r_n_200__63_, r_n_200__62_, r_n_200__61_, r_n_200__60_, r_n_200__59_, r_n_200__58_, r_n_200__57_, r_n_200__56_, r_n_200__55_, r_n_200__54_, r_n_200__53_, r_n_200__52_, r_n_200__51_, r_n_200__50_, r_n_200__49_, r_n_200__48_, r_n_200__47_, r_n_200__46_, r_n_200__45_, r_n_200__44_, r_n_200__43_, r_n_200__42_, r_n_200__41_, r_n_200__40_, r_n_200__39_, r_n_200__38_, r_n_200__37_, r_n_200__36_, r_n_200__35_, r_n_200__34_, r_n_200__33_, r_n_200__32_, r_n_200__31_, r_n_200__30_, r_n_200__29_, r_n_200__28_, r_n_200__27_, r_n_200__26_, r_n_200__25_, r_n_200__24_, r_n_200__23_, r_n_200__22_, r_n_200__21_, r_n_200__20_, r_n_200__19_, r_n_200__18_, r_n_200__17_, r_n_200__16_, r_n_200__15_, r_n_200__14_, r_n_200__13_, r_n_200__12_, r_n_200__11_, r_n_200__10_, r_n_200__9_, r_n_200__8_, r_n_200__7_, r_n_200__6_, r_n_200__5_, r_n_200__4_, r_n_200__3_, r_n_200__2_, r_n_200__1_, r_n_200__0_ } = (N400)? { r_201__63_, r_201__62_, r_201__61_, r_201__60_, r_201__59_, r_201__58_, r_201__57_, r_201__56_, r_201__55_, r_201__54_, r_201__53_, r_201__52_, r_201__51_, r_201__50_, r_201__49_, r_201__48_, r_201__47_, r_201__46_, r_201__45_, r_201__44_, r_201__43_, r_201__42_, r_201__41_, r_201__40_, r_201__39_, r_201__38_, r_201__37_, r_201__36_, r_201__35_, r_201__34_, r_201__33_, r_201__32_, r_201__31_, r_201__30_, r_201__29_, r_201__28_, r_201__27_, r_201__26_, r_201__25_, r_201__24_, r_201__23_, r_201__22_, r_201__21_, r_201__20_, r_201__19_, r_201__18_, r_201__17_, r_201__16_, r_201__15_, r_201__14_, r_201__13_, r_201__12_, r_201__11_, r_201__10_, r_201__9_, r_201__8_, r_201__7_, r_201__6_, r_201__5_, r_201__4_, r_201__3_, r_201__2_, r_201__1_, r_201__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N401)? data_i : 1'b0;
  assign N400 = sel_i[400];
  assign N401 = N2028;
  assign { r_n_201__63_, r_n_201__62_, r_n_201__61_, r_n_201__60_, r_n_201__59_, r_n_201__58_, r_n_201__57_, r_n_201__56_, r_n_201__55_, r_n_201__54_, r_n_201__53_, r_n_201__52_, r_n_201__51_, r_n_201__50_, r_n_201__49_, r_n_201__48_, r_n_201__47_, r_n_201__46_, r_n_201__45_, r_n_201__44_, r_n_201__43_, r_n_201__42_, r_n_201__41_, r_n_201__40_, r_n_201__39_, r_n_201__38_, r_n_201__37_, r_n_201__36_, r_n_201__35_, r_n_201__34_, r_n_201__33_, r_n_201__32_, r_n_201__31_, r_n_201__30_, r_n_201__29_, r_n_201__28_, r_n_201__27_, r_n_201__26_, r_n_201__25_, r_n_201__24_, r_n_201__23_, r_n_201__22_, r_n_201__21_, r_n_201__20_, r_n_201__19_, r_n_201__18_, r_n_201__17_, r_n_201__16_, r_n_201__15_, r_n_201__14_, r_n_201__13_, r_n_201__12_, r_n_201__11_, r_n_201__10_, r_n_201__9_, r_n_201__8_, r_n_201__7_, r_n_201__6_, r_n_201__5_, r_n_201__4_, r_n_201__3_, r_n_201__2_, r_n_201__1_, r_n_201__0_ } = (N402)? { r_202__63_, r_202__62_, r_202__61_, r_202__60_, r_202__59_, r_202__58_, r_202__57_, r_202__56_, r_202__55_, r_202__54_, r_202__53_, r_202__52_, r_202__51_, r_202__50_, r_202__49_, r_202__48_, r_202__47_, r_202__46_, r_202__45_, r_202__44_, r_202__43_, r_202__42_, r_202__41_, r_202__40_, r_202__39_, r_202__38_, r_202__37_, r_202__36_, r_202__35_, r_202__34_, r_202__33_, r_202__32_, r_202__31_, r_202__30_, r_202__29_, r_202__28_, r_202__27_, r_202__26_, r_202__25_, r_202__24_, r_202__23_, r_202__22_, r_202__21_, r_202__20_, r_202__19_, r_202__18_, r_202__17_, r_202__16_, r_202__15_, r_202__14_, r_202__13_, r_202__12_, r_202__11_, r_202__10_, r_202__9_, r_202__8_, r_202__7_, r_202__6_, r_202__5_, r_202__4_, r_202__3_, r_202__2_, r_202__1_, r_202__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N403)? data_i : 1'b0;
  assign N402 = sel_i[402];
  assign N403 = N2033;
  assign { r_n_202__63_, r_n_202__62_, r_n_202__61_, r_n_202__60_, r_n_202__59_, r_n_202__58_, r_n_202__57_, r_n_202__56_, r_n_202__55_, r_n_202__54_, r_n_202__53_, r_n_202__52_, r_n_202__51_, r_n_202__50_, r_n_202__49_, r_n_202__48_, r_n_202__47_, r_n_202__46_, r_n_202__45_, r_n_202__44_, r_n_202__43_, r_n_202__42_, r_n_202__41_, r_n_202__40_, r_n_202__39_, r_n_202__38_, r_n_202__37_, r_n_202__36_, r_n_202__35_, r_n_202__34_, r_n_202__33_, r_n_202__32_, r_n_202__31_, r_n_202__30_, r_n_202__29_, r_n_202__28_, r_n_202__27_, r_n_202__26_, r_n_202__25_, r_n_202__24_, r_n_202__23_, r_n_202__22_, r_n_202__21_, r_n_202__20_, r_n_202__19_, r_n_202__18_, r_n_202__17_, r_n_202__16_, r_n_202__15_, r_n_202__14_, r_n_202__13_, r_n_202__12_, r_n_202__11_, r_n_202__10_, r_n_202__9_, r_n_202__8_, r_n_202__7_, r_n_202__6_, r_n_202__5_, r_n_202__4_, r_n_202__3_, r_n_202__2_, r_n_202__1_, r_n_202__0_ } = (N404)? { r_203__63_, r_203__62_, r_203__61_, r_203__60_, r_203__59_, r_203__58_, r_203__57_, r_203__56_, r_203__55_, r_203__54_, r_203__53_, r_203__52_, r_203__51_, r_203__50_, r_203__49_, r_203__48_, r_203__47_, r_203__46_, r_203__45_, r_203__44_, r_203__43_, r_203__42_, r_203__41_, r_203__40_, r_203__39_, r_203__38_, r_203__37_, r_203__36_, r_203__35_, r_203__34_, r_203__33_, r_203__32_, r_203__31_, r_203__30_, r_203__29_, r_203__28_, r_203__27_, r_203__26_, r_203__25_, r_203__24_, r_203__23_, r_203__22_, r_203__21_, r_203__20_, r_203__19_, r_203__18_, r_203__17_, r_203__16_, r_203__15_, r_203__14_, r_203__13_, r_203__12_, r_203__11_, r_203__10_, r_203__9_, r_203__8_, r_203__7_, r_203__6_, r_203__5_, r_203__4_, r_203__3_, r_203__2_, r_203__1_, r_203__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N405)? data_i : 1'b0;
  assign N404 = sel_i[404];
  assign N405 = N2038;
  assign { r_n_203__63_, r_n_203__62_, r_n_203__61_, r_n_203__60_, r_n_203__59_, r_n_203__58_, r_n_203__57_, r_n_203__56_, r_n_203__55_, r_n_203__54_, r_n_203__53_, r_n_203__52_, r_n_203__51_, r_n_203__50_, r_n_203__49_, r_n_203__48_, r_n_203__47_, r_n_203__46_, r_n_203__45_, r_n_203__44_, r_n_203__43_, r_n_203__42_, r_n_203__41_, r_n_203__40_, r_n_203__39_, r_n_203__38_, r_n_203__37_, r_n_203__36_, r_n_203__35_, r_n_203__34_, r_n_203__33_, r_n_203__32_, r_n_203__31_, r_n_203__30_, r_n_203__29_, r_n_203__28_, r_n_203__27_, r_n_203__26_, r_n_203__25_, r_n_203__24_, r_n_203__23_, r_n_203__22_, r_n_203__21_, r_n_203__20_, r_n_203__19_, r_n_203__18_, r_n_203__17_, r_n_203__16_, r_n_203__15_, r_n_203__14_, r_n_203__13_, r_n_203__12_, r_n_203__11_, r_n_203__10_, r_n_203__9_, r_n_203__8_, r_n_203__7_, r_n_203__6_, r_n_203__5_, r_n_203__4_, r_n_203__3_, r_n_203__2_, r_n_203__1_, r_n_203__0_ } = (N406)? { r_204__63_, r_204__62_, r_204__61_, r_204__60_, r_204__59_, r_204__58_, r_204__57_, r_204__56_, r_204__55_, r_204__54_, r_204__53_, r_204__52_, r_204__51_, r_204__50_, r_204__49_, r_204__48_, r_204__47_, r_204__46_, r_204__45_, r_204__44_, r_204__43_, r_204__42_, r_204__41_, r_204__40_, r_204__39_, r_204__38_, r_204__37_, r_204__36_, r_204__35_, r_204__34_, r_204__33_, r_204__32_, r_204__31_, r_204__30_, r_204__29_, r_204__28_, r_204__27_, r_204__26_, r_204__25_, r_204__24_, r_204__23_, r_204__22_, r_204__21_, r_204__20_, r_204__19_, r_204__18_, r_204__17_, r_204__16_, r_204__15_, r_204__14_, r_204__13_, r_204__12_, r_204__11_, r_204__10_, r_204__9_, r_204__8_, r_204__7_, r_204__6_, r_204__5_, r_204__4_, r_204__3_, r_204__2_, r_204__1_, r_204__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N407)? data_i : 1'b0;
  assign N406 = sel_i[406];
  assign N407 = N2043;
  assign { r_n_204__63_, r_n_204__62_, r_n_204__61_, r_n_204__60_, r_n_204__59_, r_n_204__58_, r_n_204__57_, r_n_204__56_, r_n_204__55_, r_n_204__54_, r_n_204__53_, r_n_204__52_, r_n_204__51_, r_n_204__50_, r_n_204__49_, r_n_204__48_, r_n_204__47_, r_n_204__46_, r_n_204__45_, r_n_204__44_, r_n_204__43_, r_n_204__42_, r_n_204__41_, r_n_204__40_, r_n_204__39_, r_n_204__38_, r_n_204__37_, r_n_204__36_, r_n_204__35_, r_n_204__34_, r_n_204__33_, r_n_204__32_, r_n_204__31_, r_n_204__30_, r_n_204__29_, r_n_204__28_, r_n_204__27_, r_n_204__26_, r_n_204__25_, r_n_204__24_, r_n_204__23_, r_n_204__22_, r_n_204__21_, r_n_204__20_, r_n_204__19_, r_n_204__18_, r_n_204__17_, r_n_204__16_, r_n_204__15_, r_n_204__14_, r_n_204__13_, r_n_204__12_, r_n_204__11_, r_n_204__10_, r_n_204__9_, r_n_204__8_, r_n_204__7_, r_n_204__6_, r_n_204__5_, r_n_204__4_, r_n_204__3_, r_n_204__2_, r_n_204__1_, r_n_204__0_ } = (N408)? { r_205__63_, r_205__62_, r_205__61_, r_205__60_, r_205__59_, r_205__58_, r_205__57_, r_205__56_, r_205__55_, r_205__54_, r_205__53_, r_205__52_, r_205__51_, r_205__50_, r_205__49_, r_205__48_, r_205__47_, r_205__46_, r_205__45_, r_205__44_, r_205__43_, r_205__42_, r_205__41_, r_205__40_, r_205__39_, r_205__38_, r_205__37_, r_205__36_, r_205__35_, r_205__34_, r_205__33_, r_205__32_, r_205__31_, r_205__30_, r_205__29_, r_205__28_, r_205__27_, r_205__26_, r_205__25_, r_205__24_, r_205__23_, r_205__22_, r_205__21_, r_205__20_, r_205__19_, r_205__18_, r_205__17_, r_205__16_, r_205__15_, r_205__14_, r_205__13_, r_205__12_, r_205__11_, r_205__10_, r_205__9_, r_205__8_, r_205__7_, r_205__6_, r_205__5_, r_205__4_, r_205__3_, r_205__2_, r_205__1_, r_205__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N409)? data_i : 1'b0;
  assign N408 = sel_i[408];
  assign N409 = N2048;
  assign { r_n_205__63_, r_n_205__62_, r_n_205__61_, r_n_205__60_, r_n_205__59_, r_n_205__58_, r_n_205__57_, r_n_205__56_, r_n_205__55_, r_n_205__54_, r_n_205__53_, r_n_205__52_, r_n_205__51_, r_n_205__50_, r_n_205__49_, r_n_205__48_, r_n_205__47_, r_n_205__46_, r_n_205__45_, r_n_205__44_, r_n_205__43_, r_n_205__42_, r_n_205__41_, r_n_205__40_, r_n_205__39_, r_n_205__38_, r_n_205__37_, r_n_205__36_, r_n_205__35_, r_n_205__34_, r_n_205__33_, r_n_205__32_, r_n_205__31_, r_n_205__30_, r_n_205__29_, r_n_205__28_, r_n_205__27_, r_n_205__26_, r_n_205__25_, r_n_205__24_, r_n_205__23_, r_n_205__22_, r_n_205__21_, r_n_205__20_, r_n_205__19_, r_n_205__18_, r_n_205__17_, r_n_205__16_, r_n_205__15_, r_n_205__14_, r_n_205__13_, r_n_205__12_, r_n_205__11_, r_n_205__10_, r_n_205__9_, r_n_205__8_, r_n_205__7_, r_n_205__6_, r_n_205__5_, r_n_205__4_, r_n_205__3_, r_n_205__2_, r_n_205__1_, r_n_205__0_ } = (N410)? { r_206__63_, r_206__62_, r_206__61_, r_206__60_, r_206__59_, r_206__58_, r_206__57_, r_206__56_, r_206__55_, r_206__54_, r_206__53_, r_206__52_, r_206__51_, r_206__50_, r_206__49_, r_206__48_, r_206__47_, r_206__46_, r_206__45_, r_206__44_, r_206__43_, r_206__42_, r_206__41_, r_206__40_, r_206__39_, r_206__38_, r_206__37_, r_206__36_, r_206__35_, r_206__34_, r_206__33_, r_206__32_, r_206__31_, r_206__30_, r_206__29_, r_206__28_, r_206__27_, r_206__26_, r_206__25_, r_206__24_, r_206__23_, r_206__22_, r_206__21_, r_206__20_, r_206__19_, r_206__18_, r_206__17_, r_206__16_, r_206__15_, r_206__14_, r_206__13_, r_206__12_, r_206__11_, r_206__10_, r_206__9_, r_206__8_, r_206__7_, r_206__6_, r_206__5_, r_206__4_, r_206__3_, r_206__2_, r_206__1_, r_206__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N411)? data_i : 1'b0;
  assign N410 = sel_i[410];
  assign N411 = N2053;
  assign { r_n_206__63_, r_n_206__62_, r_n_206__61_, r_n_206__60_, r_n_206__59_, r_n_206__58_, r_n_206__57_, r_n_206__56_, r_n_206__55_, r_n_206__54_, r_n_206__53_, r_n_206__52_, r_n_206__51_, r_n_206__50_, r_n_206__49_, r_n_206__48_, r_n_206__47_, r_n_206__46_, r_n_206__45_, r_n_206__44_, r_n_206__43_, r_n_206__42_, r_n_206__41_, r_n_206__40_, r_n_206__39_, r_n_206__38_, r_n_206__37_, r_n_206__36_, r_n_206__35_, r_n_206__34_, r_n_206__33_, r_n_206__32_, r_n_206__31_, r_n_206__30_, r_n_206__29_, r_n_206__28_, r_n_206__27_, r_n_206__26_, r_n_206__25_, r_n_206__24_, r_n_206__23_, r_n_206__22_, r_n_206__21_, r_n_206__20_, r_n_206__19_, r_n_206__18_, r_n_206__17_, r_n_206__16_, r_n_206__15_, r_n_206__14_, r_n_206__13_, r_n_206__12_, r_n_206__11_, r_n_206__10_, r_n_206__9_, r_n_206__8_, r_n_206__7_, r_n_206__6_, r_n_206__5_, r_n_206__4_, r_n_206__3_, r_n_206__2_, r_n_206__1_, r_n_206__0_ } = (N412)? { r_207__63_, r_207__62_, r_207__61_, r_207__60_, r_207__59_, r_207__58_, r_207__57_, r_207__56_, r_207__55_, r_207__54_, r_207__53_, r_207__52_, r_207__51_, r_207__50_, r_207__49_, r_207__48_, r_207__47_, r_207__46_, r_207__45_, r_207__44_, r_207__43_, r_207__42_, r_207__41_, r_207__40_, r_207__39_, r_207__38_, r_207__37_, r_207__36_, r_207__35_, r_207__34_, r_207__33_, r_207__32_, r_207__31_, r_207__30_, r_207__29_, r_207__28_, r_207__27_, r_207__26_, r_207__25_, r_207__24_, r_207__23_, r_207__22_, r_207__21_, r_207__20_, r_207__19_, r_207__18_, r_207__17_, r_207__16_, r_207__15_, r_207__14_, r_207__13_, r_207__12_, r_207__11_, r_207__10_, r_207__9_, r_207__8_, r_207__7_, r_207__6_, r_207__5_, r_207__4_, r_207__3_, r_207__2_, r_207__1_, r_207__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N413)? data_i : 1'b0;
  assign N412 = sel_i[412];
  assign N413 = N2058;
  assign { r_n_207__63_, r_n_207__62_, r_n_207__61_, r_n_207__60_, r_n_207__59_, r_n_207__58_, r_n_207__57_, r_n_207__56_, r_n_207__55_, r_n_207__54_, r_n_207__53_, r_n_207__52_, r_n_207__51_, r_n_207__50_, r_n_207__49_, r_n_207__48_, r_n_207__47_, r_n_207__46_, r_n_207__45_, r_n_207__44_, r_n_207__43_, r_n_207__42_, r_n_207__41_, r_n_207__40_, r_n_207__39_, r_n_207__38_, r_n_207__37_, r_n_207__36_, r_n_207__35_, r_n_207__34_, r_n_207__33_, r_n_207__32_, r_n_207__31_, r_n_207__30_, r_n_207__29_, r_n_207__28_, r_n_207__27_, r_n_207__26_, r_n_207__25_, r_n_207__24_, r_n_207__23_, r_n_207__22_, r_n_207__21_, r_n_207__20_, r_n_207__19_, r_n_207__18_, r_n_207__17_, r_n_207__16_, r_n_207__15_, r_n_207__14_, r_n_207__13_, r_n_207__12_, r_n_207__11_, r_n_207__10_, r_n_207__9_, r_n_207__8_, r_n_207__7_, r_n_207__6_, r_n_207__5_, r_n_207__4_, r_n_207__3_, r_n_207__2_, r_n_207__1_, r_n_207__0_ } = (N414)? { r_208__63_, r_208__62_, r_208__61_, r_208__60_, r_208__59_, r_208__58_, r_208__57_, r_208__56_, r_208__55_, r_208__54_, r_208__53_, r_208__52_, r_208__51_, r_208__50_, r_208__49_, r_208__48_, r_208__47_, r_208__46_, r_208__45_, r_208__44_, r_208__43_, r_208__42_, r_208__41_, r_208__40_, r_208__39_, r_208__38_, r_208__37_, r_208__36_, r_208__35_, r_208__34_, r_208__33_, r_208__32_, r_208__31_, r_208__30_, r_208__29_, r_208__28_, r_208__27_, r_208__26_, r_208__25_, r_208__24_, r_208__23_, r_208__22_, r_208__21_, r_208__20_, r_208__19_, r_208__18_, r_208__17_, r_208__16_, r_208__15_, r_208__14_, r_208__13_, r_208__12_, r_208__11_, r_208__10_, r_208__9_, r_208__8_, r_208__7_, r_208__6_, r_208__5_, r_208__4_, r_208__3_, r_208__2_, r_208__1_, r_208__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N415)? data_i : 1'b0;
  assign N414 = sel_i[414];
  assign N415 = N2063;
  assign { r_n_208__63_, r_n_208__62_, r_n_208__61_, r_n_208__60_, r_n_208__59_, r_n_208__58_, r_n_208__57_, r_n_208__56_, r_n_208__55_, r_n_208__54_, r_n_208__53_, r_n_208__52_, r_n_208__51_, r_n_208__50_, r_n_208__49_, r_n_208__48_, r_n_208__47_, r_n_208__46_, r_n_208__45_, r_n_208__44_, r_n_208__43_, r_n_208__42_, r_n_208__41_, r_n_208__40_, r_n_208__39_, r_n_208__38_, r_n_208__37_, r_n_208__36_, r_n_208__35_, r_n_208__34_, r_n_208__33_, r_n_208__32_, r_n_208__31_, r_n_208__30_, r_n_208__29_, r_n_208__28_, r_n_208__27_, r_n_208__26_, r_n_208__25_, r_n_208__24_, r_n_208__23_, r_n_208__22_, r_n_208__21_, r_n_208__20_, r_n_208__19_, r_n_208__18_, r_n_208__17_, r_n_208__16_, r_n_208__15_, r_n_208__14_, r_n_208__13_, r_n_208__12_, r_n_208__11_, r_n_208__10_, r_n_208__9_, r_n_208__8_, r_n_208__7_, r_n_208__6_, r_n_208__5_, r_n_208__4_, r_n_208__3_, r_n_208__2_, r_n_208__1_, r_n_208__0_ } = (N416)? { r_209__63_, r_209__62_, r_209__61_, r_209__60_, r_209__59_, r_209__58_, r_209__57_, r_209__56_, r_209__55_, r_209__54_, r_209__53_, r_209__52_, r_209__51_, r_209__50_, r_209__49_, r_209__48_, r_209__47_, r_209__46_, r_209__45_, r_209__44_, r_209__43_, r_209__42_, r_209__41_, r_209__40_, r_209__39_, r_209__38_, r_209__37_, r_209__36_, r_209__35_, r_209__34_, r_209__33_, r_209__32_, r_209__31_, r_209__30_, r_209__29_, r_209__28_, r_209__27_, r_209__26_, r_209__25_, r_209__24_, r_209__23_, r_209__22_, r_209__21_, r_209__20_, r_209__19_, r_209__18_, r_209__17_, r_209__16_, r_209__15_, r_209__14_, r_209__13_, r_209__12_, r_209__11_, r_209__10_, r_209__9_, r_209__8_, r_209__7_, r_209__6_, r_209__5_, r_209__4_, r_209__3_, r_209__2_, r_209__1_, r_209__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N417)? data_i : 1'b0;
  assign N416 = sel_i[416];
  assign N417 = N2068;
  assign { r_n_209__63_, r_n_209__62_, r_n_209__61_, r_n_209__60_, r_n_209__59_, r_n_209__58_, r_n_209__57_, r_n_209__56_, r_n_209__55_, r_n_209__54_, r_n_209__53_, r_n_209__52_, r_n_209__51_, r_n_209__50_, r_n_209__49_, r_n_209__48_, r_n_209__47_, r_n_209__46_, r_n_209__45_, r_n_209__44_, r_n_209__43_, r_n_209__42_, r_n_209__41_, r_n_209__40_, r_n_209__39_, r_n_209__38_, r_n_209__37_, r_n_209__36_, r_n_209__35_, r_n_209__34_, r_n_209__33_, r_n_209__32_, r_n_209__31_, r_n_209__30_, r_n_209__29_, r_n_209__28_, r_n_209__27_, r_n_209__26_, r_n_209__25_, r_n_209__24_, r_n_209__23_, r_n_209__22_, r_n_209__21_, r_n_209__20_, r_n_209__19_, r_n_209__18_, r_n_209__17_, r_n_209__16_, r_n_209__15_, r_n_209__14_, r_n_209__13_, r_n_209__12_, r_n_209__11_, r_n_209__10_, r_n_209__9_, r_n_209__8_, r_n_209__7_, r_n_209__6_, r_n_209__5_, r_n_209__4_, r_n_209__3_, r_n_209__2_, r_n_209__1_, r_n_209__0_ } = (N418)? { r_210__63_, r_210__62_, r_210__61_, r_210__60_, r_210__59_, r_210__58_, r_210__57_, r_210__56_, r_210__55_, r_210__54_, r_210__53_, r_210__52_, r_210__51_, r_210__50_, r_210__49_, r_210__48_, r_210__47_, r_210__46_, r_210__45_, r_210__44_, r_210__43_, r_210__42_, r_210__41_, r_210__40_, r_210__39_, r_210__38_, r_210__37_, r_210__36_, r_210__35_, r_210__34_, r_210__33_, r_210__32_, r_210__31_, r_210__30_, r_210__29_, r_210__28_, r_210__27_, r_210__26_, r_210__25_, r_210__24_, r_210__23_, r_210__22_, r_210__21_, r_210__20_, r_210__19_, r_210__18_, r_210__17_, r_210__16_, r_210__15_, r_210__14_, r_210__13_, r_210__12_, r_210__11_, r_210__10_, r_210__9_, r_210__8_, r_210__7_, r_210__6_, r_210__5_, r_210__4_, r_210__3_, r_210__2_, r_210__1_, r_210__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N419)? data_i : 1'b0;
  assign N418 = sel_i[418];
  assign N419 = N2073;
  assign { r_n_210__63_, r_n_210__62_, r_n_210__61_, r_n_210__60_, r_n_210__59_, r_n_210__58_, r_n_210__57_, r_n_210__56_, r_n_210__55_, r_n_210__54_, r_n_210__53_, r_n_210__52_, r_n_210__51_, r_n_210__50_, r_n_210__49_, r_n_210__48_, r_n_210__47_, r_n_210__46_, r_n_210__45_, r_n_210__44_, r_n_210__43_, r_n_210__42_, r_n_210__41_, r_n_210__40_, r_n_210__39_, r_n_210__38_, r_n_210__37_, r_n_210__36_, r_n_210__35_, r_n_210__34_, r_n_210__33_, r_n_210__32_, r_n_210__31_, r_n_210__30_, r_n_210__29_, r_n_210__28_, r_n_210__27_, r_n_210__26_, r_n_210__25_, r_n_210__24_, r_n_210__23_, r_n_210__22_, r_n_210__21_, r_n_210__20_, r_n_210__19_, r_n_210__18_, r_n_210__17_, r_n_210__16_, r_n_210__15_, r_n_210__14_, r_n_210__13_, r_n_210__12_, r_n_210__11_, r_n_210__10_, r_n_210__9_, r_n_210__8_, r_n_210__7_, r_n_210__6_, r_n_210__5_, r_n_210__4_, r_n_210__3_, r_n_210__2_, r_n_210__1_, r_n_210__0_ } = (N420)? { r_211__63_, r_211__62_, r_211__61_, r_211__60_, r_211__59_, r_211__58_, r_211__57_, r_211__56_, r_211__55_, r_211__54_, r_211__53_, r_211__52_, r_211__51_, r_211__50_, r_211__49_, r_211__48_, r_211__47_, r_211__46_, r_211__45_, r_211__44_, r_211__43_, r_211__42_, r_211__41_, r_211__40_, r_211__39_, r_211__38_, r_211__37_, r_211__36_, r_211__35_, r_211__34_, r_211__33_, r_211__32_, r_211__31_, r_211__30_, r_211__29_, r_211__28_, r_211__27_, r_211__26_, r_211__25_, r_211__24_, r_211__23_, r_211__22_, r_211__21_, r_211__20_, r_211__19_, r_211__18_, r_211__17_, r_211__16_, r_211__15_, r_211__14_, r_211__13_, r_211__12_, r_211__11_, r_211__10_, r_211__9_, r_211__8_, r_211__7_, r_211__6_, r_211__5_, r_211__4_, r_211__3_, r_211__2_, r_211__1_, r_211__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N421)? data_i : 1'b0;
  assign N420 = sel_i[420];
  assign N421 = N2078;
  assign { r_n_211__63_, r_n_211__62_, r_n_211__61_, r_n_211__60_, r_n_211__59_, r_n_211__58_, r_n_211__57_, r_n_211__56_, r_n_211__55_, r_n_211__54_, r_n_211__53_, r_n_211__52_, r_n_211__51_, r_n_211__50_, r_n_211__49_, r_n_211__48_, r_n_211__47_, r_n_211__46_, r_n_211__45_, r_n_211__44_, r_n_211__43_, r_n_211__42_, r_n_211__41_, r_n_211__40_, r_n_211__39_, r_n_211__38_, r_n_211__37_, r_n_211__36_, r_n_211__35_, r_n_211__34_, r_n_211__33_, r_n_211__32_, r_n_211__31_, r_n_211__30_, r_n_211__29_, r_n_211__28_, r_n_211__27_, r_n_211__26_, r_n_211__25_, r_n_211__24_, r_n_211__23_, r_n_211__22_, r_n_211__21_, r_n_211__20_, r_n_211__19_, r_n_211__18_, r_n_211__17_, r_n_211__16_, r_n_211__15_, r_n_211__14_, r_n_211__13_, r_n_211__12_, r_n_211__11_, r_n_211__10_, r_n_211__9_, r_n_211__8_, r_n_211__7_, r_n_211__6_, r_n_211__5_, r_n_211__4_, r_n_211__3_, r_n_211__2_, r_n_211__1_, r_n_211__0_ } = (N422)? { r_212__63_, r_212__62_, r_212__61_, r_212__60_, r_212__59_, r_212__58_, r_212__57_, r_212__56_, r_212__55_, r_212__54_, r_212__53_, r_212__52_, r_212__51_, r_212__50_, r_212__49_, r_212__48_, r_212__47_, r_212__46_, r_212__45_, r_212__44_, r_212__43_, r_212__42_, r_212__41_, r_212__40_, r_212__39_, r_212__38_, r_212__37_, r_212__36_, r_212__35_, r_212__34_, r_212__33_, r_212__32_, r_212__31_, r_212__30_, r_212__29_, r_212__28_, r_212__27_, r_212__26_, r_212__25_, r_212__24_, r_212__23_, r_212__22_, r_212__21_, r_212__20_, r_212__19_, r_212__18_, r_212__17_, r_212__16_, r_212__15_, r_212__14_, r_212__13_, r_212__12_, r_212__11_, r_212__10_, r_212__9_, r_212__8_, r_212__7_, r_212__6_, r_212__5_, r_212__4_, r_212__3_, r_212__2_, r_212__1_, r_212__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N423)? data_i : 1'b0;
  assign N422 = sel_i[422];
  assign N423 = N2083;
  assign { r_n_212__63_, r_n_212__62_, r_n_212__61_, r_n_212__60_, r_n_212__59_, r_n_212__58_, r_n_212__57_, r_n_212__56_, r_n_212__55_, r_n_212__54_, r_n_212__53_, r_n_212__52_, r_n_212__51_, r_n_212__50_, r_n_212__49_, r_n_212__48_, r_n_212__47_, r_n_212__46_, r_n_212__45_, r_n_212__44_, r_n_212__43_, r_n_212__42_, r_n_212__41_, r_n_212__40_, r_n_212__39_, r_n_212__38_, r_n_212__37_, r_n_212__36_, r_n_212__35_, r_n_212__34_, r_n_212__33_, r_n_212__32_, r_n_212__31_, r_n_212__30_, r_n_212__29_, r_n_212__28_, r_n_212__27_, r_n_212__26_, r_n_212__25_, r_n_212__24_, r_n_212__23_, r_n_212__22_, r_n_212__21_, r_n_212__20_, r_n_212__19_, r_n_212__18_, r_n_212__17_, r_n_212__16_, r_n_212__15_, r_n_212__14_, r_n_212__13_, r_n_212__12_, r_n_212__11_, r_n_212__10_, r_n_212__9_, r_n_212__8_, r_n_212__7_, r_n_212__6_, r_n_212__5_, r_n_212__4_, r_n_212__3_, r_n_212__2_, r_n_212__1_, r_n_212__0_ } = (N424)? { r_213__63_, r_213__62_, r_213__61_, r_213__60_, r_213__59_, r_213__58_, r_213__57_, r_213__56_, r_213__55_, r_213__54_, r_213__53_, r_213__52_, r_213__51_, r_213__50_, r_213__49_, r_213__48_, r_213__47_, r_213__46_, r_213__45_, r_213__44_, r_213__43_, r_213__42_, r_213__41_, r_213__40_, r_213__39_, r_213__38_, r_213__37_, r_213__36_, r_213__35_, r_213__34_, r_213__33_, r_213__32_, r_213__31_, r_213__30_, r_213__29_, r_213__28_, r_213__27_, r_213__26_, r_213__25_, r_213__24_, r_213__23_, r_213__22_, r_213__21_, r_213__20_, r_213__19_, r_213__18_, r_213__17_, r_213__16_, r_213__15_, r_213__14_, r_213__13_, r_213__12_, r_213__11_, r_213__10_, r_213__9_, r_213__8_, r_213__7_, r_213__6_, r_213__5_, r_213__4_, r_213__3_, r_213__2_, r_213__1_, r_213__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N425)? data_i : 1'b0;
  assign N424 = sel_i[424];
  assign N425 = N2088;
  assign { r_n_213__63_, r_n_213__62_, r_n_213__61_, r_n_213__60_, r_n_213__59_, r_n_213__58_, r_n_213__57_, r_n_213__56_, r_n_213__55_, r_n_213__54_, r_n_213__53_, r_n_213__52_, r_n_213__51_, r_n_213__50_, r_n_213__49_, r_n_213__48_, r_n_213__47_, r_n_213__46_, r_n_213__45_, r_n_213__44_, r_n_213__43_, r_n_213__42_, r_n_213__41_, r_n_213__40_, r_n_213__39_, r_n_213__38_, r_n_213__37_, r_n_213__36_, r_n_213__35_, r_n_213__34_, r_n_213__33_, r_n_213__32_, r_n_213__31_, r_n_213__30_, r_n_213__29_, r_n_213__28_, r_n_213__27_, r_n_213__26_, r_n_213__25_, r_n_213__24_, r_n_213__23_, r_n_213__22_, r_n_213__21_, r_n_213__20_, r_n_213__19_, r_n_213__18_, r_n_213__17_, r_n_213__16_, r_n_213__15_, r_n_213__14_, r_n_213__13_, r_n_213__12_, r_n_213__11_, r_n_213__10_, r_n_213__9_, r_n_213__8_, r_n_213__7_, r_n_213__6_, r_n_213__5_, r_n_213__4_, r_n_213__3_, r_n_213__2_, r_n_213__1_, r_n_213__0_ } = (N426)? { r_214__63_, r_214__62_, r_214__61_, r_214__60_, r_214__59_, r_214__58_, r_214__57_, r_214__56_, r_214__55_, r_214__54_, r_214__53_, r_214__52_, r_214__51_, r_214__50_, r_214__49_, r_214__48_, r_214__47_, r_214__46_, r_214__45_, r_214__44_, r_214__43_, r_214__42_, r_214__41_, r_214__40_, r_214__39_, r_214__38_, r_214__37_, r_214__36_, r_214__35_, r_214__34_, r_214__33_, r_214__32_, r_214__31_, r_214__30_, r_214__29_, r_214__28_, r_214__27_, r_214__26_, r_214__25_, r_214__24_, r_214__23_, r_214__22_, r_214__21_, r_214__20_, r_214__19_, r_214__18_, r_214__17_, r_214__16_, r_214__15_, r_214__14_, r_214__13_, r_214__12_, r_214__11_, r_214__10_, r_214__9_, r_214__8_, r_214__7_, r_214__6_, r_214__5_, r_214__4_, r_214__3_, r_214__2_, r_214__1_, r_214__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N427)? data_i : 1'b0;
  assign N426 = sel_i[426];
  assign N427 = N2093;
  assign { r_n_214__63_, r_n_214__62_, r_n_214__61_, r_n_214__60_, r_n_214__59_, r_n_214__58_, r_n_214__57_, r_n_214__56_, r_n_214__55_, r_n_214__54_, r_n_214__53_, r_n_214__52_, r_n_214__51_, r_n_214__50_, r_n_214__49_, r_n_214__48_, r_n_214__47_, r_n_214__46_, r_n_214__45_, r_n_214__44_, r_n_214__43_, r_n_214__42_, r_n_214__41_, r_n_214__40_, r_n_214__39_, r_n_214__38_, r_n_214__37_, r_n_214__36_, r_n_214__35_, r_n_214__34_, r_n_214__33_, r_n_214__32_, r_n_214__31_, r_n_214__30_, r_n_214__29_, r_n_214__28_, r_n_214__27_, r_n_214__26_, r_n_214__25_, r_n_214__24_, r_n_214__23_, r_n_214__22_, r_n_214__21_, r_n_214__20_, r_n_214__19_, r_n_214__18_, r_n_214__17_, r_n_214__16_, r_n_214__15_, r_n_214__14_, r_n_214__13_, r_n_214__12_, r_n_214__11_, r_n_214__10_, r_n_214__9_, r_n_214__8_, r_n_214__7_, r_n_214__6_, r_n_214__5_, r_n_214__4_, r_n_214__3_, r_n_214__2_, r_n_214__1_, r_n_214__0_ } = (N428)? { r_215__63_, r_215__62_, r_215__61_, r_215__60_, r_215__59_, r_215__58_, r_215__57_, r_215__56_, r_215__55_, r_215__54_, r_215__53_, r_215__52_, r_215__51_, r_215__50_, r_215__49_, r_215__48_, r_215__47_, r_215__46_, r_215__45_, r_215__44_, r_215__43_, r_215__42_, r_215__41_, r_215__40_, r_215__39_, r_215__38_, r_215__37_, r_215__36_, r_215__35_, r_215__34_, r_215__33_, r_215__32_, r_215__31_, r_215__30_, r_215__29_, r_215__28_, r_215__27_, r_215__26_, r_215__25_, r_215__24_, r_215__23_, r_215__22_, r_215__21_, r_215__20_, r_215__19_, r_215__18_, r_215__17_, r_215__16_, r_215__15_, r_215__14_, r_215__13_, r_215__12_, r_215__11_, r_215__10_, r_215__9_, r_215__8_, r_215__7_, r_215__6_, r_215__5_, r_215__4_, r_215__3_, r_215__2_, r_215__1_, r_215__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N429)? data_i : 1'b0;
  assign N428 = sel_i[428];
  assign N429 = N2098;
  assign { r_n_215__63_, r_n_215__62_, r_n_215__61_, r_n_215__60_, r_n_215__59_, r_n_215__58_, r_n_215__57_, r_n_215__56_, r_n_215__55_, r_n_215__54_, r_n_215__53_, r_n_215__52_, r_n_215__51_, r_n_215__50_, r_n_215__49_, r_n_215__48_, r_n_215__47_, r_n_215__46_, r_n_215__45_, r_n_215__44_, r_n_215__43_, r_n_215__42_, r_n_215__41_, r_n_215__40_, r_n_215__39_, r_n_215__38_, r_n_215__37_, r_n_215__36_, r_n_215__35_, r_n_215__34_, r_n_215__33_, r_n_215__32_, r_n_215__31_, r_n_215__30_, r_n_215__29_, r_n_215__28_, r_n_215__27_, r_n_215__26_, r_n_215__25_, r_n_215__24_, r_n_215__23_, r_n_215__22_, r_n_215__21_, r_n_215__20_, r_n_215__19_, r_n_215__18_, r_n_215__17_, r_n_215__16_, r_n_215__15_, r_n_215__14_, r_n_215__13_, r_n_215__12_, r_n_215__11_, r_n_215__10_, r_n_215__9_, r_n_215__8_, r_n_215__7_, r_n_215__6_, r_n_215__5_, r_n_215__4_, r_n_215__3_, r_n_215__2_, r_n_215__1_, r_n_215__0_ } = (N430)? { r_216__63_, r_216__62_, r_216__61_, r_216__60_, r_216__59_, r_216__58_, r_216__57_, r_216__56_, r_216__55_, r_216__54_, r_216__53_, r_216__52_, r_216__51_, r_216__50_, r_216__49_, r_216__48_, r_216__47_, r_216__46_, r_216__45_, r_216__44_, r_216__43_, r_216__42_, r_216__41_, r_216__40_, r_216__39_, r_216__38_, r_216__37_, r_216__36_, r_216__35_, r_216__34_, r_216__33_, r_216__32_, r_216__31_, r_216__30_, r_216__29_, r_216__28_, r_216__27_, r_216__26_, r_216__25_, r_216__24_, r_216__23_, r_216__22_, r_216__21_, r_216__20_, r_216__19_, r_216__18_, r_216__17_, r_216__16_, r_216__15_, r_216__14_, r_216__13_, r_216__12_, r_216__11_, r_216__10_, r_216__9_, r_216__8_, r_216__7_, r_216__6_, r_216__5_, r_216__4_, r_216__3_, r_216__2_, r_216__1_, r_216__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N431)? data_i : 1'b0;
  assign N430 = sel_i[430];
  assign N431 = N2103;
  assign { r_n_216__63_, r_n_216__62_, r_n_216__61_, r_n_216__60_, r_n_216__59_, r_n_216__58_, r_n_216__57_, r_n_216__56_, r_n_216__55_, r_n_216__54_, r_n_216__53_, r_n_216__52_, r_n_216__51_, r_n_216__50_, r_n_216__49_, r_n_216__48_, r_n_216__47_, r_n_216__46_, r_n_216__45_, r_n_216__44_, r_n_216__43_, r_n_216__42_, r_n_216__41_, r_n_216__40_, r_n_216__39_, r_n_216__38_, r_n_216__37_, r_n_216__36_, r_n_216__35_, r_n_216__34_, r_n_216__33_, r_n_216__32_, r_n_216__31_, r_n_216__30_, r_n_216__29_, r_n_216__28_, r_n_216__27_, r_n_216__26_, r_n_216__25_, r_n_216__24_, r_n_216__23_, r_n_216__22_, r_n_216__21_, r_n_216__20_, r_n_216__19_, r_n_216__18_, r_n_216__17_, r_n_216__16_, r_n_216__15_, r_n_216__14_, r_n_216__13_, r_n_216__12_, r_n_216__11_, r_n_216__10_, r_n_216__9_, r_n_216__8_, r_n_216__7_, r_n_216__6_, r_n_216__5_, r_n_216__4_, r_n_216__3_, r_n_216__2_, r_n_216__1_, r_n_216__0_ } = (N432)? { r_217__63_, r_217__62_, r_217__61_, r_217__60_, r_217__59_, r_217__58_, r_217__57_, r_217__56_, r_217__55_, r_217__54_, r_217__53_, r_217__52_, r_217__51_, r_217__50_, r_217__49_, r_217__48_, r_217__47_, r_217__46_, r_217__45_, r_217__44_, r_217__43_, r_217__42_, r_217__41_, r_217__40_, r_217__39_, r_217__38_, r_217__37_, r_217__36_, r_217__35_, r_217__34_, r_217__33_, r_217__32_, r_217__31_, r_217__30_, r_217__29_, r_217__28_, r_217__27_, r_217__26_, r_217__25_, r_217__24_, r_217__23_, r_217__22_, r_217__21_, r_217__20_, r_217__19_, r_217__18_, r_217__17_, r_217__16_, r_217__15_, r_217__14_, r_217__13_, r_217__12_, r_217__11_, r_217__10_, r_217__9_, r_217__8_, r_217__7_, r_217__6_, r_217__5_, r_217__4_, r_217__3_, r_217__2_, r_217__1_, r_217__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N433)? data_i : 1'b0;
  assign N432 = sel_i[432];
  assign N433 = N2108;
  assign { r_n_217__63_, r_n_217__62_, r_n_217__61_, r_n_217__60_, r_n_217__59_, r_n_217__58_, r_n_217__57_, r_n_217__56_, r_n_217__55_, r_n_217__54_, r_n_217__53_, r_n_217__52_, r_n_217__51_, r_n_217__50_, r_n_217__49_, r_n_217__48_, r_n_217__47_, r_n_217__46_, r_n_217__45_, r_n_217__44_, r_n_217__43_, r_n_217__42_, r_n_217__41_, r_n_217__40_, r_n_217__39_, r_n_217__38_, r_n_217__37_, r_n_217__36_, r_n_217__35_, r_n_217__34_, r_n_217__33_, r_n_217__32_, r_n_217__31_, r_n_217__30_, r_n_217__29_, r_n_217__28_, r_n_217__27_, r_n_217__26_, r_n_217__25_, r_n_217__24_, r_n_217__23_, r_n_217__22_, r_n_217__21_, r_n_217__20_, r_n_217__19_, r_n_217__18_, r_n_217__17_, r_n_217__16_, r_n_217__15_, r_n_217__14_, r_n_217__13_, r_n_217__12_, r_n_217__11_, r_n_217__10_, r_n_217__9_, r_n_217__8_, r_n_217__7_, r_n_217__6_, r_n_217__5_, r_n_217__4_, r_n_217__3_, r_n_217__2_, r_n_217__1_, r_n_217__0_ } = (N434)? { r_218__63_, r_218__62_, r_218__61_, r_218__60_, r_218__59_, r_218__58_, r_218__57_, r_218__56_, r_218__55_, r_218__54_, r_218__53_, r_218__52_, r_218__51_, r_218__50_, r_218__49_, r_218__48_, r_218__47_, r_218__46_, r_218__45_, r_218__44_, r_218__43_, r_218__42_, r_218__41_, r_218__40_, r_218__39_, r_218__38_, r_218__37_, r_218__36_, r_218__35_, r_218__34_, r_218__33_, r_218__32_, r_218__31_, r_218__30_, r_218__29_, r_218__28_, r_218__27_, r_218__26_, r_218__25_, r_218__24_, r_218__23_, r_218__22_, r_218__21_, r_218__20_, r_218__19_, r_218__18_, r_218__17_, r_218__16_, r_218__15_, r_218__14_, r_218__13_, r_218__12_, r_218__11_, r_218__10_, r_218__9_, r_218__8_, r_218__7_, r_218__6_, r_218__5_, r_218__4_, r_218__3_, r_218__2_, r_218__1_, r_218__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N435)? data_i : 1'b0;
  assign N434 = sel_i[434];
  assign N435 = N2113;
  assign { r_n_218__63_, r_n_218__62_, r_n_218__61_, r_n_218__60_, r_n_218__59_, r_n_218__58_, r_n_218__57_, r_n_218__56_, r_n_218__55_, r_n_218__54_, r_n_218__53_, r_n_218__52_, r_n_218__51_, r_n_218__50_, r_n_218__49_, r_n_218__48_, r_n_218__47_, r_n_218__46_, r_n_218__45_, r_n_218__44_, r_n_218__43_, r_n_218__42_, r_n_218__41_, r_n_218__40_, r_n_218__39_, r_n_218__38_, r_n_218__37_, r_n_218__36_, r_n_218__35_, r_n_218__34_, r_n_218__33_, r_n_218__32_, r_n_218__31_, r_n_218__30_, r_n_218__29_, r_n_218__28_, r_n_218__27_, r_n_218__26_, r_n_218__25_, r_n_218__24_, r_n_218__23_, r_n_218__22_, r_n_218__21_, r_n_218__20_, r_n_218__19_, r_n_218__18_, r_n_218__17_, r_n_218__16_, r_n_218__15_, r_n_218__14_, r_n_218__13_, r_n_218__12_, r_n_218__11_, r_n_218__10_, r_n_218__9_, r_n_218__8_, r_n_218__7_, r_n_218__6_, r_n_218__5_, r_n_218__4_, r_n_218__3_, r_n_218__2_, r_n_218__1_, r_n_218__0_ } = (N436)? { r_219__63_, r_219__62_, r_219__61_, r_219__60_, r_219__59_, r_219__58_, r_219__57_, r_219__56_, r_219__55_, r_219__54_, r_219__53_, r_219__52_, r_219__51_, r_219__50_, r_219__49_, r_219__48_, r_219__47_, r_219__46_, r_219__45_, r_219__44_, r_219__43_, r_219__42_, r_219__41_, r_219__40_, r_219__39_, r_219__38_, r_219__37_, r_219__36_, r_219__35_, r_219__34_, r_219__33_, r_219__32_, r_219__31_, r_219__30_, r_219__29_, r_219__28_, r_219__27_, r_219__26_, r_219__25_, r_219__24_, r_219__23_, r_219__22_, r_219__21_, r_219__20_, r_219__19_, r_219__18_, r_219__17_, r_219__16_, r_219__15_, r_219__14_, r_219__13_, r_219__12_, r_219__11_, r_219__10_, r_219__9_, r_219__8_, r_219__7_, r_219__6_, r_219__5_, r_219__4_, r_219__3_, r_219__2_, r_219__1_, r_219__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N437)? data_i : 1'b0;
  assign N436 = sel_i[436];
  assign N437 = N2118;
  assign { r_n_219__63_, r_n_219__62_, r_n_219__61_, r_n_219__60_, r_n_219__59_, r_n_219__58_, r_n_219__57_, r_n_219__56_, r_n_219__55_, r_n_219__54_, r_n_219__53_, r_n_219__52_, r_n_219__51_, r_n_219__50_, r_n_219__49_, r_n_219__48_, r_n_219__47_, r_n_219__46_, r_n_219__45_, r_n_219__44_, r_n_219__43_, r_n_219__42_, r_n_219__41_, r_n_219__40_, r_n_219__39_, r_n_219__38_, r_n_219__37_, r_n_219__36_, r_n_219__35_, r_n_219__34_, r_n_219__33_, r_n_219__32_, r_n_219__31_, r_n_219__30_, r_n_219__29_, r_n_219__28_, r_n_219__27_, r_n_219__26_, r_n_219__25_, r_n_219__24_, r_n_219__23_, r_n_219__22_, r_n_219__21_, r_n_219__20_, r_n_219__19_, r_n_219__18_, r_n_219__17_, r_n_219__16_, r_n_219__15_, r_n_219__14_, r_n_219__13_, r_n_219__12_, r_n_219__11_, r_n_219__10_, r_n_219__9_, r_n_219__8_, r_n_219__7_, r_n_219__6_, r_n_219__5_, r_n_219__4_, r_n_219__3_, r_n_219__2_, r_n_219__1_, r_n_219__0_ } = (N438)? { r_220__63_, r_220__62_, r_220__61_, r_220__60_, r_220__59_, r_220__58_, r_220__57_, r_220__56_, r_220__55_, r_220__54_, r_220__53_, r_220__52_, r_220__51_, r_220__50_, r_220__49_, r_220__48_, r_220__47_, r_220__46_, r_220__45_, r_220__44_, r_220__43_, r_220__42_, r_220__41_, r_220__40_, r_220__39_, r_220__38_, r_220__37_, r_220__36_, r_220__35_, r_220__34_, r_220__33_, r_220__32_, r_220__31_, r_220__30_, r_220__29_, r_220__28_, r_220__27_, r_220__26_, r_220__25_, r_220__24_, r_220__23_, r_220__22_, r_220__21_, r_220__20_, r_220__19_, r_220__18_, r_220__17_, r_220__16_, r_220__15_, r_220__14_, r_220__13_, r_220__12_, r_220__11_, r_220__10_, r_220__9_, r_220__8_, r_220__7_, r_220__6_, r_220__5_, r_220__4_, r_220__3_, r_220__2_, r_220__1_, r_220__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N439)? data_i : 1'b0;
  assign N438 = sel_i[438];
  assign N439 = N2123;
  assign { r_n_220__63_, r_n_220__62_, r_n_220__61_, r_n_220__60_, r_n_220__59_, r_n_220__58_, r_n_220__57_, r_n_220__56_, r_n_220__55_, r_n_220__54_, r_n_220__53_, r_n_220__52_, r_n_220__51_, r_n_220__50_, r_n_220__49_, r_n_220__48_, r_n_220__47_, r_n_220__46_, r_n_220__45_, r_n_220__44_, r_n_220__43_, r_n_220__42_, r_n_220__41_, r_n_220__40_, r_n_220__39_, r_n_220__38_, r_n_220__37_, r_n_220__36_, r_n_220__35_, r_n_220__34_, r_n_220__33_, r_n_220__32_, r_n_220__31_, r_n_220__30_, r_n_220__29_, r_n_220__28_, r_n_220__27_, r_n_220__26_, r_n_220__25_, r_n_220__24_, r_n_220__23_, r_n_220__22_, r_n_220__21_, r_n_220__20_, r_n_220__19_, r_n_220__18_, r_n_220__17_, r_n_220__16_, r_n_220__15_, r_n_220__14_, r_n_220__13_, r_n_220__12_, r_n_220__11_, r_n_220__10_, r_n_220__9_, r_n_220__8_, r_n_220__7_, r_n_220__6_, r_n_220__5_, r_n_220__4_, r_n_220__3_, r_n_220__2_, r_n_220__1_, r_n_220__0_ } = (N440)? { r_221__63_, r_221__62_, r_221__61_, r_221__60_, r_221__59_, r_221__58_, r_221__57_, r_221__56_, r_221__55_, r_221__54_, r_221__53_, r_221__52_, r_221__51_, r_221__50_, r_221__49_, r_221__48_, r_221__47_, r_221__46_, r_221__45_, r_221__44_, r_221__43_, r_221__42_, r_221__41_, r_221__40_, r_221__39_, r_221__38_, r_221__37_, r_221__36_, r_221__35_, r_221__34_, r_221__33_, r_221__32_, r_221__31_, r_221__30_, r_221__29_, r_221__28_, r_221__27_, r_221__26_, r_221__25_, r_221__24_, r_221__23_, r_221__22_, r_221__21_, r_221__20_, r_221__19_, r_221__18_, r_221__17_, r_221__16_, r_221__15_, r_221__14_, r_221__13_, r_221__12_, r_221__11_, r_221__10_, r_221__9_, r_221__8_, r_221__7_, r_221__6_, r_221__5_, r_221__4_, r_221__3_, r_221__2_, r_221__1_, r_221__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N441)? data_i : 1'b0;
  assign N440 = sel_i[440];
  assign N441 = N2128;
  assign { r_n_221__63_, r_n_221__62_, r_n_221__61_, r_n_221__60_, r_n_221__59_, r_n_221__58_, r_n_221__57_, r_n_221__56_, r_n_221__55_, r_n_221__54_, r_n_221__53_, r_n_221__52_, r_n_221__51_, r_n_221__50_, r_n_221__49_, r_n_221__48_, r_n_221__47_, r_n_221__46_, r_n_221__45_, r_n_221__44_, r_n_221__43_, r_n_221__42_, r_n_221__41_, r_n_221__40_, r_n_221__39_, r_n_221__38_, r_n_221__37_, r_n_221__36_, r_n_221__35_, r_n_221__34_, r_n_221__33_, r_n_221__32_, r_n_221__31_, r_n_221__30_, r_n_221__29_, r_n_221__28_, r_n_221__27_, r_n_221__26_, r_n_221__25_, r_n_221__24_, r_n_221__23_, r_n_221__22_, r_n_221__21_, r_n_221__20_, r_n_221__19_, r_n_221__18_, r_n_221__17_, r_n_221__16_, r_n_221__15_, r_n_221__14_, r_n_221__13_, r_n_221__12_, r_n_221__11_, r_n_221__10_, r_n_221__9_, r_n_221__8_, r_n_221__7_, r_n_221__6_, r_n_221__5_, r_n_221__4_, r_n_221__3_, r_n_221__2_, r_n_221__1_, r_n_221__0_ } = (N442)? { r_222__63_, r_222__62_, r_222__61_, r_222__60_, r_222__59_, r_222__58_, r_222__57_, r_222__56_, r_222__55_, r_222__54_, r_222__53_, r_222__52_, r_222__51_, r_222__50_, r_222__49_, r_222__48_, r_222__47_, r_222__46_, r_222__45_, r_222__44_, r_222__43_, r_222__42_, r_222__41_, r_222__40_, r_222__39_, r_222__38_, r_222__37_, r_222__36_, r_222__35_, r_222__34_, r_222__33_, r_222__32_, r_222__31_, r_222__30_, r_222__29_, r_222__28_, r_222__27_, r_222__26_, r_222__25_, r_222__24_, r_222__23_, r_222__22_, r_222__21_, r_222__20_, r_222__19_, r_222__18_, r_222__17_, r_222__16_, r_222__15_, r_222__14_, r_222__13_, r_222__12_, r_222__11_, r_222__10_, r_222__9_, r_222__8_, r_222__7_, r_222__6_, r_222__5_, r_222__4_, r_222__3_, r_222__2_, r_222__1_, r_222__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N443)? data_i : 1'b0;
  assign N442 = sel_i[442];
  assign N443 = N2133;
  assign { r_n_222__63_, r_n_222__62_, r_n_222__61_, r_n_222__60_, r_n_222__59_, r_n_222__58_, r_n_222__57_, r_n_222__56_, r_n_222__55_, r_n_222__54_, r_n_222__53_, r_n_222__52_, r_n_222__51_, r_n_222__50_, r_n_222__49_, r_n_222__48_, r_n_222__47_, r_n_222__46_, r_n_222__45_, r_n_222__44_, r_n_222__43_, r_n_222__42_, r_n_222__41_, r_n_222__40_, r_n_222__39_, r_n_222__38_, r_n_222__37_, r_n_222__36_, r_n_222__35_, r_n_222__34_, r_n_222__33_, r_n_222__32_, r_n_222__31_, r_n_222__30_, r_n_222__29_, r_n_222__28_, r_n_222__27_, r_n_222__26_, r_n_222__25_, r_n_222__24_, r_n_222__23_, r_n_222__22_, r_n_222__21_, r_n_222__20_, r_n_222__19_, r_n_222__18_, r_n_222__17_, r_n_222__16_, r_n_222__15_, r_n_222__14_, r_n_222__13_, r_n_222__12_, r_n_222__11_, r_n_222__10_, r_n_222__9_, r_n_222__8_, r_n_222__7_, r_n_222__6_, r_n_222__5_, r_n_222__4_, r_n_222__3_, r_n_222__2_, r_n_222__1_, r_n_222__0_ } = (N444)? { r_223__63_, r_223__62_, r_223__61_, r_223__60_, r_223__59_, r_223__58_, r_223__57_, r_223__56_, r_223__55_, r_223__54_, r_223__53_, r_223__52_, r_223__51_, r_223__50_, r_223__49_, r_223__48_, r_223__47_, r_223__46_, r_223__45_, r_223__44_, r_223__43_, r_223__42_, r_223__41_, r_223__40_, r_223__39_, r_223__38_, r_223__37_, r_223__36_, r_223__35_, r_223__34_, r_223__33_, r_223__32_, r_223__31_, r_223__30_, r_223__29_, r_223__28_, r_223__27_, r_223__26_, r_223__25_, r_223__24_, r_223__23_, r_223__22_, r_223__21_, r_223__20_, r_223__19_, r_223__18_, r_223__17_, r_223__16_, r_223__15_, r_223__14_, r_223__13_, r_223__12_, r_223__11_, r_223__10_, r_223__9_, r_223__8_, r_223__7_, r_223__6_, r_223__5_, r_223__4_, r_223__3_, r_223__2_, r_223__1_, r_223__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N445)? data_i : 1'b0;
  assign N444 = sel_i[444];
  assign N445 = N2138;
  assign { r_n_223__63_, r_n_223__62_, r_n_223__61_, r_n_223__60_, r_n_223__59_, r_n_223__58_, r_n_223__57_, r_n_223__56_, r_n_223__55_, r_n_223__54_, r_n_223__53_, r_n_223__52_, r_n_223__51_, r_n_223__50_, r_n_223__49_, r_n_223__48_, r_n_223__47_, r_n_223__46_, r_n_223__45_, r_n_223__44_, r_n_223__43_, r_n_223__42_, r_n_223__41_, r_n_223__40_, r_n_223__39_, r_n_223__38_, r_n_223__37_, r_n_223__36_, r_n_223__35_, r_n_223__34_, r_n_223__33_, r_n_223__32_, r_n_223__31_, r_n_223__30_, r_n_223__29_, r_n_223__28_, r_n_223__27_, r_n_223__26_, r_n_223__25_, r_n_223__24_, r_n_223__23_, r_n_223__22_, r_n_223__21_, r_n_223__20_, r_n_223__19_, r_n_223__18_, r_n_223__17_, r_n_223__16_, r_n_223__15_, r_n_223__14_, r_n_223__13_, r_n_223__12_, r_n_223__11_, r_n_223__10_, r_n_223__9_, r_n_223__8_, r_n_223__7_, r_n_223__6_, r_n_223__5_, r_n_223__4_, r_n_223__3_, r_n_223__2_, r_n_223__1_, r_n_223__0_ } = (N446)? { r_224__63_, r_224__62_, r_224__61_, r_224__60_, r_224__59_, r_224__58_, r_224__57_, r_224__56_, r_224__55_, r_224__54_, r_224__53_, r_224__52_, r_224__51_, r_224__50_, r_224__49_, r_224__48_, r_224__47_, r_224__46_, r_224__45_, r_224__44_, r_224__43_, r_224__42_, r_224__41_, r_224__40_, r_224__39_, r_224__38_, r_224__37_, r_224__36_, r_224__35_, r_224__34_, r_224__33_, r_224__32_, r_224__31_, r_224__30_, r_224__29_, r_224__28_, r_224__27_, r_224__26_, r_224__25_, r_224__24_, r_224__23_, r_224__22_, r_224__21_, r_224__20_, r_224__19_, r_224__18_, r_224__17_, r_224__16_, r_224__15_, r_224__14_, r_224__13_, r_224__12_, r_224__11_, r_224__10_, r_224__9_, r_224__8_, r_224__7_, r_224__6_, r_224__5_, r_224__4_, r_224__3_, r_224__2_, r_224__1_, r_224__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N447)? data_i : 1'b0;
  assign N446 = sel_i[446];
  assign N447 = N2143;
  assign { r_n_224__63_, r_n_224__62_, r_n_224__61_, r_n_224__60_, r_n_224__59_, r_n_224__58_, r_n_224__57_, r_n_224__56_, r_n_224__55_, r_n_224__54_, r_n_224__53_, r_n_224__52_, r_n_224__51_, r_n_224__50_, r_n_224__49_, r_n_224__48_, r_n_224__47_, r_n_224__46_, r_n_224__45_, r_n_224__44_, r_n_224__43_, r_n_224__42_, r_n_224__41_, r_n_224__40_, r_n_224__39_, r_n_224__38_, r_n_224__37_, r_n_224__36_, r_n_224__35_, r_n_224__34_, r_n_224__33_, r_n_224__32_, r_n_224__31_, r_n_224__30_, r_n_224__29_, r_n_224__28_, r_n_224__27_, r_n_224__26_, r_n_224__25_, r_n_224__24_, r_n_224__23_, r_n_224__22_, r_n_224__21_, r_n_224__20_, r_n_224__19_, r_n_224__18_, r_n_224__17_, r_n_224__16_, r_n_224__15_, r_n_224__14_, r_n_224__13_, r_n_224__12_, r_n_224__11_, r_n_224__10_, r_n_224__9_, r_n_224__8_, r_n_224__7_, r_n_224__6_, r_n_224__5_, r_n_224__4_, r_n_224__3_, r_n_224__2_, r_n_224__1_, r_n_224__0_ } = (N448)? { r_225__63_, r_225__62_, r_225__61_, r_225__60_, r_225__59_, r_225__58_, r_225__57_, r_225__56_, r_225__55_, r_225__54_, r_225__53_, r_225__52_, r_225__51_, r_225__50_, r_225__49_, r_225__48_, r_225__47_, r_225__46_, r_225__45_, r_225__44_, r_225__43_, r_225__42_, r_225__41_, r_225__40_, r_225__39_, r_225__38_, r_225__37_, r_225__36_, r_225__35_, r_225__34_, r_225__33_, r_225__32_, r_225__31_, r_225__30_, r_225__29_, r_225__28_, r_225__27_, r_225__26_, r_225__25_, r_225__24_, r_225__23_, r_225__22_, r_225__21_, r_225__20_, r_225__19_, r_225__18_, r_225__17_, r_225__16_, r_225__15_, r_225__14_, r_225__13_, r_225__12_, r_225__11_, r_225__10_, r_225__9_, r_225__8_, r_225__7_, r_225__6_, r_225__5_, r_225__4_, r_225__3_, r_225__2_, r_225__1_, r_225__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N449)? data_i : 1'b0;
  assign N448 = sel_i[448];
  assign N449 = N2148;
  assign { r_n_225__63_, r_n_225__62_, r_n_225__61_, r_n_225__60_, r_n_225__59_, r_n_225__58_, r_n_225__57_, r_n_225__56_, r_n_225__55_, r_n_225__54_, r_n_225__53_, r_n_225__52_, r_n_225__51_, r_n_225__50_, r_n_225__49_, r_n_225__48_, r_n_225__47_, r_n_225__46_, r_n_225__45_, r_n_225__44_, r_n_225__43_, r_n_225__42_, r_n_225__41_, r_n_225__40_, r_n_225__39_, r_n_225__38_, r_n_225__37_, r_n_225__36_, r_n_225__35_, r_n_225__34_, r_n_225__33_, r_n_225__32_, r_n_225__31_, r_n_225__30_, r_n_225__29_, r_n_225__28_, r_n_225__27_, r_n_225__26_, r_n_225__25_, r_n_225__24_, r_n_225__23_, r_n_225__22_, r_n_225__21_, r_n_225__20_, r_n_225__19_, r_n_225__18_, r_n_225__17_, r_n_225__16_, r_n_225__15_, r_n_225__14_, r_n_225__13_, r_n_225__12_, r_n_225__11_, r_n_225__10_, r_n_225__9_, r_n_225__8_, r_n_225__7_, r_n_225__6_, r_n_225__5_, r_n_225__4_, r_n_225__3_, r_n_225__2_, r_n_225__1_, r_n_225__0_ } = (N450)? { r_226__63_, r_226__62_, r_226__61_, r_226__60_, r_226__59_, r_226__58_, r_226__57_, r_226__56_, r_226__55_, r_226__54_, r_226__53_, r_226__52_, r_226__51_, r_226__50_, r_226__49_, r_226__48_, r_226__47_, r_226__46_, r_226__45_, r_226__44_, r_226__43_, r_226__42_, r_226__41_, r_226__40_, r_226__39_, r_226__38_, r_226__37_, r_226__36_, r_226__35_, r_226__34_, r_226__33_, r_226__32_, r_226__31_, r_226__30_, r_226__29_, r_226__28_, r_226__27_, r_226__26_, r_226__25_, r_226__24_, r_226__23_, r_226__22_, r_226__21_, r_226__20_, r_226__19_, r_226__18_, r_226__17_, r_226__16_, r_226__15_, r_226__14_, r_226__13_, r_226__12_, r_226__11_, r_226__10_, r_226__9_, r_226__8_, r_226__7_, r_226__6_, r_226__5_, r_226__4_, r_226__3_, r_226__2_, r_226__1_, r_226__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N451)? data_i : 1'b0;
  assign N450 = sel_i[450];
  assign N451 = N2153;
  assign { r_n_226__63_, r_n_226__62_, r_n_226__61_, r_n_226__60_, r_n_226__59_, r_n_226__58_, r_n_226__57_, r_n_226__56_, r_n_226__55_, r_n_226__54_, r_n_226__53_, r_n_226__52_, r_n_226__51_, r_n_226__50_, r_n_226__49_, r_n_226__48_, r_n_226__47_, r_n_226__46_, r_n_226__45_, r_n_226__44_, r_n_226__43_, r_n_226__42_, r_n_226__41_, r_n_226__40_, r_n_226__39_, r_n_226__38_, r_n_226__37_, r_n_226__36_, r_n_226__35_, r_n_226__34_, r_n_226__33_, r_n_226__32_, r_n_226__31_, r_n_226__30_, r_n_226__29_, r_n_226__28_, r_n_226__27_, r_n_226__26_, r_n_226__25_, r_n_226__24_, r_n_226__23_, r_n_226__22_, r_n_226__21_, r_n_226__20_, r_n_226__19_, r_n_226__18_, r_n_226__17_, r_n_226__16_, r_n_226__15_, r_n_226__14_, r_n_226__13_, r_n_226__12_, r_n_226__11_, r_n_226__10_, r_n_226__9_, r_n_226__8_, r_n_226__7_, r_n_226__6_, r_n_226__5_, r_n_226__4_, r_n_226__3_, r_n_226__2_, r_n_226__1_, r_n_226__0_ } = (N452)? { r_227__63_, r_227__62_, r_227__61_, r_227__60_, r_227__59_, r_227__58_, r_227__57_, r_227__56_, r_227__55_, r_227__54_, r_227__53_, r_227__52_, r_227__51_, r_227__50_, r_227__49_, r_227__48_, r_227__47_, r_227__46_, r_227__45_, r_227__44_, r_227__43_, r_227__42_, r_227__41_, r_227__40_, r_227__39_, r_227__38_, r_227__37_, r_227__36_, r_227__35_, r_227__34_, r_227__33_, r_227__32_, r_227__31_, r_227__30_, r_227__29_, r_227__28_, r_227__27_, r_227__26_, r_227__25_, r_227__24_, r_227__23_, r_227__22_, r_227__21_, r_227__20_, r_227__19_, r_227__18_, r_227__17_, r_227__16_, r_227__15_, r_227__14_, r_227__13_, r_227__12_, r_227__11_, r_227__10_, r_227__9_, r_227__8_, r_227__7_, r_227__6_, r_227__5_, r_227__4_, r_227__3_, r_227__2_, r_227__1_, r_227__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N453)? data_i : 1'b0;
  assign N452 = sel_i[452];
  assign N453 = N2158;
  assign { r_n_227__63_, r_n_227__62_, r_n_227__61_, r_n_227__60_, r_n_227__59_, r_n_227__58_, r_n_227__57_, r_n_227__56_, r_n_227__55_, r_n_227__54_, r_n_227__53_, r_n_227__52_, r_n_227__51_, r_n_227__50_, r_n_227__49_, r_n_227__48_, r_n_227__47_, r_n_227__46_, r_n_227__45_, r_n_227__44_, r_n_227__43_, r_n_227__42_, r_n_227__41_, r_n_227__40_, r_n_227__39_, r_n_227__38_, r_n_227__37_, r_n_227__36_, r_n_227__35_, r_n_227__34_, r_n_227__33_, r_n_227__32_, r_n_227__31_, r_n_227__30_, r_n_227__29_, r_n_227__28_, r_n_227__27_, r_n_227__26_, r_n_227__25_, r_n_227__24_, r_n_227__23_, r_n_227__22_, r_n_227__21_, r_n_227__20_, r_n_227__19_, r_n_227__18_, r_n_227__17_, r_n_227__16_, r_n_227__15_, r_n_227__14_, r_n_227__13_, r_n_227__12_, r_n_227__11_, r_n_227__10_, r_n_227__9_, r_n_227__8_, r_n_227__7_, r_n_227__6_, r_n_227__5_, r_n_227__4_, r_n_227__3_, r_n_227__2_, r_n_227__1_, r_n_227__0_ } = (N454)? { r_228__63_, r_228__62_, r_228__61_, r_228__60_, r_228__59_, r_228__58_, r_228__57_, r_228__56_, r_228__55_, r_228__54_, r_228__53_, r_228__52_, r_228__51_, r_228__50_, r_228__49_, r_228__48_, r_228__47_, r_228__46_, r_228__45_, r_228__44_, r_228__43_, r_228__42_, r_228__41_, r_228__40_, r_228__39_, r_228__38_, r_228__37_, r_228__36_, r_228__35_, r_228__34_, r_228__33_, r_228__32_, r_228__31_, r_228__30_, r_228__29_, r_228__28_, r_228__27_, r_228__26_, r_228__25_, r_228__24_, r_228__23_, r_228__22_, r_228__21_, r_228__20_, r_228__19_, r_228__18_, r_228__17_, r_228__16_, r_228__15_, r_228__14_, r_228__13_, r_228__12_, r_228__11_, r_228__10_, r_228__9_, r_228__8_, r_228__7_, r_228__6_, r_228__5_, r_228__4_, r_228__3_, r_228__2_, r_228__1_, r_228__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N455)? data_i : 1'b0;
  assign N454 = sel_i[454];
  assign N455 = N2163;
  assign { r_n_228__63_, r_n_228__62_, r_n_228__61_, r_n_228__60_, r_n_228__59_, r_n_228__58_, r_n_228__57_, r_n_228__56_, r_n_228__55_, r_n_228__54_, r_n_228__53_, r_n_228__52_, r_n_228__51_, r_n_228__50_, r_n_228__49_, r_n_228__48_, r_n_228__47_, r_n_228__46_, r_n_228__45_, r_n_228__44_, r_n_228__43_, r_n_228__42_, r_n_228__41_, r_n_228__40_, r_n_228__39_, r_n_228__38_, r_n_228__37_, r_n_228__36_, r_n_228__35_, r_n_228__34_, r_n_228__33_, r_n_228__32_, r_n_228__31_, r_n_228__30_, r_n_228__29_, r_n_228__28_, r_n_228__27_, r_n_228__26_, r_n_228__25_, r_n_228__24_, r_n_228__23_, r_n_228__22_, r_n_228__21_, r_n_228__20_, r_n_228__19_, r_n_228__18_, r_n_228__17_, r_n_228__16_, r_n_228__15_, r_n_228__14_, r_n_228__13_, r_n_228__12_, r_n_228__11_, r_n_228__10_, r_n_228__9_, r_n_228__8_, r_n_228__7_, r_n_228__6_, r_n_228__5_, r_n_228__4_, r_n_228__3_, r_n_228__2_, r_n_228__1_, r_n_228__0_ } = (N456)? { r_229__63_, r_229__62_, r_229__61_, r_229__60_, r_229__59_, r_229__58_, r_229__57_, r_229__56_, r_229__55_, r_229__54_, r_229__53_, r_229__52_, r_229__51_, r_229__50_, r_229__49_, r_229__48_, r_229__47_, r_229__46_, r_229__45_, r_229__44_, r_229__43_, r_229__42_, r_229__41_, r_229__40_, r_229__39_, r_229__38_, r_229__37_, r_229__36_, r_229__35_, r_229__34_, r_229__33_, r_229__32_, r_229__31_, r_229__30_, r_229__29_, r_229__28_, r_229__27_, r_229__26_, r_229__25_, r_229__24_, r_229__23_, r_229__22_, r_229__21_, r_229__20_, r_229__19_, r_229__18_, r_229__17_, r_229__16_, r_229__15_, r_229__14_, r_229__13_, r_229__12_, r_229__11_, r_229__10_, r_229__9_, r_229__8_, r_229__7_, r_229__6_, r_229__5_, r_229__4_, r_229__3_, r_229__2_, r_229__1_, r_229__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N457)? data_i : 1'b0;
  assign N456 = sel_i[456];
  assign N457 = N2168;
  assign { r_n_229__63_, r_n_229__62_, r_n_229__61_, r_n_229__60_, r_n_229__59_, r_n_229__58_, r_n_229__57_, r_n_229__56_, r_n_229__55_, r_n_229__54_, r_n_229__53_, r_n_229__52_, r_n_229__51_, r_n_229__50_, r_n_229__49_, r_n_229__48_, r_n_229__47_, r_n_229__46_, r_n_229__45_, r_n_229__44_, r_n_229__43_, r_n_229__42_, r_n_229__41_, r_n_229__40_, r_n_229__39_, r_n_229__38_, r_n_229__37_, r_n_229__36_, r_n_229__35_, r_n_229__34_, r_n_229__33_, r_n_229__32_, r_n_229__31_, r_n_229__30_, r_n_229__29_, r_n_229__28_, r_n_229__27_, r_n_229__26_, r_n_229__25_, r_n_229__24_, r_n_229__23_, r_n_229__22_, r_n_229__21_, r_n_229__20_, r_n_229__19_, r_n_229__18_, r_n_229__17_, r_n_229__16_, r_n_229__15_, r_n_229__14_, r_n_229__13_, r_n_229__12_, r_n_229__11_, r_n_229__10_, r_n_229__9_, r_n_229__8_, r_n_229__7_, r_n_229__6_, r_n_229__5_, r_n_229__4_, r_n_229__3_, r_n_229__2_, r_n_229__1_, r_n_229__0_ } = (N458)? { r_230__63_, r_230__62_, r_230__61_, r_230__60_, r_230__59_, r_230__58_, r_230__57_, r_230__56_, r_230__55_, r_230__54_, r_230__53_, r_230__52_, r_230__51_, r_230__50_, r_230__49_, r_230__48_, r_230__47_, r_230__46_, r_230__45_, r_230__44_, r_230__43_, r_230__42_, r_230__41_, r_230__40_, r_230__39_, r_230__38_, r_230__37_, r_230__36_, r_230__35_, r_230__34_, r_230__33_, r_230__32_, r_230__31_, r_230__30_, r_230__29_, r_230__28_, r_230__27_, r_230__26_, r_230__25_, r_230__24_, r_230__23_, r_230__22_, r_230__21_, r_230__20_, r_230__19_, r_230__18_, r_230__17_, r_230__16_, r_230__15_, r_230__14_, r_230__13_, r_230__12_, r_230__11_, r_230__10_, r_230__9_, r_230__8_, r_230__7_, r_230__6_, r_230__5_, r_230__4_, r_230__3_, r_230__2_, r_230__1_, r_230__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N459)? data_i : 1'b0;
  assign N458 = sel_i[458];
  assign N459 = N2173;
  assign { r_n_230__63_, r_n_230__62_, r_n_230__61_, r_n_230__60_, r_n_230__59_, r_n_230__58_, r_n_230__57_, r_n_230__56_, r_n_230__55_, r_n_230__54_, r_n_230__53_, r_n_230__52_, r_n_230__51_, r_n_230__50_, r_n_230__49_, r_n_230__48_, r_n_230__47_, r_n_230__46_, r_n_230__45_, r_n_230__44_, r_n_230__43_, r_n_230__42_, r_n_230__41_, r_n_230__40_, r_n_230__39_, r_n_230__38_, r_n_230__37_, r_n_230__36_, r_n_230__35_, r_n_230__34_, r_n_230__33_, r_n_230__32_, r_n_230__31_, r_n_230__30_, r_n_230__29_, r_n_230__28_, r_n_230__27_, r_n_230__26_, r_n_230__25_, r_n_230__24_, r_n_230__23_, r_n_230__22_, r_n_230__21_, r_n_230__20_, r_n_230__19_, r_n_230__18_, r_n_230__17_, r_n_230__16_, r_n_230__15_, r_n_230__14_, r_n_230__13_, r_n_230__12_, r_n_230__11_, r_n_230__10_, r_n_230__9_, r_n_230__8_, r_n_230__7_, r_n_230__6_, r_n_230__5_, r_n_230__4_, r_n_230__3_, r_n_230__2_, r_n_230__1_, r_n_230__0_ } = (N460)? { r_231__63_, r_231__62_, r_231__61_, r_231__60_, r_231__59_, r_231__58_, r_231__57_, r_231__56_, r_231__55_, r_231__54_, r_231__53_, r_231__52_, r_231__51_, r_231__50_, r_231__49_, r_231__48_, r_231__47_, r_231__46_, r_231__45_, r_231__44_, r_231__43_, r_231__42_, r_231__41_, r_231__40_, r_231__39_, r_231__38_, r_231__37_, r_231__36_, r_231__35_, r_231__34_, r_231__33_, r_231__32_, r_231__31_, r_231__30_, r_231__29_, r_231__28_, r_231__27_, r_231__26_, r_231__25_, r_231__24_, r_231__23_, r_231__22_, r_231__21_, r_231__20_, r_231__19_, r_231__18_, r_231__17_, r_231__16_, r_231__15_, r_231__14_, r_231__13_, r_231__12_, r_231__11_, r_231__10_, r_231__9_, r_231__8_, r_231__7_, r_231__6_, r_231__5_, r_231__4_, r_231__3_, r_231__2_, r_231__1_, r_231__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N461)? data_i : 1'b0;
  assign N460 = sel_i[460];
  assign N461 = N2178;
  assign { r_n_231__63_, r_n_231__62_, r_n_231__61_, r_n_231__60_, r_n_231__59_, r_n_231__58_, r_n_231__57_, r_n_231__56_, r_n_231__55_, r_n_231__54_, r_n_231__53_, r_n_231__52_, r_n_231__51_, r_n_231__50_, r_n_231__49_, r_n_231__48_, r_n_231__47_, r_n_231__46_, r_n_231__45_, r_n_231__44_, r_n_231__43_, r_n_231__42_, r_n_231__41_, r_n_231__40_, r_n_231__39_, r_n_231__38_, r_n_231__37_, r_n_231__36_, r_n_231__35_, r_n_231__34_, r_n_231__33_, r_n_231__32_, r_n_231__31_, r_n_231__30_, r_n_231__29_, r_n_231__28_, r_n_231__27_, r_n_231__26_, r_n_231__25_, r_n_231__24_, r_n_231__23_, r_n_231__22_, r_n_231__21_, r_n_231__20_, r_n_231__19_, r_n_231__18_, r_n_231__17_, r_n_231__16_, r_n_231__15_, r_n_231__14_, r_n_231__13_, r_n_231__12_, r_n_231__11_, r_n_231__10_, r_n_231__9_, r_n_231__8_, r_n_231__7_, r_n_231__6_, r_n_231__5_, r_n_231__4_, r_n_231__3_, r_n_231__2_, r_n_231__1_, r_n_231__0_ } = (N462)? { r_232__63_, r_232__62_, r_232__61_, r_232__60_, r_232__59_, r_232__58_, r_232__57_, r_232__56_, r_232__55_, r_232__54_, r_232__53_, r_232__52_, r_232__51_, r_232__50_, r_232__49_, r_232__48_, r_232__47_, r_232__46_, r_232__45_, r_232__44_, r_232__43_, r_232__42_, r_232__41_, r_232__40_, r_232__39_, r_232__38_, r_232__37_, r_232__36_, r_232__35_, r_232__34_, r_232__33_, r_232__32_, r_232__31_, r_232__30_, r_232__29_, r_232__28_, r_232__27_, r_232__26_, r_232__25_, r_232__24_, r_232__23_, r_232__22_, r_232__21_, r_232__20_, r_232__19_, r_232__18_, r_232__17_, r_232__16_, r_232__15_, r_232__14_, r_232__13_, r_232__12_, r_232__11_, r_232__10_, r_232__9_, r_232__8_, r_232__7_, r_232__6_, r_232__5_, r_232__4_, r_232__3_, r_232__2_, r_232__1_, r_232__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N463)? data_i : 1'b0;
  assign N462 = sel_i[462];
  assign N463 = N2183;
  assign { r_n_232__63_, r_n_232__62_, r_n_232__61_, r_n_232__60_, r_n_232__59_, r_n_232__58_, r_n_232__57_, r_n_232__56_, r_n_232__55_, r_n_232__54_, r_n_232__53_, r_n_232__52_, r_n_232__51_, r_n_232__50_, r_n_232__49_, r_n_232__48_, r_n_232__47_, r_n_232__46_, r_n_232__45_, r_n_232__44_, r_n_232__43_, r_n_232__42_, r_n_232__41_, r_n_232__40_, r_n_232__39_, r_n_232__38_, r_n_232__37_, r_n_232__36_, r_n_232__35_, r_n_232__34_, r_n_232__33_, r_n_232__32_, r_n_232__31_, r_n_232__30_, r_n_232__29_, r_n_232__28_, r_n_232__27_, r_n_232__26_, r_n_232__25_, r_n_232__24_, r_n_232__23_, r_n_232__22_, r_n_232__21_, r_n_232__20_, r_n_232__19_, r_n_232__18_, r_n_232__17_, r_n_232__16_, r_n_232__15_, r_n_232__14_, r_n_232__13_, r_n_232__12_, r_n_232__11_, r_n_232__10_, r_n_232__9_, r_n_232__8_, r_n_232__7_, r_n_232__6_, r_n_232__5_, r_n_232__4_, r_n_232__3_, r_n_232__2_, r_n_232__1_, r_n_232__0_ } = (N464)? { r_233__63_, r_233__62_, r_233__61_, r_233__60_, r_233__59_, r_233__58_, r_233__57_, r_233__56_, r_233__55_, r_233__54_, r_233__53_, r_233__52_, r_233__51_, r_233__50_, r_233__49_, r_233__48_, r_233__47_, r_233__46_, r_233__45_, r_233__44_, r_233__43_, r_233__42_, r_233__41_, r_233__40_, r_233__39_, r_233__38_, r_233__37_, r_233__36_, r_233__35_, r_233__34_, r_233__33_, r_233__32_, r_233__31_, r_233__30_, r_233__29_, r_233__28_, r_233__27_, r_233__26_, r_233__25_, r_233__24_, r_233__23_, r_233__22_, r_233__21_, r_233__20_, r_233__19_, r_233__18_, r_233__17_, r_233__16_, r_233__15_, r_233__14_, r_233__13_, r_233__12_, r_233__11_, r_233__10_, r_233__9_, r_233__8_, r_233__7_, r_233__6_, r_233__5_, r_233__4_, r_233__3_, r_233__2_, r_233__1_, r_233__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N465)? data_i : 1'b0;
  assign N464 = sel_i[464];
  assign N465 = N2188;
  assign { r_n_233__63_, r_n_233__62_, r_n_233__61_, r_n_233__60_, r_n_233__59_, r_n_233__58_, r_n_233__57_, r_n_233__56_, r_n_233__55_, r_n_233__54_, r_n_233__53_, r_n_233__52_, r_n_233__51_, r_n_233__50_, r_n_233__49_, r_n_233__48_, r_n_233__47_, r_n_233__46_, r_n_233__45_, r_n_233__44_, r_n_233__43_, r_n_233__42_, r_n_233__41_, r_n_233__40_, r_n_233__39_, r_n_233__38_, r_n_233__37_, r_n_233__36_, r_n_233__35_, r_n_233__34_, r_n_233__33_, r_n_233__32_, r_n_233__31_, r_n_233__30_, r_n_233__29_, r_n_233__28_, r_n_233__27_, r_n_233__26_, r_n_233__25_, r_n_233__24_, r_n_233__23_, r_n_233__22_, r_n_233__21_, r_n_233__20_, r_n_233__19_, r_n_233__18_, r_n_233__17_, r_n_233__16_, r_n_233__15_, r_n_233__14_, r_n_233__13_, r_n_233__12_, r_n_233__11_, r_n_233__10_, r_n_233__9_, r_n_233__8_, r_n_233__7_, r_n_233__6_, r_n_233__5_, r_n_233__4_, r_n_233__3_, r_n_233__2_, r_n_233__1_, r_n_233__0_ } = (N466)? { r_234__63_, r_234__62_, r_234__61_, r_234__60_, r_234__59_, r_234__58_, r_234__57_, r_234__56_, r_234__55_, r_234__54_, r_234__53_, r_234__52_, r_234__51_, r_234__50_, r_234__49_, r_234__48_, r_234__47_, r_234__46_, r_234__45_, r_234__44_, r_234__43_, r_234__42_, r_234__41_, r_234__40_, r_234__39_, r_234__38_, r_234__37_, r_234__36_, r_234__35_, r_234__34_, r_234__33_, r_234__32_, r_234__31_, r_234__30_, r_234__29_, r_234__28_, r_234__27_, r_234__26_, r_234__25_, r_234__24_, r_234__23_, r_234__22_, r_234__21_, r_234__20_, r_234__19_, r_234__18_, r_234__17_, r_234__16_, r_234__15_, r_234__14_, r_234__13_, r_234__12_, r_234__11_, r_234__10_, r_234__9_, r_234__8_, r_234__7_, r_234__6_, r_234__5_, r_234__4_, r_234__3_, r_234__2_, r_234__1_, r_234__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N467)? data_i : 1'b0;
  assign N466 = sel_i[466];
  assign N467 = N2193;
  assign { r_n_234__63_, r_n_234__62_, r_n_234__61_, r_n_234__60_, r_n_234__59_, r_n_234__58_, r_n_234__57_, r_n_234__56_, r_n_234__55_, r_n_234__54_, r_n_234__53_, r_n_234__52_, r_n_234__51_, r_n_234__50_, r_n_234__49_, r_n_234__48_, r_n_234__47_, r_n_234__46_, r_n_234__45_, r_n_234__44_, r_n_234__43_, r_n_234__42_, r_n_234__41_, r_n_234__40_, r_n_234__39_, r_n_234__38_, r_n_234__37_, r_n_234__36_, r_n_234__35_, r_n_234__34_, r_n_234__33_, r_n_234__32_, r_n_234__31_, r_n_234__30_, r_n_234__29_, r_n_234__28_, r_n_234__27_, r_n_234__26_, r_n_234__25_, r_n_234__24_, r_n_234__23_, r_n_234__22_, r_n_234__21_, r_n_234__20_, r_n_234__19_, r_n_234__18_, r_n_234__17_, r_n_234__16_, r_n_234__15_, r_n_234__14_, r_n_234__13_, r_n_234__12_, r_n_234__11_, r_n_234__10_, r_n_234__9_, r_n_234__8_, r_n_234__7_, r_n_234__6_, r_n_234__5_, r_n_234__4_, r_n_234__3_, r_n_234__2_, r_n_234__1_, r_n_234__0_ } = (N468)? { r_235__63_, r_235__62_, r_235__61_, r_235__60_, r_235__59_, r_235__58_, r_235__57_, r_235__56_, r_235__55_, r_235__54_, r_235__53_, r_235__52_, r_235__51_, r_235__50_, r_235__49_, r_235__48_, r_235__47_, r_235__46_, r_235__45_, r_235__44_, r_235__43_, r_235__42_, r_235__41_, r_235__40_, r_235__39_, r_235__38_, r_235__37_, r_235__36_, r_235__35_, r_235__34_, r_235__33_, r_235__32_, r_235__31_, r_235__30_, r_235__29_, r_235__28_, r_235__27_, r_235__26_, r_235__25_, r_235__24_, r_235__23_, r_235__22_, r_235__21_, r_235__20_, r_235__19_, r_235__18_, r_235__17_, r_235__16_, r_235__15_, r_235__14_, r_235__13_, r_235__12_, r_235__11_, r_235__10_, r_235__9_, r_235__8_, r_235__7_, r_235__6_, r_235__5_, r_235__4_, r_235__3_, r_235__2_, r_235__1_, r_235__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N469)? data_i : 1'b0;
  assign N468 = sel_i[468];
  assign N469 = N2198;
  assign { r_n_235__63_, r_n_235__62_, r_n_235__61_, r_n_235__60_, r_n_235__59_, r_n_235__58_, r_n_235__57_, r_n_235__56_, r_n_235__55_, r_n_235__54_, r_n_235__53_, r_n_235__52_, r_n_235__51_, r_n_235__50_, r_n_235__49_, r_n_235__48_, r_n_235__47_, r_n_235__46_, r_n_235__45_, r_n_235__44_, r_n_235__43_, r_n_235__42_, r_n_235__41_, r_n_235__40_, r_n_235__39_, r_n_235__38_, r_n_235__37_, r_n_235__36_, r_n_235__35_, r_n_235__34_, r_n_235__33_, r_n_235__32_, r_n_235__31_, r_n_235__30_, r_n_235__29_, r_n_235__28_, r_n_235__27_, r_n_235__26_, r_n_235__25_, r_n_235__24_, r_n_235__23_, r_n_235__22_, r_n_235__21_, r_n_235__20_, r_n_235__19_, r_n_235__18_, r_n_235__17_, r_n_235__16_, r_n_235__15_, r_n_235__14_, r_n_235__13_, r_n_235__12_, r_n_235__11_, r_n_235__10_, r_n_235__9_, r_n_235__8_, r_n_235__7_, r_n_235__6_, r_n_235__5_, r_n_235__4_, r_n_235__3_, r_n_235__2_, r_n_235__1_, r_n_235__0_ } = (N470)? { r_236__63_, r_236__62_, r_236__61_, r_236__60_, r_236__59_, r_236__58_, r_236__57_, r_236__56_, r_236__55_, r_236__54_, r_236__53_, r_236__52_, r_236__51_, r_236__50_, r_236__49_, r_236__48_, r_236__47_, r_236__46_, r_236__45_, r_236__44_, r_236__43_, r_236__42_, r_236__41_, r_236__40_, r_236__39_, r_236__38_, r_236__37_, r_236__36_, r_236__35_, r_236__34_, r_236__33_, r_236__32_, r_236__31_, r_236__30_, r_236__29_, r_236__28_, r_236__27_, r_236__26_, r_236__25_, r_236__24_, r_236__23_, r_236__22_, r_236__21_, r_236__20_, r_236__19_, r_236__18_, r_236__17_, r_236__16_, r_236__15_, r_236__14_, r_236__13_, r_236__12_, r_236__11_, r_236__10_, r_236__9_, r_236__8_, r_236__7_, r_236__6_, r_236__5_, r_236__4_, r_236__3_, r_236__2_, r_236__1_, r_236__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N471)? data_i : 1'b0;
  assign N470 = sel_i[470];
  assign N471 = N2203;
  assign { r_n_236__63_, r_n_236__62_, r_n_236__61_, r_n_236__60_, r_n_236__59_, r_n_236__58_, r_n_236__57_, r_n_236__56_, r_n_236__55_, r_n_236__54_, r_n_236__53_, r_n_236__52_, r_n_236__51_, r_n_236__50_, r_n_236__49_, r_n_236__48_, r_n_236__47_, r_n_236__46_, r_n_236__45_, r_n_236__44_, r_n_236__43_, r_n_236__42_, r_n_236__41_, r_n_236__40_, r_n_236__39_, r_n_236__38_, r_n_236__37_, r_n_236__36_, r_n_236__35_, r_n_236__34_, r_n_236__33_, r_n_236__32_, r_n_236__31_, r_n_236__30_, r_n_236__29_, r_n_236__28_, r_n_236__27_, r_n_236__26_, r_n_236__25_, r_n_236__24_, r_n_236__23_, r_n_236__22_, r_n_236__21_, r_n_236__20_, r_n_236__19_, r_n_236__18_, r_n_236__17_, r_n_236__16_, r_n_236__15_, r_n_236__14_, r_n_236__13_, r_n_236__12_, r_n_236__11_, r_n_236__10_, r_n_236__9_, r_n_236__8_, r_n_236__7_, r_n_236__6_, r_n_236__5_, r_n_236__4_, r_n_236__3_, r_n_236__2_, r_n_236__1_, r_n_236__0_ } = (N472)? { r_237__63_, r_237__62_, r_237__61_, r_237__60_, r_237__59_, r_237__58_, r_237__57_, r_237__56_, r_237__55_, r_237__54_, r_237__53_, r_237__52_, r_237__51_, r_237__50_, r_237__49_, r_237__48_, r_237__47_, r_237__46_, r_237__45_, r_237__44_, r_237__43_, r_237__42_, r_237__41_, r_237__40_, r_237__39_, r_237__38_, r_237__37_, r_237__36_, r_237__35_, r_237__34_, r_237__33_, r_237__32_, r_237__31_, r_237__30_, r_237__29_, r_237__28_, r_237__27_, r_237__26_, r_237__25_, r_237__24_, r_237__23_, r_237__22_, r_237__21_, r_237__20_, r_237__19_, r_237__18_, r_237__17_, r_237__16_, r_237__15_, r_237__14_, r_237__13_, r_237__12_, r_237__11_, r_237__10_, r_237__9_, r_237__8_, r_237__7_, r_237__6_, r_237__5_, r_237__4_, r_237__3_, r_237__2_, r_237__1_, r_237__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N473)? data_i : 1'b0;
  assign N472 = sel_i[472];
  assign N473 = N2208;
  assign { r_n_237__63_, r_n_237__62_, r_n_237__61_, r_n_237__60_, r_n_237__59_, r_n_237__58_, r_n_237__57_, r_n_237__56_, r_n_237__55_, r_n_237__54_, r_n_237__53_, r_n_237__52_, r_n_237__51_, r_n_237__50_, r_n_237__49_, r_n_237__48_, r_n_237__47_, r_n_237__46_, r_n_237__45_, r_n_237__44_, r_n_237__43_, r_n_237__42_, r_n_237__41_, r_n_237__40_, r_n_237__39_, r_n_237__38_, r_n_237__37_, r_n_237__36_, r_n_237__35_, r_n_237__34_, r_n_237__33_, r_n_237__32_, r_n_237__31_, r_n_237__30_, r_n_237__29_, r_n_237__28_, r_n_237__27_, r_n_237__26_, r_n_237__25_, r_n_237__24_, r_n_237__23_, r_n_237__22_, r_n_237__21_, r_n_237__20_, r_n_237__19_, r_n_237__18_, r_n_237__17_, r_n_237__16_, r_n_237__15_, r_n_237__14_, r_n_237__13_, r_n_237__12_, r_n_237__11_, r_n_237__10_, r_n_237__9_, r_n_237__8_, r_n_237__7_, r_n_237__6_, r_n_237__5_, r_n_237__4_, r_n_237__3_, r_n_237__2_, r_n_237__1_, r_n_237__0_ } = (N474)? { r_238__63_, r_238__62_, r_238__61_, r_238__60_, r_238__59_, r_238__58_, r_238__57_, r_238__56_, r_238__55_, r_238__54_, r_238__53_, r_238__52_, r_238__51_, r_238__50_, r_238__49_, r_238__48_, r_238__47_, r_238__46_, r_238__45_, r_238__44_, r_238__43_, r_238__42_, r_238__41_, r_238__40_, r_238__39_, r_238__38_, r_238__37_, r_238__36_, r_238__35_, r_238__34_, r_238__33_, r_238__32_, r_238__31_, r_238__30_, r_238__29_, r_238__28_, r_238__27_, r_238__26_, r_238__25_, r_238__24_, r_238__23_, r_238__22_, r_238__21_, r_238__20_, r_238__19_, r_238__18_, r_238__17_, r_238__16_, r_238__15_, r_238__14_, r_238__13_, r_238__12_, r_238__11_, r_238__10_, r_238__9_, r_238__8_, r_238__7_, r_238__6_, r_238__5_, r_238__4_, r_238__3_, r_238__2_, r_238__1_, r_238__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N475)? data_i : 1'b0;
  assign N474 = sel_i[474];
  assign N475 = N2213;
  assign { r_n_238__63_, r_n_238__62_, r_n_238__61_, r_n_238__60_, r_n_238__59_, r_n_238__58_, r_n_238__57_, r_n_238__56_, r_n_238__55_, r_n_238__54_, r_n_238__53_, r_n_238__52_, r_n_238__51_, r_n_238__50_, r_n_238__49_, r_n_238__48_, r_n_238__47_, r_n_238__46_, r_n_238__45_, r_n_238__44_, r_n_238__43_, r_n_238__42_, r_n_238__41_, r_n_238__40_, r_n_238__39_, r_n_238__38_, r_n_238__37_, r_n_238__36_, r_n_238__35_, r_n_238__34_, r_n_238__33_, r_n_238__32_, r_n_238__31_, r_n_238__30_, r_n_238__29_, r_n_238__28_, r_n_238__27_, r_n_238__26_, r_n_238__25_, r_n_238__24_, r_n_238__23_, r_n_238__22_, r_n_238__21_, r_n_238__20_, r_n_238__19_, r_n_238__18_, r_n_238__17_, r_n_238__16_, r_n_238__15_, r_n_238__14_, r_n_238__13_, r_n_238__12_, r_n_238__11_, r_n_238__10_, r_n_238__9_, r_n_238__8_, r_n_238__7_, r_n_238__6_, r_n_238__5_, r_n_238__4_, r_n_238__3_, r_n_238__2_, r_n_238__1_, r_n_238__0_ } = (N476)? { r_239__63_, r_239__62_, r_239__61_, r_239__60_, r_239__59_, r_239__58_, r_239__57_, r_239__56_, r_239__55_, r_239__54_, r_239__53_, r_239__52_, r_239__51_, r_239__50_, r_239__49_, r_239__48_, r_239__47_, r_239__46_, r_239__45_, r_239__44_, r_239__43_, r_239__42_, r_239__41_, r_239__40_, r_239__39_, r_239__38_, r_239__37_, r_239__36_, r_239__35_, r_239__34_, r_239__33_, r_239__32_, r_239__31_, r_239__30_, r_239__29_, r_239__28_, r_239__27_, r_239__26_, r_239__25_, r_239__24_, r_239__23_, r_239__22_, r_239__21_, r_239__20_, r_239__19_, r_239__18_, r_239__17_, r_239__16_, r_239__15_, r_239__14_, r_239__13_, r_239__12_, r_239__11_, r_239__10_, r_239__9_, r_239__8_, r_239__7_, r_239__6_, r_239__5_, r_239__4_, r_239__3_, r_239__2_, r_239__1_, r_239__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N477)? data_i : 1'b0;
  assign N476 = sel_i[476];
  assign N477 = N2218;
  assign { r_n_239__63_, r_n_239__62_, r_n_239__61_, r_n_239__60_, r_n_239__59_, r_n_239__58_, r_n_239__57_, r_n_239__56_, r_n_239__55_, r_n_239__54_, r_n_239__53_, r_n_239__52_, r_n_239__51_, r_n_239__50_, r_n_239__49_, r_n_239__48_, r_n_239__47_, r_n_239__46_, r_n_239__45_, r_n_239__44_, r_n_239__43_, r_n_239__42_, r_n_239__41_, r_n_239__40_, r_n_239__39_, r_n_239__38_, r_n_239__37_, r_n_239__36_, r_n_239__35_, r_n_239__34_, r_n_239__33_, r_n_239__32_, r_n_239__31_, r_n_239__30_, r_n_239__29_, r_n_239__28_, r_n_239__27_, r_n_239__26_, r_n_239__25_, r_n_239__24_, r_n_239__23_, r_n_239__22_, r_n_239__21_, r_n_239__20_, r_n_239__19_, r_n_239__18_, r_n_239__17_, r_n_239__16_, r_n_239__15_, r_n_239__14_, r_n_239__13_, r_n_239__12_, r_n_239__11_, r_n_239__10_, r_n_239__9_, r_n_239__8_, r_n_239__7_, r_n_239__6_, r_n_239__5_, r_n_239__4_, r_n_239__3_, r_n_239__2_, r_n_239__1_, r_n_239__0_ } = (N478)? { r_240__63_, r_240__62_, r_240__61_, r_240__60_, r_240__59_, r_240__58_, r_240__57_, r_240__56_, r_240__55_, r_240__54_, r_240__53_, r_240__52_, r_240__51_, r_240__50_, r_240__49_, r_240__48_, r_240__47_, r_240__46_, r_240__45_, r_240__44_, r_240__43_, r_240__42_, r_240__41_, r_240__40_, r_240__39_, r_240__38_, r_240__37_, r_240__36_, r_240__35_, r_240__34_, r_240__33_, r_240__32_, r_240__31_, r_240__30_, r_240__29_, r_240__28_, r_240__27_, r_240__26_, r_240__25_, r_240__24_, r_240__23_, r_240__22_, r_240__21_, r_240__20_, r_240__19_, r_240__18_, r_240__17_, r_240__16_, r_240__15_, r_240__14_, r_240__13_, r_240__12_, r_240__11_, r_240__10_, r_240__9_, r_240__8_, r_240__7_, r_240__6_, r_240__5_, r_240__4_, r_240__3_, r_240__2_, r_240__1_, r_240__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N479)? data_i : 1'b0;
  assign N478 = sel_i[478];
  assign N479 = N2223;
  assign { r_n_240__63_, r_n_240__62_, r_n_240__61_, r_n_240__60_, r_n_240__59_, r_n_240__58_, r_n_240__57_, r_n_240__56_, r_n_240__55_, r_n_240__54_, r_n_240__53_, r_n_240__52_, r_n_240__51_, r_n_240__50_, r_n_240__49_, r_n_240__48_, r_n_240__47_, r_n_240__46_, r_n_240__45_, r_n_240__44_, r_n_240__43_, r_n_240__42_, r_n_240__41_, r_n_240__40_, r_n_240__39_, r_n_240__38_, r_n_240__37_, r_n_240__36_, r_n_240__35_, r_n_240__34_, r_n_240__33_, r_n_240__32_, r_n_240__31_, r_n_240__30_, r_n_240__29_, r_n_240__28_, r_n_240__27_, r_n_240__26_, r_n_240__25_, r_n_240__24_, r_n_240__23_, r_n_240__22_, r_n_240__21_, r_n_240__20_, r_n_240__19_, r_n_240__18_, r_n_240__17_, r_n_240__16_, r_n_240__15_, r_n_240__14_, r_n_240__13_, r_n_240__12_, r_n_240__11_, r_n_240__10_, r_n_240__9_, r_n_240__8_, r_n_240__7_, r_n_240__6_, r_n_240__5_, r_n_240__4_, r_n_240__3_, r_n_240__2_, r_n_240__1_, r_n_240__0_ } = (N480)? { r_241__63_, r_241__62_, r_241__61_, r_241__60_, r_241__59_, r_241__58_, r_241__57_, r_241__56_, r_241__55_, r_241__54_, r_241__53_, r_241__52_, r_241__51_, r_241__50_, r_241__49_, r_241__48_, r_241__47_, r_241__46_, r_241__45_, r_241__44_, r_241__43_, r_241__42_, r_241__41_, r_241__40_, r_241__39_, r_241__38_, r_241__37_, r_241__36_, r_241__35_, r_241__34_, r_241__33_, r_241__32_, r_241__31_, r_241__30_, r_241__29_, r_241__28_, r_241__27_, r_241__26_, r_241__25_, r_241__24_, r_241__23_, r_241__22_, r_241__21_, r_241__20_, r_241__19_, r_241__18_, r_241__17_, r_241__16_, r_241__15_, r_241__14_, r_241__13_, r_241__12_, r_241__11_, r_241__10_, r_241__9_, r_241__8_, r_241__7_, r_241__6_, r_241__5_, r_241__4_, r_241__3_, r_241__2_, r_241__1_, r_241__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N481)? data_i : 1'b0;
  assign N480 = sel_i[480];
  assign N481 = N2228;
  assign { r_n_241__63_, r_n_241__62_, r_n_241__61_, r_n_241__60_, r_n_241__59_, r_n_241__58_, r_n_241__57_, r_n_241__56_, r_n_241__55_, r_n_241__54_, r_n_241__53_, r_n_241__52_, r_n_241__51_, r_n_241__50_, r_n_241__49_, r_n_241__48_, r_n_241__47_, r_n_241__46_, r_n_241__45_, r_n_241__44_, r_n_241__43_, r_n_241__42_, r_n_241__41_, r_n_241__40_, r_n_241__39_, r_n_241__38_, r_n_241__37_, r_n_241__36_, r_n_241__35_, r_n_241__34_, r_n_241__33_, r_n_241__32_, r_n_241__31_, r_n_241__30_, r_n_241__29_, r_n_241__28_, r_n_241__27_, r_n_241__26_, r_n_241__25_, r_n_241__24_, r_n_241__23_, r_n_241__22_, r_n_241__21_, r_n_241__20_, r_n_241__19_, r_n_241__18_, r_n_241__17_, r_n_241__16_, r_n_241__15_, r_n_241__14_, r_n_241__13_, r_n_241__12_, r_n_241__11_, r_n_241__10_, r_n_241__9_, r_n_241__8_, r_n_241__7_, r_n_241__6_, r_n_241__5_, r_n_241__4_, r_n_241__3_, r_n_241__2_, r_n_241__1_, r_n_241__0_ } = (N482)? { r_242__63_, r_242__62_, r_242__61_, r_242__60_, r_242__59_, r_242__58_, r_242__57_, r_242__56_, r_242__55_, r_242__54_, r_242__53_, r_242__52_, r_242__51_, r_242__50_, r_242__49_, r_242__48_, r_242__47_, r_242__46_, r_242__45_, r_242__44_, r_242__43_, r_242__42_, r_242__41_, r_242__40_, r_242__39_, r_242__38_, r_242__37_, r_242__36_, r_242__35_, r_242__34_, r_242__33_, r_242__32_, r_242__31_, r_242__30_, r_242__29_, r_242__28_, r_242__27_, r_242__26_, r_242__25_, r_242__24_, r_242__23_, r_242__22_, r_242__21_, r_242__20_, r_242__19_, r_242__18_, r_242__17_, r_242__16_, r_242__15_, r_242__14_, r_242__13_, r_242__12_, r_242__11_, r_242__10_, r_242__9_, r_242__8_, r_242__7_, r_242__6_, r_242__5_, r_242__4_, r_242__3_, r_242__2_, r_242__1_, r_242__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N483)? data_i : 1'b0;
  assign N482 = sel_i[482];
  assign N483 = N2233;
  assign { r_n_242__63_, r_n_242__62_, r_n_242__61_, r_n_242__60_, r_n_242__59_, r_n_242__58_, r_n_242__57_, r_n_242__56_, r_n_242__55_, r_n_242__54_, r_n_242__53_, r_n_242__52_, r_n_242__51_, r_n_242__50_, r_n_242__49_, r_n_242__48_, r_n_242__47_, r_n_242__46_, r_n_242__45_, r_n_242__44_, r_n_242__43_, r_n_242__42_, r_n_242__41_, r_n_242__40_, r_n_242__39_, r_n_242__38_, r_n_242__37_, r_n_242__36_, r_n_242__35_, r_n_242__34_, r_n_242__33_, r_n_242__32_, r_n_242__31_, r_n_242__30_, r_n_242__29_, r_n_242__28_, r_n_242__27_, r_n_242__26_, r_n_242__25_, r_n_242__24_, r_n_242__23_, r_n_242__22_, r_n_242__21_, r_n_242__20_, r_n_242__19_, r_n_242__18_, r_n_242__17_, r_n_242__16_, r_n_242__15_, r_n_242__14_, r_n_242__13_, r_n_242__12_, r_n_242__11_, r_n_242__10_, r_n_242__9_, r_n_242__8_, r_n_242__7_, r_n_242__6_, r_n_242__5_, r_n_242__4_, r_n_242__3_, r_n_242__2_, r_n_242__1_, r_n_242__0_ } = (N484)? { r_243__63_, r_243__62_, r_243__61_, r_243__60_, r_243__59_, r_243__58_, r_243__57_, r_243__56_, r_243__55_, r_243__54_, r_243__53_, r_243__52_, r_243__51_, r_243__50_, r_243__49_, r_243__48_, r_243__47_, r_243__46_, r_243__45_, r_243__44_, r_243__43_, r_243__42_, r_243__41_, r_243__40_, r_243__39_, r_243__38_, r_243__37_, r_243__36_, r_243__35_, r_243__34_, r_243__33_, r_243__32_, r_243__31_, r_243__30_, r_243__29_, r_243__28_, r_243__27_, r_243__26_, r_243__25_, r_243__24_, r_243__23_, r_243__22_, r_243__21_, r_243__20_, r_243__19_, r_243__18_, r_243__17_, r_243__16_, r_243__15_, r_243__14_, r_243__13_, r_243__12_, r_243__11_, r_243__10_, r_243__9_, r_243__8_, r_243__7_, r_243__6_, r_243__5_, r_243__4_, r_243__3_, r_243__2_, r_243__1_, r_243__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N485)? data_i : 1'b0;
  assign N484 = sel_i[484];
  assign N485 = N2238;
  assign { r_n_243__63_, r_n_243__62_, r_n_243__61_, r_n_243__60_, r_n_243__59_, r_n_243__58_, r_n_243__57_, r_n_243__56_, r_n_243__55_, r_n_243__54_, r_n_243__53_, r_n_243__52_, r_n_243__51_, r_n_243__50_, r_n_243__49_, r_n_243__48_, r_n_243__47_, r_n_243__46_, r_n_243__45_, r_n_243__44_, r_n_243__43_, r_n_243__42_, r_n_243__41_, r_n_243__40_, r_n_243__39_, r_n_243__38_, r_n_243__37_, r_n_243__36_, r_n_243__35_, r_n_243__34_, r_n_243__33_, r_n_243__32_, r_n_243__31_, r_n_243__30_, r_n_243__29_, r_n_243__28_, r_n_243__27_, r_n_243__26_, r_n_243__25_, r_n_243__24_, r_n_243__23_, r_n_243__22_, r_n_243__21_, r_n_243__20_, r_n_243__19_, r_n_243__18_, r_n_243__17_, r_n_243__16_, r_n_243__15_, r_n_243__14_, r_n_243__13_, r_n_243__12_, r_n_243__11_, r_n_243__10_, r_n_243__9_, r_n_243__8_, r_n_243__7_, r_n_243__6_, r_n_243__5_, r_n_243__4_, r_n_243__3_, r_n_243__2_, r_n_243__1_, r_n_243__0_ } = (N486)? { r_244__63_, r_244__62_, r_244__61_, r_244__60_, r_244__59_, r_244__58_, r_244__57_, r_244__56_, r_244__55_, r_244__54_, r_244__53_, r_244__52_, r_244__51_, r_244__50_, r_244__49_, r_244__48_, r_244__47_, r_244__46_, r_244__45_, r_244__44_, r_244__43_, r_244__42_, r_244__41_, r_244__40_, r_244__39_, r_244__38_, r_244__37_, r_244__36_, r_244__35_, r_244__34_, r_244__33_, r_244__32_, r_244__31_, r_244__30_, r_244__29_, r_244__28_, r_244__27_, r_244__26_, r_244__25_, r_244__24_, r_244__23_, r_244__22_, r_244__21_, r_244__20_, r_244__19_, r_244__18_, r_244__17_, r_244__16_, r_244__15_, r_244__14_, r_244__13_, r_244__12_, r_244__11_, r_244__10_, r_244__9_, r_244__8_, r_244__7_, r_244__6_, r_244__5_, r_244__4_, r_244__3_, r_244__2_, r_244__1_, r_244__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N487)? data_i : 1'b0;
  assign N486 = sel_i[486];
  assign N487 = N2243;
  assign { r_n_244__63_, r_n_244__62_, r_n_244__61_, r_n_244__60_, r_n_244__59_, r_n_244__58_, r_n_244__57_, r_n_244__56_, r_n_244__55_, r_n_244__54_, r_n_244__53_, r_n_244__52_, r_n_244__51_, r_n_244__50_, r_n_244__49_, r_n_244__48_, r_n_244__47_, r_n_244__46_, r_n_244__45_, r_n_244__44_, r_n_244__43_, r_n_244__42_, r_n_244__41_, r_n_244__40_, r_n_244__39_, r_n_244__38_, r_n_244__37_, r_n_244__36_, r_n_244__35_, r_n_244__34_, r_n_244__33_, r_n_244__32_, r_n_244__31_, r_n_244__30_, r_n_244__29_, r_n_244__28_, r_n_244__27_, r_n_244__26_, r_n_244__25_, r_n_244__24_, r_n_244__23_, r_n_244__22_, r_n_244__21_, r_n_244__20_, r_n_244__19_, r_n_244__18_, r_n_244__17_, r_n_244__16_, r_n_244__15_, r_n_244__14_, r_n_244__13_, r_n_244__12_, r_n_244__11_, r_n_244__10_, r_n_244__9_, r_n_244__8_, r_n_244__7_, r_n_244__6_, r_n_244__5_, r_n_244__4_, r_n_244__3_, r_n_244__2_, r_n_244__1_, r_n_244__0_ } = (N488)? { r_245__63_, r_245__62_, r_245__61_, r_245__60_, r_245__59_, r_245__58_, r_245__57_, r_245__56_, r_245__55_, r_245__54_, r_245__53_, r_245__52_, r_245__51_, r_245__50_, r_245__49_, r_245__48_, r_245__47_, r_245__46_, r_245__45_, r_245__44_, r_245__43_, r_245__42_, r_245__41_, r_245__40_, r_245__39_, r_245__38_, r_245__37_, r_245__36_, r_245__35_, r_245__34_, r_245__33_, r_245__32_, r_245__31_, r_245__30_, r_245__29_, r_245__28_, r_245__27_, r_245__26_, r_245__25_, r_245__24_, r_245__23_, r_245__22_, r_245__21_, r_245__20_, r_245__19_, r_245__18_, r_245__17_, r_245__16_, r_245__15_, r_245__14_, r_245__13_, r_245__12_, r_245__11_, r_245__10_, r_245__9_, r_245__8_, r_245__7_, r_245__6_, r_245__5_, r_245__4_, r_245__3_, r_245__2_, r_245__1_, r_245__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N489)? data_i : 1'b0;
  assign N488 = sel_i[488];
  assign N489 = N2248;
  assign { r_n_245__63_, r_n_245__62_, r_n_245__61_, r_n_245__60_, r_n_245__59_, r_n_245__58_, r_n_245__57_, r_n_245__56_, r_n_245__55_, r_n_245__54_, r_n_245__53_, r_n_245__52_, r_n_245__51_, r_n_245__50_, r_n_245__49_, r_n_245__48_, r_n_245__47_, r_n_245__46_, r_n_245__45_, r_n_245__44_, r_n_245__43_, r_n_245__42_, r_n_245__41_, r_n_245__40_, r_n_245__39_, r_n_245__38_, r_n_245__37_, r_n_245__36_, r_n_245__35_, r_n_245__34_, r_n_245__33_, r_n_245__32_, r_n_245__31_, r_n_245__30_, r_n_245__29_, r_n_245__28_, r_n_245__27_, r_n_245__26_, r_n_245__25_, r_n_245__24_, r_n_245__23_, r_n_245__22_, r_n_245__21_, r_n_245__20_, r_n_245__19_, r_n_245__18_, r_n_245__17_, r_n_245__16_, r_n_245__15_, r_n_245__14_, r_n_245__13_, r_n_245__12_, r_n_245__11_, r_n_245__10_, r_n_245__9_, r_n_245__8_, r_n_245__7_, r_n_245__6_, r_n_245__5_, r_n_245__4_, r_n_245__3_, r_n_245__2_, r_n_245__1_, r_n_245__0_ } = (N490)? { r_246__63_, r_246__62_, r_246__61_, r_246__60_, r_246__59_, r_246__58_, r_246__57_, r_246__56_, r_246__55_, r_246__54_, r_246__53_, r_246__52_, r_246__51_, r_246__50_, r_246__49_, r_246__48_, r_246__47_, r_246__46_, r_246__45_, r_246__44_, r_246__43_, r_246__42_, r_246__41_, r_246__40_, r_246__39_, r_246__38_, r_246__37_, r_246__36_, r_246__35_, r_246__34_, r_246__33_, r_246__32_, r_246__31_, r_246__30_, r_246__29_, r_246__28_, r_246__27_, r_246__26_, r_246__25_, r_246__24_, r_246__23_, r_246__22_, r_246__21_, r_246__20_, r_246__19_, r_246__18_, r_246__17_, r_246__16_, r_246__15_, r_246__14_, r_246__13_, r_246__12_, r_246__11_, r_246__10_, r_246__9_, r_246__8_, r_246__7_, r_246__6_, r_246__5_, r_246__4_, r_246__3_, r_246__2_, r_246__1_, r_246__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N491)? data_i : 1'b0;
  assign N490 = sel_i[490];
  assign N491 = N2253;
  assign { r_n_246__63_, r_n_246__62_, r_n_246__61_, r_n_246__60_, r_n_246__59_, r_n_246__58_, r_n_246__57_, r_n_246__56_, r_n_246__55_, r_n_246__54_, r_n_246__53_, r_n_246__52_, r_n_246__51_, r_n_246__50_, r_n_246__49_, r_n_246__48_, r_n_246__47_, r_n_246__46_, r_n_246__45_, r_n_246__44_, r_n_246__43_, r_n_246__42_, r_n_246__41_, r_n_246__40_, r_n_246__39_, r_n_246__38_, r_n_246__37_, r_n_246__36_, r_n_246__35_, r_n_246__34_, r_n_246__33_, r_n_246__32_, r_n_246__31_, r_n_246__30_, r_n_246__29_, r_n_246__28_, r_n_246__27_, r_n_246__26_, r_n_246__25_, r_n_246__24_, r_n_246__23_, r_n_246__22_, r_n_246__21_, r_n_246__20_, r_n_246__19_, r_n_246__18_, r_n_246__17_, r_n_246__16_, r_n_246__15_, r_n_246__14_, r_n_246__13_, r_n_246__12_, r_n_246__11_, r_n_246__10_, r_n_246__9_, r_n_246__8_, r_n_246__7_, r_n_246__6_, r_n_246__5_, r_n_246__4_, r_n_246__3_, r_n_246__2_, r_n_246__1_, r_n_246__0_ } = (N492)? { r_247__63_, r_247__62_, r_247__61_, r_247__60_, r_247__59_, r_247__58_, r_247__57_, r_247__56_, r_247__55_, r_247__54_, r_247__53_, r_247__52_, r_247__51_, r_247__50_, r_247__49_, r_247__48_, r_247__47_, r_247__46_, r_247__45_, r_247__44_, r_247__43_, r_247__42_, r_247__41_, r_247__40_, r_247__39_, r_247__38_, r_247__37_, r_247__36_, r_247__35_, r_247__34_, r_247__33_, r_247__32_, r_247__31_, r_247__30_, r_247__29_, r_247__28_, r_247__27_, r_247__26_, r_247__25_, r_247__24_, r_247__23_, r_247__22_, r_247__21_, r_247__20_, r_247__19_, r_247__18_, r_247__17_, r_247__16_, r_247__15_, r_247__14_, r_247__13_, r_247__12_, r_247__11_, r_247__10_, r_247__9_, r_247__8_, r_247__7_, r_247__6_, r_247__5_, r_247__4_, r_247__3_, r_247__2_, r_247__1_, r_247__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N493)? data_i : 1'b0;
  assign N492 = sel_i[492];
  assign N493 = N2258;
  assign { r_n_247__63_, r_n_247__62_, r_n_247__61_, r_n_247__60_, r_n_247__59_, r_n_247__58_, r_n_247__57_, r_n_247__56_, r_n_247__55_, r_n_247__54_, r_n_247__53_, r_n_247__52_, r_n_247__51_, r_n_247__50_, r_n_247__49_, r_n_247__48_, r_n_247__47_, r_n_247__46_, r_n_247__45_, r_n_247__44_, r_n_247__43_, r_n_247__42_, r_n_247__41_, r_n_247__40_, r_n_247__39_, r_n_247__38_, r_n_247__37_, r_n_247__36_, r_n_247__35_, r_n_247__34_, r_n_247__33_, r_n_247__32_, r_n_247__31_, r_n_247__30_, r_n_247__29_, r_n_247__28_, r_n_247__27_, r_n_247__26_, r_n_247__25_, r_n_247__24_, r_n_247__23_, r_n_247__22_, r_n_247__21_, r_n_247__20_, r_n_247__19_, r_n_247__18_, r_n_247__17_, r_n_247__16_, r_n_247__15_, r_n_247__14_, r_n_247__13_, r_n_247__12_, r_n_247__11_, r_n_247__10_, r_n_247__9_, r_n_247__8_, r_n_247__7_, r_n_247__6_, r_n_247__5_, r_n_247__4_, r_n_247__3_, r_n_247__2_, r_n_247__1_, r_n_247__0_ } = (N494)? { r_248__63_, r_248__62_, r_248__61_, r_248__60_, r_248__59_, r_248__58_, r_248__57_, r_248__56_, r_248__55_, r_248__54_, r_248__53_, r_248__52_, r_248__51_, r_248__50_, r_248__49_, r_248__48_, r_248__47_, r_248__46_, r_248__45_, r_248__44_, r_248__43_, r_248__42_, r_248__41_, r_248__40_, r_248__39_, r_248__38_, r_248__37_, r_248__36_, r_248__35_, r_248__34_, r_248__33_, r_248__32_, r_248__31_, r_248__30_, r_248__29_, r_248__28_, r_248__27_, r_248__26_, r_248__25_, r_248__24_, r_248__23_, r_248__22_, r_248__21_, r_248__20_, r_248__19_, r_248__18_, r_248__17_, r_248__16_, r_248__15_, r_248__14_, r_248__13_, r_248__12_, r_248__11_, r_248__10_, r_248__9_, r_248__8_, r_248__7_, r_248__6_, r_248__5_, r_248__4_, r_248__3_, r_248__2_, r_248__1_, r_248__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N495)? data_i : 1'b0;
  assign N494 = sel_i[494];
  assign N495 = N2263;
  assign { r_n_248__63_, r_n_248__62_, r_n_248__61_, r_n_248__60_, r_n_248__59_, r_n_248__58_, r_n_248__57_, r_n_248__56_, r_n_248__55_, r_n_248__54_, r_n_248__53_, r_n_248__52_, r_n_248__51_, r_n_248__50_, r_n_248__49_, r_n_248__48_, r_n_248__47_, r_n_248__46_, r_n_248__45_, r_n_248__44_, r_n_248__43_, r_n_248__42_, r_n_248__41_, r_n_248__40_, r_n_248__39_, r_n_248__38_, r_n_248__37_, r_n_248__36_, r_n_248__35_, r_n_248__34_, r_n_248__33_, r_n_248__32_, r_n_248__31_, r_n_248__30_, r_n_248__29_, r_n_248__28_, r_n_248__27_, r_n_248__26_, r_n_248__25_, r_n_248__24_, r_n_248__23_, r_n_248__22_, r_n_248__21_, r_n_248__20_, r_n_248__19_, r_n_248__18_, r_n_248__17_, r_n_248__16_, r_n_248__15_, r_n_248__14_, r_n_248__13_, r_n_248__12_, r_n_248__11_, r_n_248__10_, r_n_248__9_, r_n_248__8_, r_n_248__7_, r_n_248__6_, r_n_248__5_, r_n_248__4_, r_n_248__3_, r_n_248__2_, r_n_248__1_, r_n_248__0_ } = (N496)? { r_249__63_, r_249__62_, r_249__61_, r_249__60_, r_249__59_, r_249__58_, r_249__57_, r_249__56_, r_249__55_, r_249__54_, r_249__53_, r_249__52_, r_249__51_, r_249__50_, r_249__49_, r_249__48_, r_249__47_, r_249__46_, r_249__45_, r_249__44_, r_249__43_, r_249__42_, r_249__41_, r_249__40_, r_249__39_, r_249__38_, r_249__37_, r_249__36_, r_249__35_, r_249__34_, r_249__33_, r_249__32_, r_249__31_, r_249__30_, r_249__29_, r_249__28_, r_249__27_, r_249__26_, r_249__25_, r_249__24_, r_249__23_, r_249__22_, r_249__21_, r_249__20_, r_249__19_, r_249__18_, r_249__17_, r_249__16_, r_249__15_, r_249__14_, r_249__13_, r_249__12_, r_249__11_, r_249__10_, r_249__9_, r_249__8_, r_249__7_, r_249__6_, r_249__5_, r_249__4_, r_249__3_, r_249__2_, r_249__1_, r_249__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N497)? data_i : 1'b0;
  assign N496 = sel_i[496];
  assign N497 = N2268;
  assign { r_n_249__63_, r_n_249__62_, r_n_249__61_, r_n_249__60_, r_n_249__59_, r_n_249__58_, r_n_249__57_, r_n_249__56_, r_n_249__55_, r_n_249__54_, r_n_249__53_, r_n_249__52_, r_n_249__51_, r_n_249__50_, r_n_249__49_, r_n_249__48_, r_n_249__47_, r_n_249__46_, r_n_249__45_, r_n_249__44_, r_n_249__43_, r_n_249__42_, r_n_249__41_, r_n_249__40_, r_n_249__39_, r_n_249__38_, r_n_249__37_, r_n_249__36_, r_n_249__35_, r_n_249__34_, r_n_249__33_, r_n_249__32_, r_n_249__31_, r_n_249__30_, r_n_249__29_, r_n_249__28_, r_n_249__27_, r_n_249__26_, r_n_249__25_, r_n_249__24_, r_n_249__23_, r_n_249__22_, r_n_249__21_, r_n_249__20_, r_n_249__19_, r_n_249__18_, r_n_249__17_, r_n_249__16_, r_n_249__15_, r_n_249__14_, r_n_249__13_, r_n_249__12_, r_n_249__11_, r_n_249__10_, r_n_249__9_, r_n_249__8_, r_n_249__7_, r_n_249__6_, r_n_249__5_, r_n_249__4_, r_n_249__3_, r_n_249__2_, r_n_249__1_, r_n_249__0_ } = (N498)? { r_250__63_, r_250__62_, r_250__61_, r_250__60_, r_250__59_, r_250__58_, r_250__57_, r_250__56_, r_250__55_, r_250__54_, r_250__53_, r_250__52_, r_250__51_, r_250__50_, r_250__49_, r_250__48_, r_250__47_, r_250__46_, r_250__45_, r_250__44_, r_250__43_, r_250__42_, r_250__41_, r_250__40_, r_250__39_, r_250__38_, r_250__37_, r_250__36_, r_250__35_, r_250__34_, r_250__33_, r_250__32_, r_250__31_, r_250__30_, r_250__29_, r_250__28_, r_250__27_, r_250__26_, r_250__25_, r_250__24_, r_250__23_, r_250__22_, r_250__21_, r_250__20_, r_250__19_, r_250__18_, r_250__17_, r_250__16_, r_250__15_, r_250__14_, r_250__13_, r_250__12_, r_250__11_, r_250__10_, r_250__9_, r_250__8_, r_250__7_, r_250__6_, r_250__5_, r_250__4_, r_250__3_, r_250__2_, r_250__1_, r_250__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N499)? data_i : 1'b0;
  assign N498 = sel_i[498];
  assign N499 = N2273;
  assign { r_n_250__63_, r_n_250__62_, r_n_250__61_, r_n_250__60_, r_n_250__59_, r_n_250__58_, r_n_250__57_, r_n_250__56_, r_n_250__55_, r_n_250__54_, r_n_250__53_, r_n_250__52_, r_n_250__51_, r_n_250__50_, r_n_250__49_, r_n_250__48_, r_n_250__47_, r_n_250__46_, r_n_250__45_, r_n_250__44_, r_n_250__43_, r_n_250__42_, r_n_250__41_, r_n_250__40_, r_n_250__39_, r_n_250__38_, r_n_250__37_, r_n_250__36_, r_n_250__35_, r_n_250__34_, r_n_250__33_, r_n_250__32_, r_n_250__31_, r_n_250__30_, r_n_250__29_, r_n_250__28_, r_n_250__27_, r_n_250__26_, r_n_250__25_, r_n_250__24_, r_n_250__23_, r_n_250__22_, r_n_250__21_, r_n_250__20_, r_n_250__19_, r_n_250__18_, r_n_250__17_, r_n_250__16_, r_n_250__15_, r_n_250__14_, r_n_250__13_, r_n_250__12_, r_n_250__11_, r_n_250__10_, r_n_250__9_, r_n_250__8_, r_n_250__7_, r_n_250__6_, r_n_250__5_, r_n_250__4_, r_n_250__3_, r_n_250__2_, r_n_250__1_, r_n_250__0_ } = (N500)? { r_251__63_, r_251__62_, r_251__61_, r_251__60_, r_251__59_, r_251__58_, r_251__57_, r_251__56_, r_251__55_, r_251__54_, r_251__53_, r_251__52_, r_251__51_, r_251__50_, r_251__49_, r_251__48_, r_251__47_, r_251__46_, r_251__45_, r_251__44_, r_251__43_, r_251__42_, r_251__41_, r_251__40_, r_251__39_, r_251__38_, r_251__37_, r_251__36_, r_251__35_, r_251__34_, r_251__33_, r_251__32_, r_251__31_, r_251__30_, r_251__29_, r_251__28_, r_251__27_, r_251__26_, r_251__25_, r_251__24_, r_251__23_, r_251__22_, r_251__21_, r_251__20_, r_251__19_, r_251__18_, r_251__17_, r_251__16_, r_251__15_, r_251__14_, r_251__13_, r_251__12_, r_251__11_, r_251__10_, r_251__9_, r_251__8_, r_251__7_, r_251__6_, r_251__5_, r_251__4_, r_251__3_, r_251__2_, r_251__1_, r_251__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N501)? data_i : 1'b0;
  assign N500 = sel_i[500];
  assign N501 = N2278;
  assign { r_n_251__63_, r_n_251__62_, r_n_251__61_, r_n_251__60_, r_n_251__59_, r_n_251__58_, r_n_251__57_, r_n_251__56_, r_n_251__55_, r_n_251__54_, r_n_251__53_, r_n_251__52_, r_n_251__51_, r_n_251__50_, r_n_251__49_, r_n_251__48_, r_n_251__47_, r_n_251__46_, r_n_251__45_, r_n_251__44_, r_n_251__43_, r_n_251__42_, r_n_251__41_, r_n_251__40_, r_n_251__39_, r_n_251__38_, r_n_251__37_, r_n_251__36_, r_n_251__35_, r_n_251__34_, r_n_251__33_, r_n_251__32_, r_n_251__31_, r_n_251__30_, r_n_251__29_, r_n_251__28_, r_n_251__27_, r_n_251__26_, r_n_251__25_, r_n_251__24_, r_n_251__23_, r_n_251__22_, r_n_251__21_, r_n_251__20_, r_n_251__19_, r_n_251__18_, r_n_251__17_, r_n_251__16_, r_n_251__15_, r_n_251__14_, r_n_251__13_, r_n_251__12_, r_n_251__11_, r_n_251__10_, r_n_251__9_, r_n_251__8_, r_n_251__7_, r_n_251__6_, r_n_251__5_, r_n_251__4_, r_n_251__3_, r_n_251__2_, r_n_251__1_, r_n_251__0_ } = (N502)? { r_252__63_, r_252__62_, r_252__61_, r_252__60_, r_252__59_, r_252__58_, r_252__57_, r_252__56_, r_252__55_, r_252__54_, r_252__53_, r_252__52_, r_252__51_, r_252__50_, r_252__49_, r_252__48_, r_252__47_, r_252__46_, r_252__45_, r_252__44_, r_252__43_, r_252__42_, r_252__41_, r_252__40_, r_252__39_, r_252__38_, r_252__37_, r_252__36_, r_252__35_, r_252__34_, r_252__33_, r_252__32_, r_252__31_, r_252__30_, r_252__29_, r_252__28_, r_252__27_, r_252__26_, r_252__25_, r_252__24_, r_252__23_, r_252__22_, r_252__21_, r_252__20_, r_252__19_, r_252__18_, r_252__17_, r_252__16_, r_252__15_, r_252__14_, r_252__13_, r_252__12_, r_252__11_, r_252__10_, r_252__9_, r_252__8_, r_252__7_, r_252__6_, r_252__5_, r_252__4_, r_252__3_, r_252__2_, r_252__1_, r_252__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N503)? data_i : 1'b0;
  assign N502 = sel_i[502];
  assign N503 = N2283;
  assign { r_n_252__63_, r_n_252__62_, r_n_252__61_, r_n_252__60_, r_n_252__59_, r_n_252__58_, r_n_252__57_, r_n_252__56_, r_n_252__55_, r_n_252__54_, r_n_252__53_, r_n_252__52_, r_n_252__51_, r_n_252__50_, r_n_252__49_, r_n_252__48_, r_n_252__47_, r_n_252__46_, r_n_252__45_, r_n_252__44_, r_n_252__43_, r_n_252__42_, r_n_252__41_, r_n_252__40_, r_n_252__39_, r_n_252__38_, r_n_252__37_, r_n_252__36_, r_n_252__35_, r_n_252__34_, r_n_252__33_, r_n_252__32_, r_n_252__31_, r_n_252__30_, r_n_252__29_, r_n_252__28_, r_n_252__27_, r_n_252__26_, r_n_252__25_, r_n_252__24_, r_n_252__23_, r_n_252__22_, r_n_252__21_, r_n_252__20_, r_n_252__19_, r_n_252__18_, r_n_252__17_, r_n_252__16_, r_n_252__15_, r_n_252__14_, r_n_252__13_, r_n_252__12_, r_n_252__11_, r_n_252__10_, r_n_252__9_, r_n_252__8_, r_n_252__7_, r_n_252__6_, r_n_252__5_, r_n_252__4_, r_n_252__3_, r_n_252__2_, r_n_252__1_, r_n_252__0_ } = (N504)? { r_253__63_, r_253__62_, r_253__61_, r_253__60_, r_253__59_, r_253__58_, r_253__57_, r_253__56_, r_253__55_, r_253__54_, r_253__53_, r_253__52_, r_253__51_, r_253__50_, r_253__49_, r_253__48_, r_253__47_, r_253__46_, r_253__45_, r_253__44_, r_253__43_, r_253__42_, r_253__41_, r_253__40_, r_253__39_, r_253__38_, r_253__37_, r_253__36_, r_253__35_, r_253__34_, r_253__33_, r_253__32_, r_253__31_, r_253__30_, r_253__29_, r_253__28_, r_253__27_, r_253__26_, r_253__25_, r_253__24_, r_253__23_, r_253__22_, r_253__21_, r_253__20_, r_253__19_, r_253__18_, r_253__17_, r_253__16_, r_253__15_, r_253__14_, r_253__13_, r_253__12_, r_253__11_, r_253__10_, r_253__9_, r_253__8_, r_253__7_, r_253__6_, r_253__5_, r_253__4_, r_253__3_, r_253__2_, r_253__1_, r_253__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N505)? data_i : 1'b0;
  assign N504 = sel_i[504];
  assign N505 = N2288;
  assign { r_n_253__63_, r_n_253__62_, r_n_253__61_, r_n_253__60_, r_n_253__59_, r_n_253__58_, r_n_253__57_, r_n_253__56_, r_n_253__55_, r_n_253__54_, r_n_253__53_, r_n_253__52_, r_n_253__51_, r_n_253__50_, r_n_253__49_, r_n_253__48_, r_n_253__47_, r_n_253__46_, r_n_253__45_, r_n_253__44_, r_n_253__43_, r_n_253__42_, r_n_253__41_, r_n_253__40_, r_n_253__39_, r_n_253__38_, r_n_253__37_, r_n_253__36_, r_n_253__35_, r_n_253__34_, r_n_253__33_, r_n_253__32_, r_n_253__31_, r_n_253__30_, r_n_253__29_, r_n_253__28_, r_n_253__27_, r_n_253__26_, r_n_253__25_, r_n_253__24_, r_n_253__23_, r_n_253__22_, r_n_253__21_, r_n_253__20_, r_n_253__19_, r_n_253__18_, r_n_253__17_, r_n_253__16_, r_n_253__15_, r_n_253__14_, r_n_253__13_, r_n_253__12_, r_n_253__11_, r_n_253__10_, r_n_253__9_, r_n_253__8_, r_n_253__7_, r_n_253__6_, r_n_253__5_, r_n_253__4_, r_n_253__3_, r_n_253__2_, r_n_253__1_, r_n_253__0_ } = (N506)? { r_254__63_, r_254__62_, r_254__61_, r_254__60_, r_254__59_, r_254__58_, r_254__57_, r_254__56_, r_254__55_, r_254__54_, r_254__53_, r_254__52_, r_254__51_, r_254__50_, r_254__49_, r_254__48_, r_254__47_, r_254__46_, r_254__45_, r_254__44_, r_254__43_, r_254__42_, r_254__41_, r_254__40_, r_254__39_, r_254__38_, r_254__37_, r_254__36_, r_254__35_, r_254__34_, r_254__33_, r_254__32_, r_254__31_, r_254__30_, r_254__29_, r_254__28_, r_254__27_, r_254__26_, r_254__25_, r_254__24_, r_254__23_, r_254__22_, r_254__21_, r_254__20_, r_254__19_, r_254__18_, r_254__17_, r_254__16_, r_254__15_, r_254__14_, r_254__13_, r_254__12_, r_254__11_, r_254__10_, r_254__9_, r_254__8_, r_254__7_, r_254__6_, r_254__5_, r_254__4_, r_254__3_, r_254__2_, r_254__1_, r_254__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N507)? data_i : 1'b0;
  assign N506 = sel_i[506];
  assign N507 = N2293;
  assign { r_n_254__63_, r_n_254__62_, r_n_254__61_, r_n_254__60_, r_n_254__59_, r_n_254__58_, r_n_254__57_, r_n_254__56_, r_n_254__55_, r_n_254__54_, r_n_254__53_, r_n_254__52_, r_n_254__51_, r_n_254__50_, r_n_254__49_, r_n_254__48_, r_n_254__47_, r_n_254__46_, r_n_254__45_, r_n_254__44_, r_n_254__43_, r_n_254__42_, r_n_254__41_, r_n_254__40_, r_n_254__39_, r_n_254__38_, r_n_254__37_, r_n_254__36_, r_n_254__35_, r_n_254__34_, r_n_254__33_, r_n_254__32_, r_n_254__31_, r_n_254__30_, r_n_254__29_, r_n_254__28_, r_n_254__27_, r_n_254__26_, r_n_254__25_, r_n_254__24_, r_n_254__23_, r_n_254__22_, r_n_254__21_, r_n_254__20_, r_n_254__19_, r_n_254__18_, r_n_254__17_, r_n_254__16_, r_n_254__15_, r_n_254__14_, r_n_254__13_, r_n_254__12_, r_n_254__11_, r_n_254__10_, r_n_254__9_, r_n_254__8_, r_n_254__7_, r_n_254__6_, r_n_254__5_, r_n_254__4_, r_n_254__3_, r_n_254__2_, r_n_254__1_, r_n_254__0_ } = (N508)? { r_255__63_, r_255__62_, r_255__61_, r_255__60_, r_255__59_, r_255__58_, r_255__57_, r_255__56_, r_255__55_, r_255__54_, r_255__53_, r_255__52_, r_255__51_, r_255__50_, r_255__49_, r_255__48_, r_255__47_, r_255__46_, r_255__45_, r_255__44_, r_255__43_, r_255__42_, r_255__41_, r_255__40_, r_255__39_, r_255__38_, r_255__37_, r_255__36_, r_255__35_, r_255__34_, r_255__33_, r_255__32_, r_255__31_, r_255__30_, r_255__29_, r_255__28_, r_255__27_, r_255__26_, r_255__25_, r_255__24_, r_255__23_, r_255__22_, r_255__21_, r_255__20_, r_255__19_, r_255__18_, r_255__17_, r_255__16_, r_255__15_, r_255__14_, r_255__13_, r_255__12_, r_255__11_, r_255__10_, r_255__9_, r_255__8_, r_255__7_, r_255__6_, r_255__5_, r_255__4_, r_255__3_, r_255__2_, r_255__1_, r_255__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N509)? data_i : 1'b0;
  assign N508 = sel_i[508];
  assign N509 = N2298;
  assign { r_n_255__63_, r_n_255__62_, r_n_255__61_, r_n_255__60_, r_n_255__59_, r_n_255__58_, r_n_255__57_, r_n_255__56_, r_n_255__55_, r_n_255__54_, r_n_255__53_, r_n_255__52_, r_n_255__51_, r_n_255__50_, r_n_255__49_, r_n_255__48_, r_n_255__47_, r_n_255__46_, r_n_255__45_, r_n_255__44_, r_n_255__43_, r_n_255__42_, r_n_255__41_, r_n_255__40_, r_n_255__39_, r_n_255__38_, r_n_255__37_, r_n_255__36_, r_n_255__35_, r_n_255__34_, r_n_255__33_, r_n_255__32_, r_n_255__31_, r_n_255__30_, r_n_255__29_, r_n_255__28_, r_n_255__27_, r_n_255__26_, r_n_255__25_, r_n_255__24_, r_n_255__23_, r_n_255__22_, r_n_255__21_, r_n_255__20_, r_n_255__19_, r_n_255__18_, r_n_255__17_, r_n_255__16_, r_n_255__15_, r_n_255__14_, r_n_255__13_, r_n_255__12_, r_n_255__11_, r_n_255__10_, r_n_255__9_, r_n_255__8_, r_n_255__7_, r_n_255__6_, r_n_255__5_, r_n_255__4_, r_n_255__3_, r_n_255__2_, r_n_255__1_, r_n_255__0_ } = (N510)? { r_256__63_, r_256__62_, r_256__61_, r_256__60_, r_256__59_, r_256__58_, r_256__57_, r_256__56_, r_256__55_, r_256__54_, r_256__53_, r_256__52_, r_256__51_, r_256__50_, r_256__49_, r_256__48_, r_256__47_, r_256__46_, r_256__45_, r_256__44_, r_256__43_, r_256__42_, r_256__41_, r_256__40_, r_256__39_, r_256__38_, r_256__37_, r_256__36_, r_256__35_, r_256__34_, r_256__33_, r_256__32_, r_256__31_, r_256__30_, r_256__29_, r_256__28_, r_256__27_, r_256__26_, r_256__25_, r_256__24_, r_256__23_, r_256__22_, r_256__21_, r_256__20_, r_256__19_, r_256__18_, r_256__17_, r_256__16_, r_256__15_, r_256__14_, r_256__13_, r_256__12_, r_256__11_, r_256__10_, r_256__9_, r_256__8_, r_256__7_, r_256__6_, r_256__5_, r_256__4_, r_256__3_, r_256__2_, r_256__1_, r_256__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N511)? data_i : 1'b0;
  assign N510 = sel_i[510];
  assign N511 = N2303;
  assign { r_n_256__63_, r_n_256__62_, r_n_256__61_, r_n_256__60_, r_n_256__59_, r_n_256__58_, r_n_256__57_, r_n_256__56_, r_n_256__55_, r_n_256__54_, r_n_256__53_, r_n_256__52_, r_n_256__51_, r_n_256__50_, r_n_256__49_, r_n_256__48_, r_n_256__47_, r_n_256__46_, r_n_256__45_, r_n_256__44_, r_n_256__43_, r_n_256__42_, r_n_256__41_, r_n_256__40_, r_n_256__39_, r_n_256__38_, r_n_256__37_, r_n_256__36_, r_n_256__35_, r_n_256__34_, r_n_256__33_, r_n_256__32_, r_n_256__31_, r_n_256__30_, r_n_256__29_, r_n_256__28_, r_n_256__27_, r_n_256__26_, r_n_256__25_, r_n_256__24_, r_n_256__23_, r_n_256__22_, r_n_256__21_, r_n_256__20_, r_n_256__19_, r_n_256__18_, r_n_256__17_, r_n_256__16_, r_n_256__15_, r_n_256__14_, r_n_256__13_, r_n_256__12_, r_n_256__11_, r_n_256__10_, r_n_256__9_, r_n_256__8_, r_n_256__7_, r_n_256__6_, r_n_256__5_, r_n_256__4_, r_n_256__3_, r_n_256__2_, r_n_256__1_, r_n_256__0_ } = (N512)? { r_257__63_, r_257__62_, r_257__61_, r_257__60_, r_257__59_, r_257__58_, r_257__57_, r_257__56_, r_257__55_, r_257__54_, r_257__53_, r_257__52_, r_257__51_, r_257__50_, r_257__49_, r_257__48_, r_257__47_, r_257__46_, r_257__45_, r_257__44_, r_257__43_, r_257__42_, r_257__41_, r_257__40_, r_257__39_, r_257__38_, r_257__37_, r_257__36_, r_257__35_, r_257__34_, r_257__33_, r_257__32_, r_257__31_, r_257__30_, r_257__29_, r_257__28_, r_257__27_, r_257__26_, r_257__25_, r_257__24_, r_257__23_, r_257__22_, r_257__21_, r_257__20_, r_257__19_, r_257__18_, r_257__17_, r_257__16_, r_257__15_, r_257__14_, r_257__13_, r_257__12_, r_257__11_, r_257__10_, r_257__9_, r_257__8_, r_257__7_, r_257__6_, r_257__5_, r_257__4_, r_257__3_, r_257__2_, r_257__1_, r_257__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N513)? data_i : 1'b0;
  assign N512 = sel_i[512];
  assign N513 = N2308;
  assign { r_n_257__63_, r_n_257__62_, r_n_257__61_, r_n_257__60_, r_n_257__59_, r_n_257__58_, r_n_257__57_, r_n_257__56_, r_n_257__55_, r_n_257__54_, r_n_257__53_, r_n_257__52_, r_n_257__51_, r_n_257__50_, r_n_257__49_, r_n_257__48_, r_n_257__47_, r_n_257__46_, r_n_257__45_, r_n_257__44_, r_n_257__43_, r_n_257__42_, r_n_257__41_, r_n_257__40_, r_n_257__39_, r_n_257__38_, r_n_257__37_, r_n_257__36_, r_n_257__35_, r_n_257__34_, r_n_257__33_, r_n_257__32_, r_n_257__31_, r_n_257__30_, r_n_257__29_, r_n_257__28_, r_n_257__27_, r_n_257__26_, r_n_257__25_, r_n_257__24_, r_n_257__23_, r_n_257__22_, r_n_257__21_, r_n_257__20_, r_n_257__19_, r_n_257__18_, r_n_257__17_, r_n_257__16_, r_n_257__15_, r_n_257__14_, r_n_257__13_, r_n_257__12_, r_n_257__11_, r_n_257__10_, r_n_257__9_, r_n_257__8_, r_n_257__7_, r_n_257__6_, r_n_257__5_, r_n_257__4_, r_n_257__3_, r_n_257__2_, r_n_257__1_, r_n_257__0_ } = (N514)? { r_258__63_, r_258__62_, r_258__61_, r_258__60_, r_258__59_, r_258__58_, r_258__57_, r_258__56_, r_258__55_, r_258__54_, r_258__53_, r_258__52_, r_258__51_, r_258__50_, r_258__49_, r_258__48_, r_258__47_, r_258__46_, r_258__45_, r_258__44_, r_258__43_, r_258__42_, r_258__41_, r_258__40_, r_258__39_, r_258__38_, r_258__37_, r_258__36_, r_258__35_, r_258__34_, r_258__33_, r_258__32_, r_258__31_, r_258__30_, r_258__29_, r_258__28_, r_258__27_, r_258__26_, r_258__25_, r_258__24_, r_258__23_, r_258__22_, r_258__21_, r_258__20_, r_258__19_, r_258__18_, r_258__17_, r_258__16_, r_258__15_, r_258__14_, r_258__13_, r_258__12_, r_258__11_, r_258__10_, r_258__9_, r_258__8_, r_258__7_, r_258__6_, r_258__5_, r_258__4_, r_258__3_, r_258__2_, r_258__1_, r_258__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N515)? data_i : 1'b0;
  assign N514 = sel_i[514];
  assign N515 = N2313;
  assign { r_n_258__63_, r_n_258__62_, r_n_258__61_, r_n_258__60_, r_n_258__59_, r_n_258__58_, r_n_258__57_, r_n_258__56_, r_n_258__55_, r_n_258__54_, r_n_258__53_, r_n_258__52_, r_n_258__51_, r_n_258__50_, r_n_258__49_, r_n_258__48_, r_n_258__47_, r_n_258__46_, r_n_258__45_, r_n_258__44_, r_n_258__43_, r_n_258__42_, r_n_258__41_, r_n_258__40_, r_n_258__39_, r_n_258__38_, r_n_258__37_, r_n_258__36_, r_n_258__35_, r_n_258__34_, r_n_258__33_, r_n_258__32_, r_n_258__31_, r_n_258__30_, r_n_258__29_, r_n_258__28_, r_n_258__27_, r_n_258__26_, r_n_258__25_, r_n_258__24_, r_n_258__23_, r_n_258__22_, r_n_258__21_, r_n_258__20_, r_n_258__19_, r_n_258__18_, r_n_258__17_, r_n_258__16_, r_n_258__15_, r_n_258__14_, r_n_258__13_, r_n_258__12_, r_n_258__11_, r_n_258__10_, r_n_258__9_, r_n_258__8_, r_n_258__7_, r_n_258__6_, r_n_258__5_, r_n_258__4_, r_n_258__3_, r_n_258__2_, r_n_258__1_, r_n_258__0_ } = (N516)? { r_259__63_, r_259__62_, r_259__61_, r_259__60_, r_259__59_, r_259__58_, r_259__57_, r_259__56_, r_259__55_, r_259__54_, r_259__53_, r_259__52_, r_259__51_, r_259__50_, r_259__49_, r_259__48_, r_259__47_, r_259__46_, r_259__45_, r_259__44_, r_259__43_, r_259__42_, r_259__41_, r_259__40_, r_259__39_, r_259__38_, r_259__37_, r_259__36_, r_259__35_, r_259__34_, r_259__33_, r_259__32_, r_259__31_, r_259__30_, r_259__29_, r_259__28_, r_259__27_, r_259__26_, r_259__25_, r_259__24_, r_259__23_, r_259__22_, r_259__21_, r_259__20_, r_259__19_, r_259__18_, r_259__17_, r_259__16_, r_259__15_, r_259__14_, r_259__13_, r_259__12_, r_259__11_, r_259__10_, r_259__9_, r_259__8_, r_259__7_, r_259__6_, r_259__5_, r_259__4_, r_259__3_, r_259__2_, r_259__1_, r_259__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N517)? data_i : 1'b0;
  assign N516 = sel_i[516];
  assign N517 = N2318;
  assign { r_n_259__63_, r_n_259__62_, r_n_259__61_, r_n_259__60_, r_n_259__59_, r_n_259__58_, r_n_259__57_, r_n_259__56_, r_n_259__55_, r_n_259__54_, r_n_259__53_, r_n_259__52_, r_n_259__51_, r_n_259__50_, r_n_259__49_, r_n_259__48_, r_n_259__47_, r_n_259__46_, r_n_259__45_, r_n_259__44_, r_n_259__43_, r_n_259__42_, r_n_259__41_, r_n_259__40_, r_n_259__39_, r_n_259__38_, r_n_259__37_, r_n_259__36_, r_n_259__35_, r_n_259__34_, r_n_259__33_, r_n_259__32_, r_n_259__31_, r_n_259__30_, r_n_259__29_, r_n_259__28_, r_n_259__27_, r_n_259__26_, r_n_259__25_, r_n_259__24_, r_n_259__23_, r_n_259__22_, r_n_259__21_, r_n_259__20_, r_n_259__19_, r_n_259__18_, r_n_259__17_, r_n_259__16_, r_n_259__15_, r_n_259__14_, r_n_259__13_, r_n_259__12_, r_n_259__11_, r_n_259__10_, r_n_259__9_, r_n_259__8_, r_n_259__7_, r_n_259__6_, r_n_259__5_, r_n_259__4_, r_n_259__3_, r_n_259__2_, r_n_259__1_, r_n_259__0_ } = (N518)? { r_260__63_, r_260__62_, r_260__61_, r_260__60_, r_260__59_, r_260__58_, r_260__57_, r_260__56_, r_260__55_, r_260__54_, r_260__53_, r_260__52_, r_260__51_, r_260__50_, r_260__49_, r_260__48_, r_260__47_, r_260__46_, r_260__45_, r_260__44_, r_260__43_, r_260__42_, r_260__41_, r_260__40_, r_260__39_, r_260__38_, r_260__37_, r_260__36_, r_260__35_, r_260__34_, r_260__33_, r_260__32_, r_260__31_, r_260__30_, r_260__29_, r_260__28_, r_260__27_, r_260__26_, r_260__25_, r_260__24_, r_260__23_, r_260__22_, r_260__21_, r_260__20_, r_260__19_, r_260__18_, r_260__17_, r_260__16_, r_260__15_, r_260__14_, r_260__13_, r_260__12_, r_260__11_, r_260__10_, r_260__9_, r_260__8_, r_260__7_, r_260__6_, r_260__5_, r_260__4_, r_260__3_, r_260__2_, r_260__1_, r_260__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N519)? data_i : 1'b0;
  assign N518 = sel_i[518];
  assign N519 = N2323;
  assign { r_n_260__63_, r_n_260__62_, r_n_260__61_, r_n_260__60_, r_n_260__59_, r_n_260__58_, r_n_260__57_, r_n_260__56_, r_n_260__55_, r_n_260__54_, r_n_260__53_, r_n_260__52_, r_n_260__51_, r_n_260__50_, r_n_260__49_, r_n_260__48_, r_n_260__47_, r_n_260__46_, r_n_260__45_, r_n_260__44_, r_n_260__43_, r_n_260__42_, r_n_260__41_, r_n_260__40_, r_n_260__39_, r_n_260__38_, r_n_260__37_, r_n_260__36_, r_n_260__35_, r_n_260__34_, r_n_260__33_, r_n_260__32_, r_n_260__31_, r_n_260__30_, r_n_260__29_, r_n_260__28_, r_n_260__27_, r_n_260__26_, r_n_260__25_, r_n_260__24_, r_n_260__23_, r_n_260__22_, r_n_260__21_, r_n_260__20_, r_n_260__19_, r_n_260__18_, r_n_260__17_, r_n_260__16_, r_n_260__15_, r_n_260__14_, r_n_260__13_, r_n_260__12_, r_n_260__11_, r_n_260__10_, r_n_260__9_, r_n_260__8_, r_n_260__7_, r_n_260__6_, r_n_260__5_, r_n_260__4_, r_n_260__3_, r_n_260__2_, r_n_260__1_, r_n_260__0_ } = (N520)? { r_261__63_, r_261__62_, r_261__61_, r_261__60_, r_261__59_, r_261__58_, r_261__57_, r_261__56_, r_261__55_, r_261__54_, r_261__53_, r_261__52_, r_261__51_, r_261__50_, r_261__49_, r_261__48_, r_261__47_, r_261__46_, r_261__45_, r_261__44_, r_261__43_, r_261__42_, r_261__41_, r_261__40_, r_261__39_, r_261__38_, r_261__37_, r_261__36_, r_261__35_, r_261__34_, r_261__33_, r_261__32_, r_261__31_, r_261__30_, r_261__29_, r_261__28_, r_261__27_, r_261__26_, r_261__25_, r_261__24_, r_261__23_, r_261__22_, r_261__21_, r_261__20_, r_261__19_, r_261__18_, r_261__17_, r_261__16_, r_261__15_, r_261__14_, r_261__13_, r_261__12_, r_261__11_, r_261__10_, r_261__9_, r_261__8_, r_261__7_, r_261__6_, r_261__5_, r_261__4_, r_261__3_, r_261__2_, r_261__1_, r_261__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N521)? data_i : 1'b0;
  assign N520 = sel_i[520];
  assign N521 = N2328;
  assign { r_n_261__63_, r_n_261__62_, r_n_261__61_, r_n_261__60_, r_n_261__59_, r_n_261__58_, r_n_261__57_, r_n_261__56_, r_n_261__55_, r_n_261__54_, r_n_261__53_, r_n_261__52_, r_n_261__51_, r_n_261__50_, r_n_261__49_, r_n_261__48_, r_n_261__47_, r_n_261__46_, r_n_261__45_, r_n_261__44_, r_n_261__43_, r_n_261__42_, r_n_261__41_, r_n_261__40_, r_n_261__39_, r_n_261__38_, r_n_261__37_, r_n_261__36_, r_n_261__35_, r_n_261__34_, r_n_261__33_, r_n_261__32_, r_n_261__31_, r_n_261__30_, r_n_261__29_, r_n_261__28_, r_n_261__27_, r_n_261__26_, r_n_261__25_, r_n_261__24_, r_n_261__23_, r_n_261__22_, r_n_261__21_, r_n_261__20_, r_n_261__19_, r_n_261__18_, r_n_261__17_, r_n_261__16_, r_n_261__15_, r_n_261__14_, r_n_261__13_, r_n_261__12_, r_n_261__11_, r_n_261__10_, r_n_261__9_, r_n_261__8_, r_n_261__7_, r_n_261__6_, r_n_261__5_, r_n_261__4_, r_n_261__3_, r_n_261__2_, r_n_261__1_, r_n_261__0_ } = (N522)? { r_262__63_, r_262__62_, r_262__61_, r_262__60_, r_262__59_, r_262__58_, r_262__57_, r_262__56_, r_262__55_, r_262__54_, r_262__53_, r_262__52_, r_262__51_, r_262__50_, r_262__49_, r_262__48_, r_262__47_, r_262__46_, r_262__45_, r_262__44_, r_262__43_, r_262__42_, r_262__41_, r_262__40_, r_262__39_, r_262__38_, r_262__37_, r_262__36_, r_262__35_, r_262__34_, r_262__33_, r_262__32_, r_262__31_, r_262__30_, r_262__29_, r_262__28_, r_262__27_, r_262__26_, r_262__25_, r_262__24_, r_262__23_, r_262__22_, r_262__21_, r_262__20_, r_262__19_, r_262__18_, r_262__17_, r_262__16_, r_262__15_, r_262__14_, r_262__13_, r_262__12_, r_262__11_, r_262__10_, r_262__9_, r_262__8_, r_262__7_, r_262__6_, r_262__5_, r_262__4_, r_262__3_, r_262__2_, r_262__1_, r_262__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N523)? data_i : 1'b0;
  assign N522 = sel_i[522];
  assign N523 = N2333;
  assign { r_n_262__63_, r_n_262__62_, r_n_262__61_, r_n_262__60_, r_n_262__59_, r_n_262__58_, r_n_262__57_, r_n_262__56_, r_n_262__55_, r_n_262__54_, r_n_262__53_, r_n_262__52_, r_n_262__51_, r_n_262__50_, r_n_262__49_, r_n_262__48_, r_n_262__47_, r_n_262__46_, r_n_262__45_, r_n_262__44_, r_n_262__43_, r_n_262__42_, r_n_262__41_, r_n_262__40_, r_n_262__39_, r_n_262__38_, r_n_262__37_, r_n_262__36_, r_n_262__35_, r_n_262__34_, r_n_262__33_, r_n_262__32_, r_n_262__31_, r_n_262__30_, r_n_262__29_, r_n_262__28_, r_n_262__27_, r_n_262__26_, r_n_262__25_, r_n_262__24_, r_n_262__23_, r_n_262__22_, r_n_262__21_, r_n_262__20_, r_n_262__19_, r_n_262__18_, r_n_262__17_, r_n_262__16_, r_n_262__15_, r_n_262__14_, r_n_262__13_, r_n_262__12_, r_n_262__11_, r_n_262__10_, r_n_262__9_, r_n_262__8_, r_n_262__7_, r_n_262__6_, r_n_262__5_, r_n_262__4_, r_n_262__3_, r_n_262__2_, r_n_262__1_, r_n_262__0_ } = (N524)? { r_263__63_, r_263__62_, r_263__61_, r_263__60_, r_263__59_, r_263__58_, r_263__57_, r_263__56_, r_263__55_, r_263__54_, r_263__53_, r_263__52_, r_263__51_, r_263__50_, r_263__49_, r_263__48_, r_263__47_, r_263__46_, r_263__45_, r_263__44_, r_263__43_, r_263__42_, r_263__41_, r_263__40_, r_263__39_, r_263__38_, r_263__37_, r_263__36_, r_263__35_, r_263__34_, r_263__33_, r_263__32_, r_263__31_, r_263__30_, r_263__29_, r_263__28_, r_263__27_, r_263__26_, r_263__25_, r_263__24_, r_263__23_, r_263__22_, r_263__21_, r_263__20_, r_263__19_, r_263__18_, r_263__17_, r_263__16_, r_263__15_, r_263__14_, r_263__13_, r_263__12_, r_263__11_, r_263__10_, r_263__9_, r_263__8_, r_263__7_, r_263__6_, r_263__5_, r_263__4_, r_263__3_, r_263__2_, r_263__1_, r_263__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N525)? data_i : 1'b0;
  assign N524 = sel_i[524];
  assign N525 = N2338;
  assign { r_n_263__63_, r_n_263__62_, r_n_263__61_, r_n_263__60_, r_n_263__59_, r_n_263__58_, r_n_263__57_, r_n_263__56_, r_n_263__55_, r_n_263__54_, r_n_263__53_, r_n_263__52_, r_n_263__51_, r_n_263__50_, r_n_263__49_, r_n_263__48_, r_n_263__47_, r_n_263__46_, r_n_263__45_, r_n_263__44_, r_n_263__43_, r_n_263__42_, r_n_263__41_, r_n_263__40_, r_n_263__39_, r_n_263__38_, r_n_263__37_, r_n_263__36_, r_n_263__35_, r_n_263__34_, r_n_263__33_, r_n_263__32_, r_n_263__31_, r_n_263__30_, r_n_263__29_, r_n_263__28_, r_n_263__27_, r_n_263__26_, r_n_263__25_, r_n_263__24_, r_n_263__23_, r_n_263__22_, r_n_263__21_, r_n_263__20_, r_n_263__19_, r_n_263__18_, r_n_263__17_, r_n_263__16_, r_n_263__15_, r_n_263__14_, r_n_263__13_, r_n_263__12_, r_n_263__11_, r_n_263__10_, r_n_263__9_, r_n_263__8_, r_n_263__7_, r_n_263__6_, r_n_263__5_, r_n_263__4_, r_n_263__3_, r_n_263__2_, r_n_263__1_, r_n_263__0_ } = (N526)? { r_264__63_, r_264__62_, r_264__61_, r_264__60_, r_264__59_, r_264__58_, r_264__57_, r_264__56_, r_264__55_, r_264__54_, r_264__53_, r_264__52_, r_264__51_, r_264__50_, r_264__49_, r_264__48_, r_264__47_, r_264__46_, r_264__45_, r_264__44_, r_264__43_, r_264__42_, r_264__41_, r_264__40_, r_264__39_, r_264__38_, r_264__37_, r_264__36_, r_264__35_, r_264__34_, r_264__33_, r_264__32_, r_264__31_, r_264__30_, r_264__29_, r_264__28_, r_264__27_, r_264__26_, r_264__25_, r_264__24_, r_264__23_, r_264__22_, r_264__21_, r_264__20_, r_264__19_, r_264__18_, r_264__17_, r_264__16_, r_264__15_, r_264__14_, r_264__13_, r_264__12_, r_264__11_, r_264__10_, r_264__9_, r_264__8_, r_264__7_, r_264__6_, r_264__5_, r_264__4_, r_264__3_, r_264__2_, r_264__1_, r_264__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N527)? data_i : 1'b0;
  assign N526 = sel_i[526];
  assign N527 = N2343;
  assign { r_n_264__63_, r_n_264__62_, r_n_264__61_, r_n_264__60_, r_n_264__59_, r_n_264__58_, r_n_264__57_, r_n_264__56_, r_n_264__55_, r_n_264__54_, r_n_264__53_, r_n_264__52_, r_n_264__51_, r_n_264__50_, r_n_264__49_, r_n_264__48_, r_n_264__47_, r_n_264__46_, r_n_264__45_, r_n_264__44_, r_n_264__43_, r_n_264__42_, r_n_264__41_, r_n_264__40_, r_n_264__39_, r_n_264__38_, r_n_264__37_, r_n_264__36_, r_n_264__35_, r_n_264__34_, r_n_264__33_, r_n_264__32_, r_n_264__31_, r_n_264__30_, r_n_264__29_, r_n_264__28_, r_n_264__27_, r_n_264__26_, r_n_264__25_, r_n_264__24_, r_n_264__23_, r_n_264__22_, r_n_264__21_, r_n_264__20_, r_n_264__19_, r_n_264__18_, r_n_264__17_, r_n_264__16_, r_n_264__15_, r_n_264__14_, r_n_264__13_, r_n_264__12_, r_n_264__11_, r_n_264__10_, r_n_264__9_, r_n_264__8_, r_n_264__7_, r_n_264__6_, r_n_264__5_, r_n_264__4_, r_n_264__3_, r_n_264__2_, r_n_264__1_, r_n_264__0_ } = (N528)? { r_265__63_, r_265__62_, r_265__61_, r_265__60_, r_265__59_, r_265__58_, r_265__57_, r_265__56_, r_265__55_, r_265__54_, r_265__53_, r_265__52_, r_265__51_, r_265__50_, r_265__49_, r_265__48_, r_265__47_, r_265__46_, r_265__45_, r_265__44_, r_265__43_, r_265__42_, r_265__41_, r_265__40_, r_265__39_, r_265__38_, r_265__37_, r_265__36_, r_265__35_, r_265__34_, r_265__33_, r_265__32_, r_265__31_, r_265__30_, r_265__29_, r_265__28_, r_265__27_, r_265__26_, r_265__25_, r_265__24_, r_265__23_, r_265__22_, r_265__21_, r_265__20_, r_265__19_, r_265__18_, r_265__17_, r_265__16_, r_265__15_, r_265__14_, r_265__13_, r_265__12_, r_265__11_, r_265__10_, r_265__9_, r_265__8_, r_265__7_, r_265__6_, r_265__5_, r_265__4_, r_265__3_, r_265__2_, r_265__1_, r_265__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N529)? data_i : 1'b0;
  assign N528 = sel_i[528];
  assign N529 = N2348;
  assign { r_n_265__63_, r_n_265__62_, r_n_265__61_, r_n_265__60_, r_n_265__59_, r_n_265__58_, r_n_265__57_, r_n_265__56_, r_n_265__55_, r_n_265__54_, r_n_265__53_, r_n_265__52_, r_n_265__51_, r_n_265__50_, r_n_265__49_, r_n_265__48_, r_n_265__47_, r_n_265__46_, r_n_265__45_, r_n_265__44_, r_n_265__43_, r_n_265__42_, r_n_265__41_, r_n_265__40_, r_n_265__39_, r_n_265__38_, r_n_265__37_, r_n_265__36_, r_n_265__35_, r_n_265__34_, r_n_265__33_, r_n_265__32_, r_n_265__31_, r_n_265__30_, r_n_265__29_, r_n_265__28_, r_n_265__27_, r_n_265__26_, r_n_265__25_, r_n_265__24_, r_n_265__23_, r_n_265__22_, r_n_265__21_, r_n_265__20_, r_n_265__19_, r_n_265__18_, r_n_265__17_, r_n_265__16_, r_n_265__15_, r_n_265__14_, r_n_265__13_, r_n_265__12_, r_n_265__11_, r_n_265__10_, r_n_265__9_, r_n_265__8_, r_n_265__7_, r_n_265__6_, r_n_265__5_, r_n_265__4_, r_n_265__3_, r_n_265__2_, r_n_265__1_, r_n_265__0_ } = (N530)? { r_266__63_, r_266__62_, r_266__61_, r_266__60_, r_266__59_, r_266__58_, r_266__57_, r_266__56_, r_266__55_, r_266__54_, r_266__53_, r_266__52_, r_266__51_, r_266__50_, r_266__49_, r_266__48_, r_266__47_, r_266__46_, r_266__45_, r_266__44_, r_266__43_, r_266__42_, r_266__41_, r_266__40_, r_266__39_, r_266__38_, r_266__37_, r_266__36_, r_266__35_, r_266__34_, r_266__33_, r_266__32_, r_266__31_, r_266__30_, r_266__29_, r_266__28_, r_266__27_, r_266__26_, r_266__25_, r_266__24_, r_266__23_, r_266__22_, r_266__21_, r_266__20_, r_266__19_, r_266__18_, r_266__17_, r_266__16_, r_266__15_, r_266__14_, r_266__13_, r_266__12_, r_266__11_, r_266__10_, r_266__9_, r_266__8_, r_266__7_, r_266__6_, r_266__5_, r_266__4_, r_266__3_, r_266__2_, r_266__1_, r_266__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N531)? data_i : 1'b0;
  assign N530 = sel_i[530];
  assign N531 = N2353;
  assign { r_n_266__63_, r_n_266__62_, r_n_266__61_, r_n_266__60_, r_n_266__59_, r_n_266__58_, r_n_266__57_, r_n_266__56_, r_n_266__55_, r_n_266__54_, r_n_266__53_, r_n_266__52_, r_n_266__51_, r_n_266__50_, r_n_266__49_, r_n_266__48_, r_n_266__47_, r_n_266__46_, r_n_266__45_, r_n_266__44_, r_n_266__43_, r_n_266__42_, r_n_266__41_, r_n_266__40_, r_n_266__39_, r_n_266__38_, r_n_266__37_, r_n_266__36_, r_n_266__35_, r_n_266__34_, r_n_266__33_, r_n_266__32_, r_n_266__31_, r_n_266__30_, r_n_266__29_, r_n_266__28_, r_n_266__27_, r_n_266__26_, r_n_266__25_, r_n_266__24_, r_n_266__23_, r_n_266__22_, r_n_266__21_, r_n_266__20_, r_n_266__19_, r_n_266__18_, r_n_266__17_, r_n_266__16_, r_n_266__15_, r_n_266__14_, r_n_266__13_, r_n_266__12_, r_n_266__11_, r_n_266__10_, r_n_266__9_, r_n_266__8_, r_n_266__7_, r_n_266__6_, r_n_266__5_, r_n_266__4_, r_n_266__3_, r_n_266__2_, r_n_266__1_, r_n_266__0_ } = (N532)? { r_267__63_, r_267__62_, r_267__61_, r_267__60_, r_267__59_, r_267__58_, r_267__57_, r_267__56_, r_267__55_, r_267__54_, r_267__53_, r_267__52_, r_267__51_, r_267__50_, r_267__49_, r_267__48_, r_267__47_, r_267__46_, r_267__45_, r_267__44_, r_267__43_, r_267__42_, r_267__41_, r_267__40_, r_267__39_, r_267__38_, r_267__37_, r_267__36_, r_267__35_, r_267__34_, r_267__33_, r_267__32_, r_267__31_, r_267__30_, r_267__29_, r_267__28_, r_267__27_, r_267__26_, r_267__25_, r_267__24_, r_267__23_, r_267__22_, r_267__21_, r_267__20_, r_267__19_, r_267__18_, r_267__17_, r_267__16_, r_267__15_, r_267__14_, r_267__13_, r_267__12_, r_267__11_, r_267__10_, r_267__9_, r_267__8_, r_267__7_, r_267__6_, r_267__5_, r_267__4_, r_267__3_, r_267__2_, r_267__1_, r_267__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N533)? data_i : 1'b0;
  assign N532 = sel_i[532];
  assign N533 = N2358;
  assign { r_n_267__63_, r_n_267__62_, r_n_267__61_, r_n_267__60_, r_n_267__59_, r_n_267__58_, r_n_267__57_, r_n_267__56_, r_n_267__55_, r_n_267__54_, r_n_267__53_, r_n_267__52_, r_n_267__51_, r_n_267__50_, r_n_267__49_, r_n_267__48_, r_n_267__47_, r_n_267__46_, r_n_267__45_, r_n_267__44_, r_n_267__43_, r_n_267__42_, r_n_267__41_, r_n_267__40_, r_n_267__39_, r_n_267__38_, r_n_267__37_, r_n_267__36_, r_n_267__35_, r_n_267__34_, r_n_267__33_, r_n_267__32_, r_n_267__31_, r_n_267__30_, r_n_267__29_, r_n_267__28_, r_n_267__27_, r_n_267__26_, r_n_267__25_, r_n_267__24_, r_n_267__23_, r_n_267__22_, r_n_267__21_, r_n_267__20_, r_n_267__19_, r_n_267__18_, r_n_267__17_, r_n_267__16_, r_n_267__15_, r_n_267__14_, r_n_267__13_, r_n_267__12_, r_n_267__11_, r_n_267__10_, r_n_267__9_, r_n_267__8_, r_n_267__7_, r_n_267__6_, r_n_267__5_, r_n_267__4_, r_n_267__3_, r_n_267__2_, r_n_267__1_, r_n_267__0_ } = (N534)? { r_268__63_, r_268__62_, r_268__61_, r_268__60_, r_268__59_, r_268__58_, r_268__57_, r_268__56_, r_268__55_, r_268__54_, r_268__53_, r_268__52_, r_268__51_, r_268__50_, r_268__49_, r_268__48_, r_268__47_, r_268__46_, r_268__45_, r_268__44_, r_268__43_, r_268__42_, r_268__41_, r_268__40_, r_268__39_, r_268__38_, r_268__37_, r_268__36_, r_268__35_, r_268__34_, r_268__33_, r_268__32_, r_268__31_, r_268__30_, r_268__29_, r_268__28_, r_268__27_, r_268__26_, r_268__25_, r_268__24_, r_268__23_, r_268__22_, r_268__21_, r_268__20_, r_268__19_, r_268__18_, r_268__17_, r_268__16_, r_268__15_, r_268__14_, r_268__13_, r_268__12_, r_268__11_, r_268__10_, r_268__9_, r_268__8_, r_268__7_, r_268__6_, r_268__5_, r_268__4_, r_268__3_, r_268__2_, r_268__1_, r_268__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N535)? data_i : 1'b0;
  assign N534 = sel_i[534];
  assign N535 = N2363;
  assign { r_n_268__63_, r_n_268__62_, r_n_268__61_, r_n_268__60_, r_n_268__59_, r_n_268__58_, r_n_268__57_, r_n_268__56_, r_n_268__55_, r_n_268__54_, r_n_268__53_, r_n_268__52_, r_n_268__51_, r_n_268__50_, r_n_268__49_, r_n_268__48_, r_n_268__47_, r_n_268__46_, r_n_268__45_, r_n_268__44_, r_n_268__43_, r_n_268__42_, r_n_268__41_, r_n_268__40_, r_n_268__39_, r_n_268__38_, r_n_268__37_, r_n_268__36_, r_n_268__35_, r_n_268__34_, r_n_268__33_, r_n_268__32_, r_n_268__31_, r_n_268__30_, r_n_268__29_, r_n_268__28_, r_n_268__27_, r_n_268__26_, r_n_268__25_, r_n_268__24_, r_n_268__23_, r_n_268__22_, r_n_268__21_, r_n_268__20_, r_n_268__19_, r_n_268__18_, r_n_268__17_, r_n_268__16_, r_n_268__15_, r_n_268__14_, r_n_268__13_, r_n_268__12_, r_n_268__11_, r_n_268__10_, r_n_268__9_, r_n_268__8_, r_n_268__7_, r_n_268__6_, r_n_268__5_, r_n_268__4_, r_n_268__3_, r_n_268__2_, r_n_268__1_, r_n_268__0_ } = (N536)? { r_269__63_, r_269__62_, r_269__61_, r_269__60_, r_269__59_, r_269__58_, r_269__57_, r_269__56_, r_269__55_, r_269__54_, r_269__53_, r_269__52_, r_269__51_, r_269__50_, r_269__49_, r_269__48_, r_269__47_, r_269__46_, r_269__45_, r_269__44_, r_269__43_, r_269__42_, r_269__41_, r_269__40_, r_269__39_, r_269__38_, r_269__37_, r_269__36_, r_269__35_, r_269__34_, r_269__33_, r_269__32_, r_269__31_, r_269__30_, r_269__29_, r_269__28_, r_269__27_, r_269__26_, r_269__25_, r_269__24_, r_269__23_, r_269__22_, r_269__21_, r_269__20_, r_269__19_, r_269__18_, r_269__17_, r_269__16_, r_269__15_, r_269__14_, r_269__13_, r_269__12_, r_269__11_, r_269__10_, r_269__9_, r_269__8_, r_269__7_, r_269__6_, r_269__5_, r_269__4_, r_269__3_, r_269__2_, r_269__1_, r_269__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N537)? data_i : 1'b0;
  assign N536 = sel_i[536];
  assign N537 = N2368;
  assign { r_n_269__63_, r_n_269__62_, r_n_269__61_, r_n_269__60_, r_n_269__59_, r_n_269__58_, r_n_269__57_, r_n_269__56_, r_n_269__55_, r_n_269__54_, r_n_269__53_, r_n_269__52_, r_n_269__51_, r_n_269__50_, r_n_269__49_, r_n_269__48_, r_n_269__47_, r_n_269__46_, r_n_269__45_, r_n_269__44_, r_n_269__43_, r_n_269__42_, r_n_269__41_, r_n_269__40_, r_n_269__39_, r_n_269__38_, r_n_269__37_, r_n_269__36_, r_n_269__35_, r_n_269__34_, r_n_269__33_, r_n_269__32_, r_n_269__31_, r_n_269__30_, r_n_269__29_, r_n_269__28_, r_n_269__27_, r_n_269__26_, r_n_269__25_, r_n_269__24_, r_n_269__23_, r_n_269__22_, r_n_269__21_, r_n_269__20_, r_n_269__19_, r_n_269__18_, r_n_269__17_, r_n_269__16_, r_n_269__15_, r_n_269__14_, r_n_269__13_, r_n_269__12_, r_n_269__11_, r_n_269__10_, r_n_269__9_, r_n_269__8_, r_n_269__7_, r_n_269__6_, r_n_269__5_, r_n_269__4_, r_n_269__3_, r_n_269__2_, r_n_269__1_, r_n_269__0_ } = (N538)? { r_270__63_, r_270__62_, r_270__61_, r_270__60_, r_270__59_, r_270__58_, r_270__57_, r_270__56_, r_270__55_, r_270__54_, r_270__53_, r_270__52_, r_270__51_, r_270__50_, r_270__49_, r_270__48_, r_270__47_, r_270__46_, r_270__45_, r_270__44_, r_270__43_, r_270__42_, r_270__41_, r_270__40_, r_270__39_, r_270__38_, r_270__37_, r_270__36_, r_270__35_, r_270__34_, r_270__33_, r_270__32_, r_270__31_, r_270__30_, r_270__29_, r_270__28_, r_270__27_, r_270__26_, r_270__25_, r_270__24_, r_270__23_, r_270__22_, r_270__21_, r_270__20_, r_270__19_, r_270__18_, r_270__17_, r_270__16_, r_270__15_, r_270__14_, r_270__13_, r_270__12_, r_270__11_, r_270__10_, r_270__9_, r_270__8_, r_270__7_, r_270__6_, r_270__5_, r_270__4_, r_270__3_, r_270__2_, r_270__1_, r_270__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N539)? data_i : 1'b0;
  assign N538 = sel_i[538];
  assign N539 = N2373;
  assign { r_n_270__63_, r_n_270__62_, r_n_270__61_, r_n_270__60_, r_n_270__59_, r_n_270__58_, r_n_270__57_, r_n_270__56_, r_n_270__55_, r_n_270__54_, r_n_270__53_, r_n_270__52_, r_n_270__51_, r_n_270__50_, r_n_270__49_, r_n_270__48_, r_n_270__47_, r_n_270__46_, r_n_270__45_, r_n_270__44_, r_n_270__43_, r_n_270__42_, r_n_270__41_, r_n_270__40_, r_n_270__39_, r_n_270__38_, r_n_270__37_, r_n_270__36_, r_n_270__35_, r_n_270__34_, r_n_270__33_, r_n_270__32_, r_n_270__31_, r_n_270__30_, r_n_270__29_, r_n_270__28_, r_n_270__27_, r_n_270__26_, r_n_270__25_, r_n_270__24_, r_n_270__23_, r_n_270__22_, r_n_270__21_, r_n_270__20_, r_n_270__19_, r_n_270__18_, r_n_270__17_, r_n_270__16_, r_n_270__15_, r_n_270__14_, r_n_270__13_, r_n_270__12_, r_n_270__11_, r_n_270__10_, r_n_270__9_, r_n_270__8_, r_n_270__7_, r_n_270__6_, r_n_270__5_, r_n_270__4_, r_n_270__3_, r_n_270__2_, r_n_270__1_, r_n_270__0_ } = (N540)? { r_271__63_, r_271__62_, r_271__61_, r_271__60_, r_271__59_, r_271__58_, r_271__57_, r_271__56_, r_271__55_, r_271__54_, r_271__53_, r_271__52_, r_271__51_, r_271__50_, r_271__49_, r_271__48_, r_271__47_, r_271__46_, r_271__45_, r_271__44_, r_271__43_, r_271__42_, r_271__41_, r_271__40_, r_271__39_, r_271__38_, r_271__37_, r_271__36_, r_271__35_, r_271__34_, r_271__33_, r_271__32_, r_271__31_, r_271__30_, r_271__29_, r_271__28_, r_271__27_, r_271__26_, r_271__25_, r_271__24_, r_271__23_, r_271__22_, r_271__21_, r_271__20_, r_271__19_, r_271__18_, r_271__17_, r_271__16_, r_271__15_, r_271__14_, r_271__13_, r_271__12_, r_271__11_, r_271__10_, r_271__9_, r_271__8_, r_271__7_, r_271__6_, r_271__5_, r_271__4_, r_271__3_, r_271__2_, r_271__1_, r_271__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N541)? data_i : 1'b0;
  assign N540 = sel_i[540];
  assign N541 = N2378;
  assign { r_n_271__63_, r_n_271__62_, r_n_271__61_, r_n_271__60_, r_n_271__59_, r_n_271__58_, r_n_271__57_, r_n_271__56_, r_n_271__55_, r_n_271__54_, r_n_271__53_, r_n_271__52_, r_n_271__51_, r_n_271__50_, r_n_271__49_, r_n_271__48_, r_n_271__47_, r_n_271__46_, r_n_271__45_, r_n_271__44_, r_n_271__43_, r_n_271__42_, r_n_271__41_, r_n_271__40_, r_n_271__39_, r_n_271__38_, r_n_271__37_, r_n_271__36_, r_n_271__35_, r_n_271__34_, r_n_271__33_, r_n_271__32_, r_n_271__31_, r_n_271__30_, r_n_271__29_, r_n_271__28_, r_n_271__27_, r_n_271__26_, r_n_271__25_, r_n_271__24_, r_n_271__23_, r_n_271__22_, r_n_271__21_, r_n_271__20_, r_n_271__19_, r_n_271__18_, r_n_271__17_, r_n_271__16_, r_n_271__15_, r_n_271__14_, r_n_271__13_, r_n_271__12_, r_n_271__11_, r_n_271__10_, r_n_271__9_, r_n_271__8_, r_n_271__7_, r_n_271__6_, r_n_271__5_, r_n_271__4_, r_n_271__3_, r_n_271__2_, r_n_271__1_, r_n_271__0_ } = (N542)? { r_272__63_, r_272__62_, r_272__61_, r_272__60_, r_272__59_, r_272__58_, r_272__57_, r_272__56_, r_272__55_, r_272__54_, r_272__53_, r_272__52_, r_272__51_, r_272__50_, r_272__49_, r_272__48_, r_272__47_, r_272__46_, r_272__45_, r_272__44_, r_272__43_, r_272__42_, r_272__41_, r_272__40_, r_272__39_, r_272__38_, r_272__37_, r_272__36_, r_272__35_, r_272__34_, r_272__33_, r_272__32_, r_272__31_, r_272__30_, r_272__29_, r_272__28_, r_272__27_, r_272__26_, r_272__25_, r_272__24_, r_272__23_, r_272__22_, r_272__21_, r_272__20_, r_272__19_, r_272__18_, r_272__17_, r_272__16_, r_272__15_, r_272__14_, r_272__13_, r_272__12_, r_272__11_, r_272__10_, r_272__9_, r_272__8_, r_272__7_, r_272__6_, r_272__5_, r_272__4_, r_272__3_, r_272__2_, r_272__1_, r_272__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N543)? data_i : 1'b0;
  assign N542 = sel_i[542];
  assign N543 = N2383;
  assign { r_n_272__63_, r_n_272__62_, r_n_272__61_, r_n_272__60_, r_n_272__59_, r_n_272__58_, r_n_272__57_, r_n_272__56_, r_n_272__55_, r_n_272__54_, r_n_272__53_, r_n_272__52_, r_n_272__51_, r_n_272__50_, r_n_272__49_, r_n_272__48_, r_n_272__47_, r_n_272__46_, r_n_272__45_, r_n_272__44_, r_n_272__43_, r_n_272__42_, r_n_272__41_, r_n_272__40_, r_n_272__39_, r_n_272__38_, r_n_272__37_, r_n_272__36_, r_n_272__35_, r_n_272__34_, r_n_272__33_, r_n_272__32_, r_n_272__31_, r_n_272__30_, r_n_272__29_, r_n_272__28_, r_n_272__27_, r_n_272__26_, r_n_272__25_, r_n_272__24_, r_n_272__23_, r_n_272__22_, r_n_272__21_, r_n_272__20_, r_n_272__19_, r_n_272__18_, r_n_272__17_, r_n_272__16_, r_n_272__15_, r_n_272__14_, r_n_272__13_, r_n_272__12_, r_n_272__11_, r_n_272__10_, r_n_272__9_, r_n_272__8_, r_n_272__7_, r_n_272__6_, r_n_272__5_, r_n_272__4_, r_n_272__3_, r_n_272__2_, r_n_272__1_, r_n_272__0_ } = (N544)? { r_273__63_, r_273__62_, r_273__61_, r_273__60_, r_273__59_, r_273__58_, r_273__57_, r_273__56_, r_273__55_, r_273__54_, r_273__53_, r_273__52_, r_273__51_, r_273__50_, r_273__49_, r_273__48_, r_273__47_, r_273__46_, r_273__45_, r_273__44_, r_273__43_, r_273__42_, r_273__41_, r_273__40_, r_273__39_, r_273__38_, r_273__37_, r_273__36_, r_273__35_, r_273__34_, r_273__33_, r_273__32_, r_273__31_, r_273__30_, r_273__29_, r_273__28_, r_273__27_, r_273__26_, r_273__25_, r_273__24_, r_273__23_, r_273__22_, r_273__21_, r_273__20_, r_273__19_, r_273__18_, r_273__17_, r_273__16_, r_273__15_, r_273__14_, r_273__13_, r_273__12_, r_273__11_, r_273__10_, r_273__9_, r_273__8_, r_273__7_, r_273__6_, r_273__5_, r_273__4_, r_273__3_, r_273__2_, r_273__1_, r_273__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N545)? data_i : 1'b0;
  assign N544 = sel_i[544];
  assign N545 = N2388;
  assign { r_n_273__63_, r_n_273__62_, r_n_273__61_, r_n_273__60_, r_n_273__59_, r_n_273__58_, r_n_273__57_, r_n_273__56_, r_n_273__55_, r_n_273__54_, r_n_273__53_, r_n_273__52_, r_n_273__51_, r_n_273__50_, r_n_273__49_, r_n_273__48_, r_n_273__47_, r_n_273__46_, r_n_273__45_, r_n_273__44_, r_n_273__43_, r_n_273__42_, r_n_273__41_, r_n_273__40_, r_n_273__39_, r_n_273__38_, r_n_273__37_, r_n_273__36_, r_n_273__35_, r_n_273__34_, r_n_273__33_, r_n_273__32_, r_n_273__31_, r_n_273__30_, r_n_273__29_, r_n_273__28_, r_n_273__27_, r_n_273__26_, r_n_273__25_, r_n_273__24_, r_n_273__23_, r_n_273__22_, r_n_273__21_, r_n_273__20_, r_n_273__19_, r_n_273__18_, r_n_273__17_, r_n_273__16_, r_n_273__15_, r_n_273__14_, r_n_273__13_, r_n_273__12_, r_n_273__11_, r_n_273__10_, r_n_273__9_, r_n_273__8_, r_n_273__7_, r_n_273__6_, r_n_273__5_, r_n_273__4_, r_n_273__3_, r_n_273__2_, r_n_273__1_, r_n_273__0_ } = (N546)? { r_274__63_, r_274__62_, r_274__61_, r_274__60_, r_274__59_, r_274__58_, r_274__57_, r_274__56_, r_274__55_, r_274__54_, r_274__53_, r_274__52_, r_274__51_, r_274__50_, r_274__49_, r_274__48_, r_274__47_, r_274__46_, r_274__45_, r_274__44_, r_274__43_, r_274__42_, r_274__41_, r_274__40_, r_274__39_, r_274__38_, r_274__37_, r_274__36_, r_274__35_, r_274__34_, r_274__33_, r_274__32_, r_274__31_, r_274__30_, r_274__29_, r_274__28_, r_274__27_, r_274__26_, r_274__25_, r_274__24_, r_274__23_, r_274__22_, r_274__21_, r_274__20_, r_274__19_, r_274__18_, r_274__17_, r_274__16_, r_274__15_, r_274__14_, r_274__13_, r_274__12_, r_274__11_, r_274__10_, r_274__9_, r_274__8_, r_274__7_, r_274__6_, r_274__5_, r_274__4_, r_274__3_, r_274__2_, r_274__1_, r_274__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N547)? data_i : 1'b0;
  assign N546 = sel_i[546];
  assign N547 = N2393;
  assign { r_n_274__63_, r_n_274__62_, r_n_274__61_, r_n_274__60_, r_n_274__59_, r_n_274__58_, r_n_274__57_, r_n_274__56_, r_n_274__55_, r_n_274__54_, r_n_274__53_, r_n_274__52_, r_n_274__51_, r_n_274__50_, r_n_274__49_, r_n_274__48_, r_n_274__47_, r_n_274__46_, r_n_274__45_, r_n_274__44_, r_n_274__43_, r_n_274__42_, r_n_274__41_, r_n_274__40_, r_n_274__39_, r_n_274__38_, r_n_274__37_, r_n_274__36_, r_n_274__35_, r_n_274__34_, r_n_274__33_, r_n_274__32_, r_n_274__31_, r_n_274__30_, r_n_274__29_, r_n_274__28_, r_n_274__27_, r_n_274__26_, r_n_274__25_, r_n_274__24_, r_n_274__23_, r_n_274__22_, r_n_274__21_, r_n_274__20_, r_n_274__19_, r_n_274__18_, r_n_274__17_, r_n_274__16_, r_n_274__15_, r_n_274__14_, r_n_274__13_, r_n_274__12_, r_n_274__11_, r_n_274__10_, r_n_274__9_, r_n_274__8_, r_n_274__7_, r_n_274__6_, r_n_274__5_, r_n_274__4_, r_n_274__3_, r_n_274__2_, r_n_274__1_, r_n_274__0_ } = (N548)? { r_275__63_, r_275__62_, r_275__61_, r_275__60_, r_275__59_, r_275__58_, r_275__57_, r_275__56_, r_275__55_, r_275__54_, r_275__53_, r_275__52_, r_275__51_, r_275__50_, r_275__49_, r_275__48_, r_275__47_, r_275__46_, r_275__45_, r_275__44_, r_275__43_, r_275__42_, r_275__41_, r_275__40_, r_275__39_, r_275__38_, r_275__37_, r_275__36_, r_275__35_, r_275__34_, r_275__33_, r_275__32_, r_275__31_, r_275__30_, r_275__29_, r_275__28_, r_275__27_, r_275__26_, r_275__25_, r_275__24_, r_275__23_, r_275__22_, r_275__21_, r_275__20_, r_275__19_, r_275__18_, r_275__17_, r_275__16_, r_275__15_, r_275__14_, r_275__13_, r_275__12_, r_275__11_, r_275__10_, r_275__9_, r_275__8_, r_275__7_, r_275__6_, r_275__5_, r_275__4_, r_275__3_, r_275__2_, r_275__1_, r_275__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N549)? data_i : 1'b0;
  assign N548 = sel_i[548];
  assign N549 = N2398;
  assign { r_n_275__63_, r_n_275__62_, r_n_275__61_, r_n_275__60_, r_n_275__59_, r_n_275__58_, r_n_275__57_, r_n_275__56_, r_n_275__55_, r_n_275__54_, r_n_275__53_, r_n_275__52_, r_n_275__51_, r_n_275__50_, r_n_275__49_, r_n_275__48_, r_n_275__47_, r_n_275__46_, r_n_275__45_, r_n_275__44_, r_n_275__43_, r_n_275__42_, r_n_275__41_, r_n_275__40_, r_n_275__39_, r_n_275__38_, r_n_275__37_, r_n_275__36_, r_n_275__35_, r_n_275__34_, r_n_275__33_, r_n_275__32_, r_n_275__31_, r_n_275__30_, r_n_275__29_, r_n_275__28_, r_n_275__27_, r_n_275__26_, r_n_275__25_, r_n_275__24_, r_n_275__23_, r_n_275__22_, r_n_275__21_, r_n_275__20_, r_n_275__19_, r_n_275__18_, r_n_275__17_, r_n_275__16_, r_n_275__15_, r_n_275__14_, r_n_275__13_, r_n_275__12_, r_n_275__11_, r_n_275__10_, r_n_275__9_, r_n_275__8_, r_n_275__7_, r_n_275__6_, r_n_275__5_, r_n_275__4_, r_n_275__3_, r_n_275__2_, r_n_275__1_, r_n_275__0_ } = (N550)? { r_276__63_, r_276__62_, r_276__61_, r_276__60_, r_276__59_, r_276__58_, r_276__57_, r_276__56_, r_276__55_, r_276__54_, r_276__53_, r_276__52_, r_276__51_, r_276__50_, r_276__49_, r_276__48_, r_276__47_, r_276__46_, r_276__45_, r_276__44_, r_276__43_, r_276__42_, r_276__41_, r_276__40_, r_276__39_, r_276__38_, r_276__37_, r_276__36_, r_276__35_, r_276__34_, r_276__33_, r_276__32_, r_276__31_, r_276__30_, r_276__29_, r_276__28_, r_276__27_, r_276__26_, r_276__25_, r_276__24_, r_276__23_, r_276__22_, r_276__21_, r_276__20_, r_276__19_, r_276__18_, r_276__17_, r_276__16_, r_276__15_, r_276__14_, r_276__13_, r_276__12_, r_276__11_, r_276__10_, r_276__9_, r_276__8_, r_276__7_, r_276__6_, r_276__5_, r_276__4_, r_276__3_, r_276__2_, r_276__1_, r_276__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N551)? data_i : 1'b0;
  assign N550 = sel_i[550];
  assign N551 = N2403;
  assign { r_n_276__63_, r_n_276__62_, r_n_276__61_, r_n_276__60_, r_n_276__59_, r_n_276__58_, r_n_276__57_, r_n_276__56_, r_n_276__55_, r_n_276__54_, r_n_276__53_, r_n_276__52_, r_n_276__51_, r_n_276__50_, r_n_276__49_, r_n_276__48_, r_n_276__47_, r_n_276__46_, r_n_276__45_, r_n_276__44_, r_n_276__43_, r_n_276__42_, r_n_276__41_, r_n_276__40_, r_n_276__39_, r_n_276__38_, r_n_276__37_, r_n_276__36_, r_n_276__35_, r_n_276__34_, r_n_276__33_, r_n_276__32_, r_n_276__31_, r_n_276__30_, r_n_276__29_, r_n_276__28_, r_n_276__27_, r_n_276__26_, r_n_276__25_, r_n_276__24_, r_n_276__23_, r_n_276__22_, r_n_276__21_, r_n_276__20_, r_n_276__19_, r_n_276__18_, r_n_276__17_, r_n_276__16_, r_n_276__15_, r_n_276__14_, r_n_276__13_, r_n_276__12_, r_n_276__11_, r_n_276__10_, r_n_276__9_, r_n_276__8_, r_n_276__7_, r_n_276__6_, r_n_276__5_, r_n_276__4_, r_n_276__3_, r_n_276__2_, r_n_276__1_, r_n_276__0_ } = (N552)? { r_277__63_, r_277__62_, r_277__61_, r_277__60_, r_277__59_, r_277__58_, r_277__57_, r_277__56_, r_277__55_, r_277__54_, r_277__53_, r_277__52_, r_277__51_, r_277__50_, r_277__49_, r_277__48_, r_277__47_, r_277__46_, r_277__45_, r_277__44_, r_277__43_, r_277__42_, r_277__41_, r_277__40_, r_277__39_, r_277__38_, r_277__37_, r_277__36_, r_277__35_, r_277__34_, r_277__33_, r_277__32_, r_277__31_, r_277__30_, r_277__29_, r_277__28_, r_277__27_, r_277__26_, r_277__25_, r_277__24_, r_277__23_, r_277__22_, r_277__21_, r_277__20_, r_277__19_, r_277__18_, r_277__17_, r_277__16_, r_277__15_, r_277__14_, r_277__13_, r_277__12_, r_277__11_, r_277__10_, r_277__9_, r_277__8_, r_277__7_, r_277__6_, r_277__5_, r_277__4_, r_277__3_, r_277__2_, r_277__1_, r_277__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N553)? data_i : 1'b0;
  assign N552 = sel_i[552];
  assign N553 = N2408;
  assign { r_n_277__63_, r_n_277__62_, r_n_277__61_, r_n_277__60_, r_n_277__59_, r_n_277__58_, r_n_277__57_, r_n_277__56_, r_n_277__55_, r_n_277__54_, r_n_277__53_, r_n_277__52_, r_n_277__51_, r_n_277__50_, r_n_277__49_, r_n_277__48_, r_n_277__47_, r_n_277__46_, r_n_277__45_, r_n_277__44_, r_n_277__43_, r_n_277__42_, r_n_277__41_, r_n_277__40_, r_n_277__39_, r_n_277__38_, r_n_277__37_, r_n_277__36_, r_n_277__35_, r_n_277__34_, r_n_277__33_, r_n_277__32_, r_n_277__31_, r_n_277__30_, r_n_277__29_, r_n_277__28_, r_n_277__27_, r_n_277__26_, r_n_277__25_, r_n_277__24_, r_n_277__23_, r_n_277__22_, r_n_277__21_, r_n_277__20_, r_n_277__19_, r_n_277__18_, r_n_277__17_, r_n_277__16_, r_n_277__15_, r_n_277__14_, r_n_277__13_, r_n_277__12_, r_n_277__11_, r_n_277__10_, r_n_277__9_, r_n_277__8_, r_n_277__7_, r_n_277__6_, r_n_277__5_, r_n_277__4_, r_n_277__3_, r_n_277__2_, r_n_277__1_, r_n_277__0_ } = (N554)? { r_278__63_, r_278__62_, r_278__61_, r_278__60_, r_278__59_, r_278__58_, r_278__57_, r_278__56_, r_278__55_, r_278__54_, r_278__53_, r_278__52_, r_278__51_, r_278__50_, r_278__49_, r_278__48_, r_278__47_, r_278__46_, r_278__45_, r_278__44_, r_278__43_, r_278__42_, r_278__41_, r_278__40_, r_278__39_, r_278__38_, r_278__37_, r_278__36_, r_278__35_, r_278__34_, r_278__33_, r_278__32_, r_278__31_, r_278__30_, r_278__29_, r_278__28_, r_278__27_, r_278__26_, r_278__25_, r_278__24_, r_278__23_, r_278__22_, r_278__21_, r_278__20_, r_278__19_, r_278__18_, r_278__17_, r_278__16_, r_278__15_, r_278__14_, r_278__13_, r_278__12_, r_278__11_, r_278__10_, r_278__9_, r_278__8_, r_278__7_, r_278__6_, r_278__5_, r_278__4_, r_278__3_, r_278__2_, r_278__1_, r_278__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N555)? data_i : 1'b0;
  assign N554 = sel_i[554];
  assign N555 = N2413;
  assign { r_n_278__63_, r_n_278__62_, r_n_278__61_, r_n_278__60_, r_n_278__59_, r_n_278__58_, r_n_278__57_, r_n_278__56_, r_n_278__55_, r_n_278__54_, r_n_278__53_, r_n_278__52_, r_n_278__51_, r_n_278__50_, r_n_278__49_, r_n_278__48_, r_n_278__47_, r_n_278__46_, r_n_278__45_, r_n_278__44_, r_n_278__43_, r_n_278__42_, r_n_278__41_, r_n_278__40_, r_n_278__39_, r_n_278__38_, r_n_278__37_, r_n_278__36_, r_n_278__35_, r_n_278__34_, r_n_278__33_, r_n_278__32_, r_n_278__31_, r_n_278__30_, r_n_278__29_, r_n_278__28_, r_n_278__27_, r_n_278__26_, r_n_278__25_, r_n_278__24_, r_n_278__23_, r_n_278__22_, r_n_278__21_, r_n_278__20_, r_n_278__19_, r_n_278__18_, r_n_278__17_, r_n_278__16_, r_n_278__15_, r_n_278__14_, r_n_278__13_, r_n_278__12_, r_n_278__11_, r_n_278__10_, r_n_278__9_, r_n_278__8_, r_n_278__7_, r_n_278__6_, r_n_278__5_, r_n_278__4_, r_n_278__3_, r_n_278__2_, r_n_278__1_, r_n_278__0_ } = (N556)? { r_279__63_, r_279__62_, r_279__61_, r_279__60_, r_279__59_, r_279__58_, r_279__57_, r_279__56_, r_279__55_, r_279__54_, r_279__53_, r_279__52_, r_279__51_, r_279__50_, r_279__49_, r_279__48_, r_279__47_, r_279__46_, r_279__45_, r_279__44_, r_279__43_, r_279__42_, r_279__41_, r_279__40_, r_279__39_, r_279__38_, r_279__37_, r_279__36_, r_279__35_, r_279__34_, r_279__33_, r_279__32_, r_279__31_, r_279__30_, r_279__29_, r_279__28_, r_279__27_, r_279__26_, r_279__25_, r_279__24_, r_279__23_, r_279__22_, r_279__21_, r_279__20_, r_279__19_, r_279__18_, r_279__17_, r_279__16_, r_279__15_, r_279__14_, r_279__13_, r_279__12_, r_279__11_, r_279__10_, r_279__9_, r_279__8_, r_279__7_, r_279__6_, r_279__5_, r_279__4_, r_279__3_, r_279__2_, r_279__1_, r_279__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N557)? data_i : 1'b0;
  assign N556 = sel_i[556];
  assign N557 = N2418;
  assign { r_n_279__63_, r_n_279__62_, r_n_279__61_, r_n_279__60_, r_n_279__59_, r_n_279__58_, r_n_279__57_, r_n_279__56_, r_n_279__55_, r_n_279__54_, r_n_279__53_, r_n_279__52_, r_n_279__51_, r_n_279__50_, r_n_279__49_, r_n_279__48_, r_n_279__47_, r_n_279__46_, r_n_279__45_, r_n_279__44_, r_n_279__43_, r_n_279__42_, r_n_279__41_, r_n_279__40_, r_n_279__39_, r_n_279__38_, r_n_279__37_, r_n_279__36_, r_n_279__35_, r_n_279__34_, r_n_279__33_, r_n_279__32_, r_n_279__31_, r_n_279__30_, r_n_279__29_, r_n_279__28_, r_n_279__27_, r_n_279__26_, r_n_279__25_, r_n_279__24_, r_n_279__23_, r_n_279__22_, r_n_279__21_, r_n_279__20_, r_n_279__19_, r_n_279__18_, r_n_279__17_, r_n_279__16_, r_n_279__15_, r_n_279__14_, r_n_279__13_, r_n_279__12_, r_n_279__11_, r_n_279__10_, r_n_279__9_, r_n_279__8_, r_n_279__7_, r_n_279__6_, r_n_279__5_, r_n_279__4_, r_n_279__3_, r_n_279__2_, r_n_279__1_, r_n_279__0_ } = (N558)? { r_280__63_, r_280__62_, r_280__61_, r_280__60_, r_280__59_, r_280__58_, r_280__57_, r_280__56_, r_280__55_, r_280__54_, r_280__53_, r_280__52_, r_280__51_, r_280__50_, r_280__49_, r_280__48_, r_280__47_, r_280__46_, r_280__45_, r_280__44_, r_280__43_, r_280__42_, r_280__41_, r_280__40_, r_280__39_, r_280__38_, r_280__37_, r_280__36_, r_280__35_, r_280__34_, r_280__33_, r_280__32_, r_280__31_, r_280__30_, r_280__29_, r_280__28_, r_280__27_, r_280__26_, r_280__25_, r_280__24_, r_280__23_, r_280__22_, r_280__21_, r_280__20_, r_280__19_, r_280__18_, r_280__17_, r_280__16_, r_280__15_, r_280__14_, r_280__13_, r_280__12_, r_280__11_, r_280__10_, r_280__9_, r_280__8_, r_280__7_, r_280__6_, r_280__5_, r_280__4_, r_280__3_, r_280__2_, r_280__1_, r_280__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N559)? data_i : 1'b0;
  assign N558 = sel_i[558];
  assign N559 = N2423;
  assign { r_n_280__63_, r_n_280__62_, r_n_280__61_, r_n_280__60_, r_n_280__59_, r_n_280__58_, r_n_280__57_, r_n_280__56_, r_n_280__55_, r_n_280__54_, r_n_280__53_, r_n_280__52_, r_n_280__51_, r_n_280__50_, r_n_280__49_, r_n_280__48_, r_n_280__47_, r_n_280__46_, r_n_280__45_, r_n_280__44_, r_n_280__43_, r_n_280__42_, r_n_280__41_, r_n_280__40_, r_n_280__39_, r_n_280__38_, r_n_280__37_, r_n_280__36_, r_n_280__35_, r_n_280__34_, r_n_280__33_, r_n_280__32_, r_n_280__31_, r_n_280__30_, r_n_280__29_, r_n_280__28_, r_n_280__27_, r_n_280__26_, r_n_280__25_, r_n_280__24_, r_n_280__23_, r_n_280__22_, r_n_280__21_, r_n_280__20_, r_n_280__19_, r_n_280__18_, r_n_280__17_, r_n_280__16_, r_n_280__15_, r_n_280__14_, r_n_280__13_, r_n_280__12_, r_n_280__11_, r_n_280__10_, r_n_280__9_, r_n_280__8_, r_n_280__7_, r_n_280__6_, r_n_280__5_, r_n_280__4_, r_n_280__3_, r_n_280__2_, r_n_280__1_, r_n_280__0_ } = (N560)? { r_281__63_, r_281__62_, r_281__61_, r_281__60_, r_281__59_, r_281__58_, r_281__57_, r_281__56_, r_281__55_, r_281__54_, r_281__53_, r_281__52_, r_281__51_, r_281__50_, r_281__49_, r_281__48_, r_281__47_, r_281__46_, r_281__45_, r_281__44_, r_281__43_, r_281__42_, r_281__41_, r_281__40_, r_281__39_, r_281__38_, r_281__37_, r_281__36_, r_281__35_, r_281__34_, r_281__33_, r_281__32_, r_281__31_, r_281__30_, r_281__29_, r_281__28_, r_281__27_, r_281__26_, r_281__25_, r_281__24_, r_281__23_, r_281__22_, r_281__21_, r_281__20_, r_281__19_, r_281__18_, r_281__17_, r_281__16_, r_281__15_, r_281__14_, r_281__13_, r_281__12_, r_281__11_, r_281__10_, r_281__9_, r_281__8_, r_281__7_, r_281__6_, r_281__5_, r_281__4_, r_281__3_, r_281__2_, r_281__1_, r_281__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N561)? data_i : 1'b0;
  assign N560 = sel_i[560];
  assign N561 = N2428;
  assign { r_n_281__63_, r_n_281__62_, r_n_281__61_, r_n_281__60_, r_n_281__59_, r_n_281__58_, r_n_281__57_, r_n_281__56_, r_n_281__55_, r_n_281__54_, r_n_281__53_, r_n_281__52_, r_n_281__51_, r_n_281__50_, r_n_281__49_, r_n_281__48_, r_n_281__47_, r_n_281__46_, r_n_281__45_, r_n_281__44_, r_n_281__43_, r_n_281__42_, r_n_281__41_, r_n_281__40_, r_n_281__39_, r_n_281__38_, r_n_281__37_, r_n_281__36_, r_n_281__35_, r_n_281__34_, r_n_281__33_, r_n_281__32_, r_n_281__31_, r_n_281__30_, r_n_281__29_, r_n_281__28_, r_n_281__27_, r_n_281__26_, r_n_281__25_, r_n_281__24_, r_n_281__23_, r_n_281__22_, r_n_281__21_, r_n_281__20_, r_n_281__19_, r_n_281__18_, r_n_281__17_, r_n_281__16_, r_n_281__15_, r_n_281__14_, r_n_281__13_, r_n_281__12_, r_n_281__11_, r_n_281__10_, r_n_281__9_, r_n_281__8_, r_n_281__7_, r_n_281__6_, r_n_281__5_, r_n_281__4_, r_n_281__3_, r_n_281__2_, r_n_281__1_, r_n_281__0_ } = (N562)? { r_282__63_, r_282__62_, r_282__61_, r_282__60_, r_282__59_, r_282__58_, r_282__57_, r_282__56_, r_282__55_, r_282__54_, r_282__53_, r_282__52_, r_282__51_, r_282__50_, r_282__49_, r_282__48_, r_282__47_, r_282__46_, r_282__45_, r_282__44_, r_282__43_, r_282__42_, r_282__41_, r_282__40_, r_282__39_, r_282__38_, r_282__37_, r_282__36_, r_282__35_, r_282__34_, r_282__33_, r_282__32_, r_282__31_, r_282__30_, r_282__29_, r_282__28_, r_282__27_, r_282__26_, r_282__25_, r_282__24_, r_282__23_, r_282__22_, r_282__21_, r_282__20_, r_282__19_, r_282__18_, r_282__17_, r_282__16_, r_282__15_, r_282__14_, r_282__13_, r_282__12_, r_282__11_, r_282__10_, r_282__9_, r_282__8_, r_282__7_, r_282__6_, r_282__5_, r_282__4_, r_282__3_, r_282__2_, r_282__1_, r_282__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N563)? data_i : 1'b0;
  assign N562 = sel_i[562];
  assign N563 = N2433;
  assign { r_n_282__63_, r_n_282__62_, r_n_282__61_, r_n_282__60_, r_n_282__59_, r_n_282__58_, r_n_282__57_, r_n_282__56_, r_n_282__55_, r_n_282__54_, r_n_282__53_, r_n_282__52_, r_n_282__51_, r_n_282__50_, r_n_282__49_, r_n_282__48_, r_n_282__47_, r_n_282__46_, r_n_282__45_, r_n_282__44_, r_n_282__43_, r_n_282__42_, r_n_282__41_, r_n_282__40_, r_n_282__39_, r_n_282__38_, r_n_282__37_, r_n_282__36_, r_n_282__35_, r_n_282__34_, r_n_282__33_, r_n_282__32_, r_n_282__31_, r_n_282__30_, r_n_282__29_, r_n_282__28_, r_n_282__27_, r_n_282__26_, r_n_282__25_, r_n_282__24_, r_n_282__23_, r_n_282__22_, r_n_282__21_, r_n_282__20_, r_n_282__19_, r_n_282__18_, r_n_282__17_, r_n_282__16_, r_n_282__15_, r_n_282__14_, r_n_282__13_, r_n_282__12_, r_n_282__11_, r_n_282__10_, r_n_282__9_, r_n_282__8_, r_n_282__7_, r_n_282__6_, r_n_282__5_, r_n_282__4_, r_n_282__3_, r_n_282__2_, r_n_282__1_, r_n_282__0_ } = (N564)? { r_283__63_, r_283__62_, r_283__61_, r_283__60_, r_283__59_, r_283__58_, r_283__57_, r_283__56_, r_283__55_, r_283__54_, r_283__53_, r_283__52_, r_283__51_, r_283__50_, r_283__49_, r_283__48_, r_283__47_, r_283__46_, r_283__45_, r_283__44_, r_283__43_, r_283__42_, r_283__41_, r_283__40_, r_283__39_, r_283__38_, r_283__37_, r_283__36_, r_283__35_, r_283__34_, r_283__33_, r_283__32_, r_283__31_, r_283__30_, r_283__29_, r_283__28_, r_283__27_, r_283__26_, r_283__25_, r_283__24_, r_283__23_, r_283__22_, r_283__21_, r_283__20_, r_283__19_, r_283__18_, r_283__17_, r_283__16_, r_283__15_, r_283__14_, r_283__13_, r_283__12_, r_283__11_, r_283__10_, r_283__9_, r_283__8_, r_283__7_, r_283__6_, r_283__5_, r_283__4_, r_283__3_, r_283__2_, r_283__1_, r_283__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N565)? data_i : 1'b0;
  assign N564 = sel_i[564];
  assign N565 = N2438;
  assign { r_n_283__63_, r_n_283__62_, r_n_283__61_, r_n_283__60_, r_n_283__59_, r_n_283__58_, r_n_283__57_, r_n_283__56_, r_n_283__55_, r_n_283__54_, r_n_283__53_, r_n_283__52_, r_n_283__51_, r_n_283__50_, r_n_283__49_, r_n_283__48_, r_n_283__47_, r_n_283__46_, r_n_283__45_, r_n_283__44_, r_n_283__43_, r_n_283__42_, r_n_283__41_, r_n_283__40_, r_n_283__39_, r_n_283__38_, r_n_283__37_, r_n_283__36_, r_n_283__35_, r_n_283__34_, r_n_283__33_, r_n_283__32_, r_n_283__31_, r_n_283__30_, r_n_283__29_, r_n_283__28_, r_n_283__27_, r_n_283__26_, r_n_283__25_, r_n_283__24_, r_n_283__23_, r_n_283__22_, r_n_283__21_, r_n_283__20_, r_n_283__19_, r_n_283__18_, r_n_283__17_, r_n_283__16_, r_n_283__15_, r_n_283__14_, r_n_283__13_, r_n_283__12_, r_n_283__11_, r_n_283__10_, r_n_283__9_, r_n_283__8_, r_n_283__7_, r_n_283__6_, r_n_283__5_, r_n_283__4_, r_n_283__3_, r_n_283__2_, r_n_283__1_, r_n_283__0_ } = (N566)? { r_284__63_, r_284__62_, r_284__61_, r_284__60_, r_284__59_, r_284__58_, r_284__57_, r_284__56_, r_284__55_, r_284__54_, r_284__53_, r_284__52_, r_284__51_, r_284__50_, r_284__49_, r_284__48_, r_284__47_, r_284__46_, r_284__45_, r_284__44_, r_284__43_, r_284__42_, r_284__41_, r_284__40_, r_284__39_, r_284__38_, r_284__37_, r_284__36_, r_284__35_, r_284__34_, r_284__33_, r_284__32_, r_284__31_, r_284__30_, r_284__29_, r_284__28_, r_284__27_, r_284__26_, r_284__25_, r_284__24_, r_284__23_, r_284__22_, r_284__21_, r_284__20_, r_284__19_, r_284__18_, r_284__17_, r_284__16_, r_284__15_, r_284__14_, r_284__13_, r_284__12_, r_284__11_, r_284__10_, r_284__9_, r_284__8_, r_284__7_, r_284__6_, r_284__5_, r_284__4_, r_284__3_, r_284__2_, r_284__1_, r_284__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N567)? data_i : 1'b0;
  assign N566 = sel_i[566];
  assign N567 = N2443;
  assign { r_n_284__63_, r_n_284__62_, r_n_284__61_, r_n_284__60_, r_n_284__59_, r_n_284__58_, r_n_284__57_, r_n_284__56_, r_n_284__55_, r_n_284__54_, r_n_284__53_, r_n_284__52_, r_n_284__51_, r_n_284__50_, r_n_284__49_, r_n_284__48_, r_n_284__47_, r_n_284__46_, r_n_284__45_, r_n_284__44_, r_n_284__43_, r_n_284__42_, r_n_284__41_, r_n_284__40_, r_n_284__39_, r_n_284__38_, r_n_284__37_, r_n_284__36_, r_n_284__35_, r_n_284__34_, r_n_284__33_, r_n_284__32_, r_n_284__31_, r_n_284__30_, r_n_284__29_, r_n_284__28_, r_n_284__27_, r_n_284__26_, r_n_284__25_, r_n_284__24_, r_n_284__23_, r_n_284__22_, r_n_284__21_, r_n_284__20_, r_n_284__19_, r_n_284__18_, r_n_284__17_, r_n_284__16_, r_n_284__15_, r_n_284__14_, r_n_284__13_, r_n_284__12_, r_n_284__11_, r_n_284__10_, r_n_284__9_, r_n_284__8_, r_n_284__7_, r_n_284__6_, r_n_284__5_, r_n_284__4_, r_n_284__3_, r_n_284__2_, r_n_284__1_, r_n_284__0_ } = (N568)? { r_285__63_, r_285__62_, r_285__61_, r_285__60_, r_285__59_, r_285__58_, r_285__57_, r_285__56_, r_285__55_, r_285__54_, r_285__53_, r_285__52_, r_285__51_, r_285__50_, r_285__49_, r_285__48_, r_285__47_, r_285__46_, r_285__45_, r_285__44_, r_285__43_, r_285__42_, r_285__41_, r_285__40_, r_285__39_, r_285__38_, r_285__37_, r_285__36_, r_285__35_, r_285__34_, r_285__33_, r_285__32_, r_285__31_, r_285__30_, r_285__29_, r_285__28_, r_285__27_, r_285__26_, r_285__25_, r_285__24_, r_285__23_, r_285__22_, r_285__21_, r_285__20_, r_285__19_, r_285__18_, r_285__17_, r_285__16_, r_285__15_, r_285__14_, r_285__13_, r_285__12_, r_285__11_, r_285__10_, r_285__9_, r_285__8_, r_285__7_, r_285__6_, r_285__5_, r_285__4_, r_285__3_, r_285__2_, r_285__1_, r_285__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N569)? data_i : 1'b0;
  assign N568 = sel_i[568];
  assign N569 = N2448;
  assign { r_n_285__63_, r_n_285__62_, r_n_285__61_, r_n_285__60_, r_n_285__59_, r_n_285__58_, r_n_285__57_, r_n_285__56_, r_n_285__55_, r_n_285__54_, r_n_285__53_, r_n_285__52_, r_n_285__51_, r_n_285__50_, r_n_285__49_, r_n_285__48_, r_n_285__47_, r_n_285__46_, r_n_285__45_, r_n_285__44_, r_n_285__43_, r_n_285__42_, r_n_285__41_, r_n_285__40_, r_n_285__39_, r_n_285__38_, r_n_285__37_, r_n_285__36_, r_n_285__35_, r_n_285__34_, r_n_285__33_, r_n_285__32_, r_n_285__31_, r_n_285__30_, r_n_285__29_, r_n_285__28_, r_n_285__27_, r_n_285__26_, r_n_285__25_, r_n_285__24_, r_n_285__23_, r_n_285__22_, r_n_285__21_, r_n_285__20_, r_n_285__19_, r_n_285__18_, r_n_285__17_, r_n_285__16_, r_n_285__15_, r_n_285__14_, r_n_285__13_, r_n_285__12_, r_n_285__11_, r_n_285__10_, r_n_285__9_, r_n_285__8_, r_n_285__7_, r_n_285__6_, r_n_285__5_, r_n_285__4_, r_n_285__3_, r_n_285__2_, r_n_285__1_, r_n_285__0_ } = (N570)? { r_286__63_, r_286__62_, r_286__61_, r_286__60_, r_286__59_, r_286__58_, r_286__57_, r_286__56_, r_286__55_, r_286__54_, r_286__53_, r_286__52_, r_286__51_, r_286__50_, r_286__49_, r_286__48_, r_286__47_, r_286__46_, r_286__45_, r_286__44_, r_286__43_, r_286__42_, r_286__41_, r_286__40_, r_286__39_, r_286__38_, r_286__37_, r_286__36_, r_286__35_, r_286__34_, r_286__33_, r_286__32_, r_286__31_, r_286__30_, r_286__29_, r_286__28_, r_286__27_, r_286__26_, r_286__25_, r_286__24_, r_286__23_, r_286__22_, r_286__21_, r_286__20_, r_286__19_, r_286__18_, r_286__17_, r_286__16_, r_286__15_, r_286__14_, r_286__13_, r_286__12_, r_286__11_, r_286__10_, r_286__9_, r_286__8_, r_286__7_, r_286__6_, r_286__5_, r_286__4_, r_286__3_, r_286__2_, r_286__1_, r_286__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N571)? data_i : 1'b0;
  assign N570 = sel_i[570];
  assign N571 = N2453;
  assign { r_n_286__63_, r_n_286__62_, r_n_286__61_, r_n_286__60_, r_n_286__59_, r_n_286__58_, r_n_286__57_, r_n_286__56_, r_n_286__55_, r_n_286__54_, r_n_286__53_, r_n_286__52_, r_n_286__51_, r_n_286__50_, r_n_286__49_, r_n_286__48_, r_n_286__47_, r_n_286__46_, r_n_286__45_, r_n_286__44_, r_n_286__43_, r_n_286__42_, r_n_286__41_, r_n_286__40_, r_n_286__39_, r_n_286__38_, r_n_286__37_, r_n_286__36_, r_n_286__35_, r_n_286__34_, r_n_286__33_, r_n_286__32_, r_n_286__31_, r_n_286__30_, r_n_286__29_, r_n_286__28_, r_n_286__27_, r_n_286__26_, r_n_286__25_, r_n_286__24_, r_n_286__23_, r_n_286__22_, r_n_286__21_, r_n_286__20_, r_n_286__19_, r_n_286__18_, r_n_286__17_, r_n_286__16_, r_n_286__15_, r_n_286__14_, r_n_286__13_, r_n_286__12_, r_n_286__11_, r_n_286__10_, r_n_286__9_, r_n_286__8_, r_n_286__7_, r_n_286__6_, r_n_286__5_, r_n_286__4_, r_n_286__3_, r_n_286__2_, r_n_286__1_, r_n_286__0_ } = (N572)? { r_287__63_, r_287__62_, r_287__61_, r_287__60_, r_287__59_, r_287__58_, r_287__57_, r_287__56_, r_287__55_, r_287__54_, r_287__53_, r_287__52_, r_287__51_, r_287__50_, r_287__49_, r_287__48_, r_287__47_, r_287__46_, r_287__45_, r_287__44_, r_287__43_, r_287__42_, r_287__41_, r_287__40_, r_287__39_, r_287__38_, r_287__37_, r_287__36_, r_287__35_, r_287__34_, r_287__33_, r_287__32_, r_287__31_, r_287__30_, r_287__29_, r_287__28_, r_287__27_, r_287__26_, r_287__25_, r_287__24_, r_287__23_, r_287__22_, r_287__21_, r_287__20_, r_287__19_, r_287__18_, r_287__17_, r_287__16_, r_287__15_, r_287__14_, r_287__13_, r_287__12_, r_287__11_, r_287__10_, r_287__9_, r_287__8_, r_287__7_, r_287__6_, r_287__5_, r_287__4_, r_287__3_, r_287__2_, r_287__1_, r_287__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N573)? data_i : 1'b0;
  assign N572 = sel_i[572];
  assign N573 = N2458;
  assign { r_n_287__63_, r_n_287__62_, r_n_287__61_, r_n_287__60_, r_n_287__59_, r_n_287__58_, r_n_287__57_, r_n_287__56_, r_n_287__55_, r_n_287__54_, r_n_287__53_, r_n_287__52_, r_n_287__51_, r_n_287__50_, r_n_287__49_, r_n_287__48_, r_n_287__47_, r_n_287__46_, r_n_287__45_, r_n_287__44_, r_n_287__43_, r_n_287__42_, r_n_287__41_, r_n_287__40_, r_n_287__39_, r_n_287__38_, r_n_287__37_, r_n_287__36_, r_n_287__35_, r_n_287__34_, r_n_287__33_, r_n_287__32_, r_n_287__31_, r_n_287__30_, r_n_287__29_, r_n_287__28_, r_n_287__27_, r_n_287__26_, r_n_287__25_, r_n_287__24_, r_n_287__23_, r_n_287__22_, r_n_287__21_, r_n_287__20_, r_n_287__19_, r_n_287__18_, r_n_287__17_, r_n_287__16_, r_n_287__15_, r_n_287__14_, r_n_287__13_, r_n_287__12_, r_n_287__11_, r_n_287__10_, r_n_287__9_, r_n_287__8_, r_n_287__7_, r_n_287__6_, r_n_287__5_, r_n_287__4_, r_n_287__3_, r_n_287__2_, r_n_287__1_, r_n_287__0_ } = (N574)? { r_288__63_, r_288__62_, r_288__61_, r_288__60_, r_288__59_, r_288__58_, r_288__57_, r_288__56_, r_288__55_, r_288__54_, r_288__53_, r_288__52_, r_288__51_, r_288__50_, r_288__49_, r_288__48_, r_288__47_, r_288__46_, r_288__45_, r_288__44_, r_288__43_, r_288__42_, r_288__41_, r_288__40_, r_288__39_, r_288__38_, r_288__37_, r_288__36_, r_288__35_, r_288__34_, r_288__33_, r_288__32_, r_288__31_, r_288__30_, r_288__29_, r_288__28_, r_288__27_, r_288__26_, r_288__25_, r_288__24_, r_288__23_, r_288__22_, r_288__21_, r_288__20_, r_288__19_, r_288__18_, r_288__17_, r_288__16_, r_288__15_, r_288__14_, r_288__13_, r_288__12_, r_288__11_, r_288__10_, r_288__9_, r_288__8_, r_288__7_, r_288__6_, r_288__5_, r_288__4_, r_288__3_, r_288__2_, r_288__1_, r_288__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N575)? data_i : 1'b0;
  assign N574 = sel_i[574];
  assign N575 = N2463;
  assign { r_n_288__63_, r_n_288__62_, r_n_288__61_, r_n_288__60_, r_n_288__59_, r_n_288__58_, r_n_288__57_, r_n_288__56_, r_n_288__55_, r_n_288__54_, r_n_288__53_, r_n_288__52_, r_n_288__51_, r_n_288__50_, r_n_288__49_, r_n_288__48_, r_n_288__47_, r_n_288__46_, r_n_288__45_, r_n_288__44_, r_n_288__43_, r_n_288__42_, r_n_288__41_, r_n_288__40_, r_n_288__39_, r_n_288__38_, r_n_288__37_, r_n_288__36_, r_n_288__35_, r_n_288__34_, r_n_288__33_, r_n_288__32_, r_n_288__31_, r_n_288__30_, r_n_288__29_, r_n_288__28_, r_n_288__27_, r_n_288__26_, r_n_288__25_, r_n_288__24_, r_n_288__23_, r_n_288__22_, r_n_288__21_, r_n_288__20_, r_n_288__19_, r_n_288__18_, r_n_288__17_, r_n_288__16_, r_n_288__15_, r_n_288__14_, r_n_288__13_, r_n_288__12_, r_n_288__11_, r_n_288__10_, r_n_288__9_, r_n_288__8_, r_n_288__7_, r_n_288__6_, r_n_288__5_, r_n_288__4_, r_n_288__3_, r_n_288__2_, r_n_288__1_, r_n_288__0_ } = (N576)? { r_289__63_, r_289__62_, r_289__61_, r_289__60_, r_289__59_, r_289__58_, r_289__57_, r_289__56_, r_289__55_, r_289__54_, r_289__53_, r_289__52_, r_289__51_, r_289__50_, r_289__49_, r_289__48_, r_289__47_, r_289__46_, r_289__45_, r_289__44_, r_289__43_, r_289__42_, r_289__41_, r_289__40_, r_289__39_, r_289__38_, r_289__37_, r_289__36_, r_289__35_, r_289__34_, r_289__33_, r_289__32_, r_289__31_, r_289__30_, r_289__29_, r_289__28_, r_289__27_, r_289__26_, r_289__25_, r_289__24_, r_289__23_, r_289__22_, r_289__21_, r_289__20_, r_289__19_, r_289__18_, r_289__17_, r_289__16_, r_289__15_, r_289__14_, r_289__13_, r_289__12_, r_289__11_, r_289__10_, r_289__9_, r_289__8_, r_289__7_, r_289__6_, r_289__5_, r_289__4_, r_289__3_, r_289__2_, r_289__1_, r_289__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N577)? data_i : 1'b0;
  assign N576 = sel_i[576];
  assign N577 = N2468;
  assign { r_n_289__63_, r_n_289__62_, r_n_289__61_, r_n_289__60_, r_n_289__59_, r_n_289__58_, r_n_289__57_, r_n_289__56_, r_n_289__55_, r_n_289__54_, r_n_289__53_, r_n_289__52_, r_n_289__51_, r_n_289__50_, r_n_289__49_, r_n_289__48_, r_n_289__47_, r_n_289__46_, r_n_289__45_, r_n_289__44_, r_n_289__43_, r_n_289__42_, r_n_289__41_, r_n_289__40_, r_n_289__39_, r_n_289__38_, r_n_289__37_, r_n_289__36_, r_n_289__35_, r_n_289__34_, r_n_289__33_, r_n_289__32_, r_n_289__31_, r_n_289__30_, r_n_289__29_, r_n_289__28_, r_n_289__27_, r_n_289__26_, r_n_289__25_, r_n_289__24_, r_n_289__23_, r_n_289__22_, r_n_289__21_, r_n_289__20_, r_n_289__19_, r_n_289__18_, r_n_289__17_, r_n_289__16_, r_n_289__15_, r_n_289__14_, r_n_289__13_, r_n_289__12_, r_n_289__11_, r_n_289__10_, r_n_289__9_, r_n_289__8_, r_n_289__7_, r_n_289__6_, r_n_289__5_, r_n_289__4_, r_n_289__3_, r_n_289__2_, r_n_289__1_, r_n_289__0_ } = (N578)? { r_290__63_, r_290__62_, r_290__61_, r_290__60_, r_290__59_, r_290__58_, r_290__57_, r_290__56_, r_290__55_, r_290__54_, r_290__53_, r_290__52_, r_290__51_, r_290__50_, r_290__49_, r_290__48_, r_290__47_, r_290__46_, r_290__45_, r_290__44_, r_290__43_, r_290__42_, r_290__41_, r_290__40_, r_290__39_, r_290__38_, r_290__37_, r_290__36_, r_290__35_, r_290__34_, r_290__33_, r_290__32_, r_290__31_, r_290__30_, r_290__29_, r_290__28_, r_290__27_, r_290__26_, r_290__25_, r_290__24_, r_290__23_, r_290__22_, r_290__21_, r_290__20_, r_290__19_, r_290__18_, r_290__17_, r_290__16_, r_290__15_, r_290__14_, r_290__13_, r_290__12_, r_290__11_, r_290__10_, r_290__9_, r_290__8_, r_290__7_, r_290__6_, r_290__5_, r_290__4_, r_290__3_, r_290__2_, r_290__1_, r_290__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N579)? data_i : 1'b0;
  assign N578 = sel_i[578];
  assign N579 = N2473;
  assign { r_n_290__63_, r_n_290__62_, r_n_290__61_, r_n_290__60_, r_n_290__59_, r_n_290__58_, r_n_290__57_, r_n_290__56_, r_n_290__55_, r_n_290__54_, r_n_290__53_, r_n_290__52_, r_n_290__51_, r_n_290__50_, r_n_290__49_, r_n_290__48_, r_n_290__47_, r_n_290__46_, r_n_290__45_, r_n_290__44_, r_n_290__43_, r_n_290__42_, r_n_290__41_, r_n_290__40_, r_n_290__39_, r_n_290__38_, r_n_290__37_, r_n_290__36_, r_n_290__35_, r_n_290__34_, r_n_290__33_, r_n_290__32_, r_n_290__31_, r_n_290__30_, r_n_290__29_, r_n_290__28_, r_n_290__27_, r_n_290__26_, r_n_290__25_, r_n_290__24_, r_n_290__23_, r_n_290__22_, r_n_290__21_, r_n_290__20_, r_n_290__19_, r_n_290__18_, r_n_290__17_, r_n_290__16_, r_n_290__15_, r_n_290__14_, r_n_290__13_, r_n_290__12_, r_n_290__11_, r_n_290__10_, r_n_290__9_, r_n_290__8_, r_n_290__7_, r_n_290__6_, r_n_290__5_, r_n_290__4_, r_n_290__3_, r_n_290__2_, r_n_290__1_, r_n_290__0_ } = (N580)? { r_291__63_, r_291__62_, r_291__61_, r_291__60_, r_291__59_, r_291__58_, r_291__57_, r_291__56_, r_291__55_, r_291__54_, r_291__53_, r_291__52_, r_291__51_, r_291__50_, r_291__49_, r_291__48_, r_291__47_, r_291__46_, r_291__45_, r_291__44_, r_291__43_, r_291__42_, r_291__41_, r_291__40_, r_291__39_, r_291__38_, r_291__37_, r_291__36_, r_291__35_, r_291__34_, r_291__33_, r_291__32_, r_291__31_, r_291__30_, r_291__29_, r_291__28_, r_291__27_, r_291__26_, r_291__25_, r_291__24_, r_291__23_, r_291__22_, r_291__21_, r_291__20_, r_291__19_, r_291__18_, r_291__17_, r_291__16_, r_291__15_, r_291__14_, r_291__13_, r_291__12_, r_291__11_, r_291__10_, r_291__9_, r_291__8_, r_291__7_, r_291__6_, r_291__5_, r_291__4_, r_291__3_, r_291__2_, r_291__1_, r_291__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N581)? data_i : 1'b0;
  assign N580 = sel_i[580];
  assign N581 = N2478;
  assign { r_n_291__63_, r_n_291__62_, r_n_291__61_, r_n_291__60_, r_n_291__59_, r_n_291__58_, r_n_291__57_, r_n_291__56_, r_n_291__55_, r_n_291__54_, r_n_291__53_, r_n_291__52_, r_n_291__51_, r_n_291__50_, r_n_291__49_, r_n_291__48_, r_n_291__47_, r_n_291__46_, r_n_291__45_, r_n_291__44_, r_n_291__43_, r_n_291__42_, r_n_291__41_, r_n_291__40_, r_n_291__39_, r_n_291__38_, r_n_291__37_, r_n_291__36_, r_n_291__35_, r_n_291__34_, r_n_291__33_, r_n_291__32_, r_n_291__31_, r_n_291__30_, r_n_291__29_, r_n_291__28_, r_n_291__27_, r_n_291__26_, r_n_291__25_, r_n_291__24_, r_n_291__23_, r_n_291__22_, r_n_291__21_, r_n_291__20_, r_n_291__19_, r_n_291__18_, r_n_291__17_, r_n_291__16_, r_n_291__15_, r_n_291__14_, r_n_291__13_, r_n_291__12_, r_n_291__11_, r_n_291__10_, r_n_291__9_, r_n_291__8_, r_n_291__7_, r_n_291__6_, r_n_291__5_, r_n_291__4_, r_n_291__3_, r_n_291__2_, r_n_291__1_, r_n_291__0_ } = (N582)? { r_292__63_, r_292__62_, r_292__61_, r_292__60_, r_292__59_, r_292__58_, r_292__57_, r_292__56_, r_292__55_, r_292__54_, r_292__53_, r_292__52_, r_292__51_, r_292__50_, r_292__49_, r_292__48_, r_292__47_, r_292__46_, r_292__45_, r_292__44_, r_292__43_, r_292__42_, r_292__41_, r_292__40_, r_292__39_, r_292__38_, r_292__37_, r_292__36_, r_292__35_, r_292__34_, r_292__33_, r_292__32_, r_292__31_, r_292__30_, r_292__29_, r_292__28_, r_292__27_, r_292__26_, r_292__25_, r_292__24_, r_292__23_, r_292__22_, r_292__21_, r_292__20_, r_292__19_, r_292__18_, r_292__17_, r_292__16_, r_292__15_, r_292__14_, r_292__13_, r_292__12_, r_292__11_, r_292__10_, r_292__9_, r_292__8_, r_292__7_, r_292__6_, r_292__5_, r_292__4_, r_292__3_, r_292__2_, r_292__1_, r_292__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N583)? data_i : 1'b0;
  assign N582 = sel_i[582];
  assign N583 = N2483;
  assign { r_n_292__63_, r_n_292__62_, r_n_292__61_, r_n_292__60_, r_n_292__59_, r_n_292__58_, r_n_292__57_, r_n_292__56_, r_n_292__55_, r_n_292__54_, r_n_292__53_, r_n_292__52_, r_n_292__51_, r_n_292__50_, r_n_292__49_, r_n_292__48_, r_n_292__47_, r_n_292__46_, r_n_292__45_, r_n_292__44_, r_n_292__43_, r_n_292__42_, r_n_292__41_, r_n_292__40_, r_n_292__39_, r_n_292__38_, r_n_292__37_, r_n_292__36_, r_n_292__35_, r_n_292__34_, r_n_292__33_, r_n_292__32_, r_n_292__31_, r_n_292__30_, r_n_292__29_, r_n_292__28_, r_n_292__27_, r_n_292__26_, r_n_292__25_, r_n_292__24_, r_n_292__23_, r_n_292__22_, r_n_292__21_, r_n_292__20_, r_n_292__19_, r_n_292__18_, r_n_292__17_, r_n_292__16_, r_n_292__15_, r_n_292__14_, r_n_292__13_, r_n_292__12_, r_n_292__11_, r_n_292__10_, r_n_292__9_, r_n_292__8_, r_n_292__7_, r_n_292__6_, r_n_292__5_, r_n_292__4_, r_n_292__3_, r_n_292__2_, r_n_292__1_, r_n_292__0_ } = (N584)? { r_293__63_, r_293__62_, r_293__61_, r_293__60_, r_293__59_, r_293__58_, r_293__57_, r_293__56_, r_293__55_, r_293__54_, r_293__53_, r_293__52_, r_293__51_, r_293__50_, r_293__49_, r_293__48_, r_293__47_, r_293__46_, r_293__45_, r_293__44_, r_293__43_, r_293__42_, r_293__41_, r_293__40_, r_293__39_, r_293__38_, r_293__37_, r_293__36_, r_293__35_, r_293__34_, r_293__33_, r_293__32_, r_293__31_, r_293__30_, r_293__29_, r_293__28_, r_293__27_, r_293__26_, r_293__25_, r_293__24_, r_293__23_, r_293__22_, r_293__21_, r_293__20_, r_293__19_, r_293__18_, r_293__17_, r_293__16_, r_293__15_, r_293__14_, r_293__13_, r_293__12_, r_293__11_, r_293__10_, r_293__9_, r_293__8_, r_293__7_, r_293__6_, r_293__5_, r_293__4_, r_293__3_, r_293__2_, r_293__1_, r_293__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N585)? data_i : 1'b0;
  assign N584 = sel_i[584];
  assign N585 = N2488;
  assign { r_n_293__63_, r_n_293__62_, r_n_293__61_, r_n_293__60_, r_n_293__59_, r_n_293__58_, r_n_293__57_, r_n_293__56_, r_n_293__55_, r_n_293__54_, r_n_293__53_, r_n_293__52_, r_n_293__51_, r_n_293__50_, r_n_293__49_, r_n_293__48_, r_n_293__47_, r_n_293__46_, r_n_293__45_, r_n_293__44_, r_n_293__43_, r_n_293__42_, r_n_293__41_, r_n_293__40_, r_n_293__39_, r_n_293__38_, r_n_293__37_, r_n_293__36_, r_n_293__35_, r_n_293__34_, r_n_293__33_, r_n_293__32_, r_n_293__31_, r_n_293__30_, r_n_293__29_, r_n_293__28_, r_n_293__27_, r_n_293__26_, r_n_293__25_, r_n_293__24_, r_n_293__23_, r_n_293__22_, r_n_293__21_, r_n_293__20_, r_n_293__19_, r_n_293__18_, r_n_293__17_, r_n_293__16_, r_n_293__15_, r_n_293__14_, r_n_293__13_, r_n_293__12_, r_n_293__11_, r_n_293__10_, r_n_293__9_, r_n_293__8_, r_n_293__7_, r_n_293__6_, r_n_293__5_, r_n_293__4_, r_n_293__3_, r_n_293__2_, r_n_293__1_, r_n_293__0_ } = (N586)? { r_294__63_, r_294__62_, r_294__61_, r_294__60_, r_294__59_, r_294__58_, r_294__57_, r_294__56_, r_294__55_, r_294__54_, r_294__53_, r_294__52_, r_294__51_, r_294__50_, r_294__49_, r_294__48_, r_294__47_, r_294__46_, r_294__45_, r_294__44_, r_294__43_, r_294__42_, r_294__41_, r_294__40_, r_294__39_, r_294__38_, r_294__37_, r_294__36_, r_294__35_, r_294__34_, r_294__33_, r_294__32_, r_294__31_, r_294__30_, r_294__29_, r_294__28_, r_294__27_, r_294__26_, r_294__25_, r_294__24_, r_294__23_, r_294__22_, r_294__21_, r_294__20_, r_294__19_, r_294__18_, r_294__17_, r_294__16_, r_294__15_, r_294__14_, r_294__13_, r_294__12_, r_294__11_, r_294__10_, r_294__9_, r_294__8_, r_294__7_, r_294__6_, r_294__5_, r_294__4_, r_294__3_, r_294__2_, r_294__1_, r_294__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N587)? data_i : 1'b0;
  assign N586 = sel_i[586];
  assign N587 = N2493;
  assign { r_n_294__63_, r_n_294__62_, r_n_294__61_, r_n_294__60_, r_n_294__59_, r_n_294__58_, r_n_294__57_, r_n_294__56_, r_n_294__55_, r_n_294__54_, r_n_294__53_, r_n_294__52_, r_n_294__51_, r_n_294__50_, r_n_294__49_, r_n_294__48_, r_n_294__47_, r_n_294__46_, r_n_294__45_, r_n_294__44_, r_n_294__43_, r_n_294__42_, r_n_294__41_, r_n_294__40_, r_n_294__39_, r_n_294__38_, r_n_294__37_, r_n_294__36_, r_n_294__35_, r_n_294__34_, r_n_294__33_, r_n_294__32_, r_n_294__31_, r_n_294__30_, r_n_294__29_, r_n_294__28_, r_n_294__27_, r_n_294__26_, r_n_294__25_, r_n_294__24_, r_n_294__23_, r_n_294__22_, r_n_294__21_, r_n_294__20_, r_n_294__19_, r_n_294__18_, r_n_294__17_, r_n_294__16_, r_n_294__15_, r_n_294__14_, r_n_294__13_, r_n_294__12_, r_n_294__11_, r_n_294__10_, r_n_294__9_, r_n_294__8_, r_n_294__7_, r_n_294__6_, r_n_294__5_, r_n_294__4_, r_n_294__3_, r_n_294__2_, r_n_294__1_, r_n_294__0_ } = (N588)? { r_295__63_, r_295__62_, r_295__61_, r_295__60_, r_295__59_, r_295__58_, r_295__57_, r_295__56_, r_295__55_, r_295__54_, r_295__53_, r_295__52_, r_295__51_, r_295__50_, r_295__49_, r_295__48_, r_295__47_, r_295__46_, r_295__45_, r_295__44_, r_295__43_, r_295__42_, r_295__41_, r_295__40_, r_295__39_, r_295__38_, r_295__37_, r_295__36_, r_295__35_, r_295__34_, r_295__33_, r_295__32_, r_295__31_, r_295__30_, r_295__29_, r_295__28_, r_295__27_, r_295__26_, r_295__25_, r_295__24_, r_295__23_, r_295__22_, r_295__21_, r_295__20_, r_295__19_, r_295__18_, r_295__17_, r_295__16_, r_295__15_, r_295__14_, r_295__13_, r_295__12_, r_295__11_, r_295__10_, r_295__9_, r_295__8_, r_295__7_, r_295__6_, r_295__5_, r_295__4_, r_295__3_, r_295__2_, r_295__1_, r_295__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N589)? data_i : 1'b0;
  assign N588 = sel_i[588];
  assign N589 = N2498;
  assign { r_n_295__63_, r_n_295__62_, r_n_295__61_, r_n_295__60_, r_n_295__59_, r_n_295__58_, r_n_295__57_, r_n_295__56_, r_n_295__55_, r_n_295__54_, r_n_295__53_, r_n_295__52_, r_n_295__51_, r_n_295__50_, r_n_295__49_, r_n_295__48_, r_n_295__47_, r_n_295__46_, r_n_295__45_, r_n_295__44_, r_n_295__43_, r_n_295__42_, r_n_295__41_, r_n_295__40_, r_n_295__39_, r_n_295__38_, r_n_295__37_, r_n_295__36_, r_n_295__35_, r_n_295__34_, r_n_295__33_, r_n_295__32_, r_n_295__31_, r_n_295__30_, r_n_295__29_, r_n_295__28_, r_n_295__27_, r_n_295__26_, r_n_295__25_, r_n_295__24_, r_n_295__23_, r_n_295__22_, r_n_295__21_, r_n_295__20_, r_n_295__19_, r_n_295__18_, r_n_295__17_, r_n_295__16_, r_n_295__15_, r_n_295__14_, r_n_295__13_, r_n_295__12_, r_n_295__11_, r_n_295__10_, r_n_295__9_, r_n_295__8_, r_n_295__7_, r_n_295__6_, r_n_295__5_, r_n_295__4_, r_n_295__3_, r_n_295__2_, r_n_295__1_, r_n_295__0_ } = (N590)? { r_296__63_, r_296__62_, r_296__61_, r_296__60_, r_296__59_, r_296__58_, r_296__57_, r_296__56_, r_296__55_, r_296__54_, r_296__53_, r_296__52_, r_296__51_, r_296__50_, r_296__49_, r_296__48_, r_296__47_, r_296__46_, r_296__45_, r_296__44_, r_296__43_, r_296__42_, r_296__41_, r_296__40_, r_296__39_, r_296__38_, r_296__37_, r_296__36_, r_296__35_, r_296__34_, r_296__33_, r_296__32_, r_296__31_, r_296__30_, r_296__29_, r_296__28_, r_296__27_, r_296__26_, r_296__25_, r_296__24_, r_296__23_, r_296__22_, r_296__21_, r_296__20_, r_296__19_, r_296__18_, r_296__17_, r_296__16_, r_296__15_, r_296__14_, r_296__13_, r_296__12_, r_296__11_, r_296__10_, r_296__9_, r_296__8_, r_296__7_, r_296__6_, r_296__5_, r_296__4_, r_296__3_, r_296__2_, r_296__1_, r_296__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N591)? data_i : 1'b0;
  assign N590 = sel_i[590];
  assign N591 = N2503;
  assign { r_n_296__63_, r_n_296__62_, r_n_296__61_, r_n_296__60_, r_n_296__59_, r_n_296__58_, r_n_296__57_, r_n_296__56_, r_n_296__55_, r_n_296__54_, r_n_296__53_, r_n_296__52_, r_n_296__51_, r_n_296__50_, r_n_296__49_, r_n_296__48_, r_n_296__47_, r_n_296__46_, r_n_296__45_, r_n_296__44_, r_n_296__43_, r_n_296__42_, r_n_296__41_, r_n_296__40_, r_n_296__39_, r_n_296__38_, r_n_296__37_, r_n_296__36_, r_n_296__35_, r_n_296__34_, r_n_296__33_, r_n_296__32_, r_n_296__31_, r_n_296__30_, r_n_296__29_, r_n_296__28_, r_n_296__27_, r_n_296__26_, r_n_296__25_, r_n_296__24_, r_n_296__23_, r_n_296__22_, r_n_296__21_, r_n_296__20_, r_n_296__19_, r_n_296__18_, r_n_296__17_, r_n_296__16_, r_n_296__15_, r_n_296__14_, r_n_296__13_, r_n_296__12_, r_n_296__11_, r_n_296__10_, r_n_296__9_, r_n_296__8_, r_n_296__7_, r_n_296__6_, r_n_296__5_, r_n_296__4_, r_n_296__3_, r_n_296__2_, r_n_296__1_, r_n_296__0_ } = (N592)? { r_297__63_, r_297__62_, r_297__61_, r_297__60_, r_297__59_, r_297__58_, r_297__57_, r_297__56_, r_297__55_, r_297__54_, r_297__53_, r_297__52_, r_297__51_, r_297__50_, r_297__49_, r_297__48_, r_297__47_, r_297__46_, r_297__45_, r_297__44_, r_297__43_, r_297__42_, r_297__41_, r_297__40_, r_297__39_, r_297__38_, r_297__37_, r_297__36_, r_297__35_, r_297__34_, r_297__33_, r_297__32_, r_297__31_, r_297__30_, r_297__29_, r_297__28_, r_297__27_, r_297__26_, r_297__25_, r_297__24_, r_297__23_, r_297__22_, r_297__21_, r_297__20_, r_297__19_, r_297__18_, r_297__17_, r_297__16_, r_297__15_, r_297__14_, r_297__13_, r_297__12_, r_297__11_, r_297__10_, r_297__9_, r_297__8_, r_297__7_, r_297__6_, r_297__5_, r_297__4_, r_297__3_, r_297__2_, r_297__1_, r_297__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N593)? data_i : 1'b0;
  assign N592 = sel_i[592];
  assign N593 = N2508;
  assign { r_n_297__63_, r_n_297__62_, r_n_297__61_, r_n_297__60_, r_n_297__59_, r_n_297__58_, r_n_297__57_, r_n_297__56_, r_n_297__55_, r_n_297__54_, r_n_297__53_, r_n_297__52_, r_n_297__51_, r_n_297__50_, r_n_297__49_, r_n_297__48_, r_n_297__47_, r_n_297__46_, r_n_297__45_, r_n_297__44_, r_n_297__43_, r_n_297__42_, r_n_297__41_, r_n_297__40_, r_n_297__39_, r_n_297__38_, r_n_297__37_, r_n_297__36_, r_n_297__35_, r_n_297__34_, r_n_297__33_, r_n_297__32_, r_n_297__31_, r_n_297__30_, r_n_297__29_, r_n_297__28_, r_n_297__27_, r_n_297__26_, r_n_297__25_, r_n_297__24_, r_n_297__23_, r_n_297__22_, r_n_297__21_, r_n_297__20_, r_n_297__19_, r_n_297__18_, r_n_297__17_, r_n_297__16_, r_n_297__15_, r_n_297__14_, r_n_297__13_, r_n_297__12_, r_n_297__11_, r_n_297__10_, r_n_297__9_, r_n_297__8_, r_n_297__7_, r_n_297__6_, r_n_297__5_, r_n_297__4_, r_n_297__3_, r_n_297__2_, r_n_297__1_, r_n_297__0_ } = (N594)? { r_298__63_, r_298__62_, r_298__61_, r_298__60_, r_298__59_, r_298__58_, r_298__57_, r_298__56_, r_298__55_, r_298__54_, r_298__53_, r_298__52_, r_298__51_, r_298__50_, r_298__49_, r_298__48_, r_298__47_, r_298__46_, r_298__45_, r_298__44_, r_298__43_, r_298__42_, r_298__41_, r_298__40_, r_298__39_, r_298__38_, r_298__37_, r_298__36_, r_298__35_, r_298__34_, r_298__33_, r_298__32_, r_298__31_, r_298__30_, r_298__29_, r_298__28_, r_298__27_, r_298__26_, r_298__25_, r_298__24_, r_298__23_, r_298__22_, r_298__21_, r_298__20_, r_298__19_, r_298__18_, r_298__17_, r_298__16_, r_298__15_, r_298__14_, r_298__13_, r_298__12_, r_298__11_, r_298__10_, r_298__9_, r_298__8_, r_298__7_, r_298__6_, r_298__5_, r_298__4_, r_298__3_, r_298__2_, r_298__1_, r_298__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N595)? data_i : 1'b0;
  assign N594 = sel_i[594];
  assign N595 = N2513;
  assign { r_n_298__63_, r_n_298__62_, r_n_298__61_, r_n_298__60_, r_n_298__59_, r_n_298__58_, r_n_298__57_, r_n_298__56_, r_n_298__55_, r_n_298__54_, r_n_298__53_, r_n_298__52_, r_n_298__51_, r_n_298__50_, r_n_298__49_, r_n_298__48_, r_n_298__47_, r_n_298__46_, r_n_298__45_, r_n_298__44_, r_n_298__43_, r_n_298__42_, r_n_298__41_, r_n_298__40_, r_n_298__39_, r_n_298__38_, r_n_298__37_, r_n_298__36_, r_n_298__35_, r_n_298__34_, r_n_298__33_, r_n_298__32_, r_n_298__31_, r_n_298__30_, r_n_298__29_, r_n_298__28_, r_n_298__27_, r_n_298__26_, r_n_298__25_, r_n_298__24_, r_n_298__23_, r_n_298__22_, r_n_298__21_, r_n_298__20_, r_n_298__19_, r_n_298__18_, r_n_298__17_, r_n_298__16_, r_n_298__15_, r_n_298__14_, r_n_298__13_, r_n_298__12_, r_n_298__11_, r_n_298__10_, r_n_298__9_, r_n_298__8_, r_n_298__7_, r_n_298__6_, r_n_298__5_, r_n_298__4_, r_n_298__3_, r_n_298__2_, r_n_298__1_, r_n_298__0_ } = (N596)? { r_299__63_, r_299__62_, r_299__61_, r_299__60_, r_299__59_, r_299__58_, r_299__57_, r_299__56_, r_299__55_, r_299__54_, r_299__53_, r_299__52_, r_299__51_, r_299__50_, r_299__49_, r_299__48_, r_299__47_, r_299__46_, r_299__45_, r_299__44_, r_299__43_, r_299__42_, r_299__41_, r_299__40_, r_299__39_, r_299__38_, r_299__37_, r_299__36_, r_299__35_, r_299__34_, r_299__33_, r_299__32_, r_299__31_, r_299__30_, r_299__29_, r_299__28_, r_299__27_, r_299__26_, r_299__25_, r_299__24_, r_299__23_, r_299__22_, r_299__21_, r_299__20_, r_299__19_, r_299__18_, r_299__17_, r_299__16_, r_299__15_, r_299__14_, r_299__13_, r_299__12_, r_299__11_, r_299__10_, r_299__9_, r_299__8_, r_299__7_, r_299__6_, r_299__5_, r_299__4_, r_299__3_, r_299__2_, r_299__1_, r_299__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N597)? data_i : 1'b0;
  assign N596 = sel_i[596];
  assign N597 = N2518;
  assign { r_n_299__63_, r_n_299__62_, r_n_299__61_, r_n_299__60_, r_n_299__59_, r_n_299__58_, r_n_299__57_, r_n_299__56_, r_n_299__55_, r_n_299__54_, r_n_299__53_, r_n_299__52_, r_n_299__51_, r_n_299__50_, r_n_299__49_, r_n_299__48_, r_n_299__47_, r_n_299__46_, r_n_299__45_, r_n_299__44_, r_n_299__43_, r_n_299__42_, r_n_299__41_, r_n_299__40_, r_n_299__39_, r_n_299__38_, r_n_299__37_, r_n_299__36_, r_n_299__35_, r_n_299__34_, r_n_299__33_, r_n_299__32_, r_n_299__31_, r_n_299__30_, r_n_299__29_, r_n_299__28_, r_n_299__27_, r_n_299__26_, r_n_299__25_, r_n_299__24_, r_n_299__23_, r_n_299__22_, r_n_299__21_, r_n_299__20_, r_n_299__19_, r_n_299__18_, r_n_299__17_, r_n_299__16_, r_n_299__15_, r_n_299__14_, r_n_299__13_, r_n_299__12_, r_n_299__11_, r_n_299__10_, r_n_299__9_, r_n_299__8_, r_n_299__7_, r_n_299__6_, r_n_299__5_, r_n_299__4_, r_n_299__3_, r_n_299__2_, r_n_299__1_, r_n_299__0_ } = (N598)? { r_300__63_, r_300__62_, r_300__61_, r_300__60_, r_300__59_, r_300__58_, r_300__57_, r_300__56_, r_300__55_, r_300__54_, r_300__53_, r_300__52_, r_300__51_, r_300__50_, r_300__49_, r_300__48_, r_300__47_, r_300__46_, r_300__45_, r_300__44_, r_300__43_, r_300__42_, r_300__41_, r_300__40_, r_300__39_, r_300__38_, r_300__37_, r_300__36_, r_300__35_, r_300__34_, r_300__33_, r_300__32_, r_300__31_, r_300__30_, r_300__29_, r_300__28_, r_300__27_, r_300__26_, r_300__25_, r_300__24_, r_300__23_, r_300__22_, r_300__21_, r_300__20_, r_300__19_, r_300__18_, r_300__17_, r_300__16_, r_300__15_, r_300__14_, r_300__13_, r_300__12_, r_300__11_, r_300__10_, r_300__9_, r_300__8_, r_300__7_, r_300__6_, r_300__5_, r_300__4_, r_300__3_, r_300__2_, r_300__1_, r_300__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N599)? data_i : 1'b0;
  assign N598 = sel_i[598];
  assign N599 = N2523;
  assign { r_n_300__63_, r_n_300__62_, r_n_300__61_, r_n_300__60_, r_n_300__59_, r_n_300__58_, r_n_300__57_, r_n_300__56_, r_n_300__55_, r_n_300__54_, r_n_300__53_, r_n_300__52_, r_n_300__51_, r_n_300__50_, r_n_300__49_, r_n_300__48_, r_n_300__47_, r_n_300__46_, r_n_300__45_, r_n_300__44_, r_n_300__43_, r_n_300__42_, r_n_300__41_, r_n_300__40_, r_n_300__39_, r_n_300__38_, r_n_300__37_, r_n_300__36_, r_n_300__35_, r_n_300__34_, r_n_300__33_, r_n_300__32_, r_n_300__31_, r_n_300__30_, r_n_300__29_, r_n_300__28_, r_n_300__27_, r_n_300__26_, r_n_300__25_, r_n_300__24_, r_n_300__23_, r_n_300__22_, r_n_300__21_, r_n_300__20_, r_n_300__19_, r_n_300__18_, r_n_300__17_, r_n_300__16_, r_n_300__15_, r_n_300__14_, r_n_300__13_, r_n_300__12_, r_n_300__11_, r_n_300__10_, r_n_300__9_, r_n_300__8_, r_n_300__7_, r_n_300__6_, r_n_300__5_, r_n_300__4_, r_n_300__3_, r_n_300__2_, r_n_300__1_, r_n_300__0_ } = (N600)? { r_301__63_, r_301__62_, r_301__61_, r_301__60_, r_301__59_, r_301__58_, r_301__57_, r_301__56_, r_301__55_, r_301__54_, r_301__53_, r_301__52_, r_301__51_, r_301__50_, r_301__49_, r_301__48_, r_301__47_, r_301__46_, r_301__45_, r_301__44_, r_301__43_, r_301__42_, r_301__41_, r_301__40_, r_301__39_, r_301__38_, r_301__37_, r_301__36_, r_301__35_, r_301__34_, r_301__33_, r_301__32_, r_301__31_, r_301__30_, r_301__29_, r_301__28_, r_301__27_, r_301__26_, r_301__25_, r_301__24_, r_301__23_, r_301__22_, r_301__21_, r_301__20_, r_301__19_, r_301__18_, r_301__17_, r_301__16_, r_301__15_, r_301__14_, r_301__13_, r_301__12_, r_301__11_, r_301__10_, r_301__9_, r_301__8_, r_301__7_, r_301__6_, r_301__5_, r_301__4_, r_301__3_, r_301__2_, r_301__1_, r_301__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N601)? data_i : 1'b0;
  assign N600 = sel_i[600];
  assign N601 = N2528;
  assign { r_n_301__63_, r_n_301__62_, r_n_301__61_, r_n_301__60_, r_n_301__59_, r_n_301__58_, r_n_301__57_, r_n_301__56_, r_n_301__55_, r_n_301__54_, r_n_301__53_, r_n_301__52_, r_n_301__51_, r_n_301__50_, r_n_301__49_, r_n_301__48_, r_n_301__47_, r_n_301__46_, r_n_301__45_, r_n_301__44_, r_n_301__43_, r_n_301__42_, r_n_301__41_, r_n_301__40_, r_n_301__39_, r_n_301__38_, r_n_301__37_, r_n_301__36_, r_n_301__35_, r_n_301__34_, r_n_301__33_, r_n_301__32_, r_n_301__31_, r_n_301__30_, r_n_301__29_, r_n_301__28_, r_n_301__27_, r_n_301__26_, r_n_301__25_, r_n_301__24_, r_n_301__23_, r_n_301__22_, r_n_301__21_, r_n_301__20_, r_n_301__19_, r_n_301__18_, r_n_301__17_, r_n_301__16_, r_n_301__15_, r_n_301__14_, r_n_301__13_, r_n_301__12_, r_n_301__11_, r_n_301__10_, r_n_301__9_, r_n_301__8_, r_n_301__7_, r_n_301__6_, r_n_301__5_, r_n_301__4_, r_n_301__3_, r_n_301__2_, r_n_301__1_, r_n_301__0_ } = (N602)? { r_302__63_, r_302__62_, r_302__61_, r_302__60_, r_302__59_, r_302__58_, r_302__57_, r_302__56_, r_302__55_, r_302__54_, r_302__53_, r_302__52_, r_302__51_, r_302__50_, r_302__49_, r_302__48_, r_302__47_, r_302__46_, r_302__45_, r_302__44_, r_302__43_, r_302__42_, r_302__41_, r_302__40_, r_302__39_, r_302__38_, r_302__37_, r_302__36_, r_302__35_, r_302__34_, r_302__33_, r_302__32_, r_302__31_, r_302__30_, r_302__29_, r_302__28_, r_302__27_, r_302__26_, r_302__25_, r_302__24_, r_302__23_, r_302__22_, r_302__21_, r_302__20_, r_302__19_, r_302__18_, r_302__17_, r_302__16_, r_302__15_, r_302__14_, r_302__13_, r_302__12_, r_302__11_, r_302__10_, r_302__9_, r_302__8_, r_302__7_, r_302__6_, r_302__5_, r_302__4_, r_302__3_, r_302__2_, r_302__1_, r_302__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N603)? data_i : 1'b0;
  assign N602 = sel_i[602];
  assign N603 = N2533;
  assign { r_n_302__63_, r_n_302__62_, r_n_302__61_, r_n_302__60_, r_n_302__59_, r_n_302__58_, r_n_302__57_, r_n_302__56_, r_n_302__55_, r_n_302__54_, r_n_302__53_, r_n_302__52_, r_n_302__51_, r_n_302__50_, r_n_302__49_, r_n_302__48_, r_n_302__47_, r_n_302__46_, r_n_302__45_, r_n_302__44_, r_n_302__43_, r_n_302__42_, r_n_302__41_, r_n_302__40_, r_n_302__39_, r_n_302__38_, r_n_302__37_, r_n_302__36_, r_n_302__35_, r_n_302__34_, r_n_302__33_, r_n_302__32_, r_n_302__31_, r_n_302__30_, r_n_302__29_, r_n_302__28_, r_n_302__27_, r_n_302__26_, r_n_302__25_, r_n_302__24_, r_n_302__23_, r_n_302__22_, r_n_302__21_, r_n_302__20_, r_n_302__19_, r_n_302__18_, r_n_302__17_, r_n_302__16_, r_n_302__15_, r_n_302__14_, r_n_302__13_, r_n_302__12_, r_n_302__11_, r_n_302__10_, r_n_302__9_, r_n_302__8_, r_n_302__7_, r_n_302__6_, r_n_302__5_, r_n_302__4_, r_n_302__3_, r_n_302__2_, r_n_302__1_, r_n_302__0_ } = (N604)? { r_303__63_, r_303__62_, r_303__61_, r_303__60_, r_303__59_, r_303__58_, r_303__57_, r_303__56_, r_303__55_, r_303__54_, r_303__53_, r_303__52_, r_303__51_, r_303__50_, r_303__49_, r_303__48_, r_303__47_, r_303__46_, r_303__45_, r_303__44_, r_303__43_, r_303__42_, r_303__41_, r_303__40_, r_303__39_, r_303__38_, r_303__37_, r_303__36_, r_303__35_, r_303__34_, r_303__33_, r_303__32_, r_303__31_, r_303__30_, r_303__29_, r_303__28_, r_303__27_, r_303__26_, r_303__25_, r_303__24_, r_303__23_, r_303__22_, r_303__21_, r_303__20_, r_303__19_, r_303__18_, r_303__17_, r_303__16_, r_303__15_, r_303__14_, r_303__13_, r_303__12_, r_303__11_, r_303__10_, r_303__9_, r_303__8_, r_303__7_, r_303__6_, r_303__5_, r_303__4_, r_303__3_, r_303__2_, r_303__1_, r_303__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N605)? data_i : 1'b0;
  assign N604 = sel_i[604];
  assign N605 = N2538;
  assign { r_n_303__63_, r_n_303__62_, r_n_303__61_, r_n_303__60_, r_n_303__59_, r_n_303__58_, r_n_303__57_, r_n_303__56_, r_n_303__55_, r_n_303__54_, r_n_303__53_, r_n_303__52_, r_n_303__51_, r_n_303__50_, r_n_303__49_, r_n_303__48_, r_n_303__47_, r_n_303__46_, r_n_303__45_, r_n_303__44_, r_n_303__43_, r_n_303__42_, r_n_303__41_, r_n_303__40_, r_n_303__39_, r_n_303__38_, r_n_303__37_, r_n_303__36_, r_n_303__35_, r_n_303__34_, r_n_303__33_, r_n_303__32_, r_n_303__31_, r_n_303__30_, r_n_303__29_, r_n_303__28_, r_n_303__27_, r_n_303__26_, r_n_303__25_, r_n_303__24_, r_n_303__23_, r_n_303__22_, r_n_303__21_, r_n_303__20_, r_n_303__19_, r_n_303__18_, r_n_303__17_, r_n_303__16_, r_n_303__15_, r_n_303__14_, r_n_303__13_, r_n_303__12_, r_n_303__11_, r_n_303__10_, r_n_303__9_, r_n_303__8_, r_n_303__7_, r_n_303__6_, r_n_303__5_, r_n_303__4_, r_n_303__3_, r_n_303__2_, r_n_303__1_, r_n_303__0_ } = (N606)? { r_304__63_, r_304__62_, r_304__61_, r_304__60_, r_304__59_, r_304__58_, r_304__57_, r_304__56_, r_304__55_, r_304__54_, r_304__53_, r_304__52_, r_304__51_, r_304__50_, r_304__49_, r_304__48_, r_304__47_, r_304__46_, r_304__45_, r_304__44_, r_304__43_, r_304__42_, r_304__41_, r_304__40_, r_304__39_, r_304__38_, r_304__37_, r_304__36_, r_304__35_, r_304__34_, r_304__33_, r_304__32_, r_304__31_, r_304__30_, r_304__29_, r_304__28_, r_304__27_, r_304__26_, r_304__25_, r_304__24_, r_304__23_, r_304__22_, r_304__21_, r_304__20_, r_304__19_, r_304__18_, r_304__17_, r_304__16_, r_304__15_, r_304__14_, r_304__13_, r_304__12_, r_304__11_, r_304__10_, r_304__9_, r_304__8_, r_304__7_, r_304__6_, r_304__5_, r_304__4_, r_304__3_, r_304__2_, r_304__1_, r_304__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N607)? data_i : 1'b0;
  assign N606 = sel_i[606];
  assign N607 = N2543;
  assign { r_n_304__63_, r_n_304__62_, r_n_304__61_, r_n_304__60_, r_n_304__59_, r_n_304__58_, r_n_304__57_, r_n_304__56_, r_n_304__55_, r_n_304__54_, r_n_304__53_, r_n_304__52_, r_n_304__51_, r_n_304__50_, r_n_304__49_, r_n_304__48_, r_n_304__47_, r_n_304__46_, r_n_304__45_, r_n_304__44_, r_n_304__43_, r_n_304__42_, r_n_304__41_, r_n_304__40_, r_n_304__39_, r_n_304__38_, r_n_304__37_, r_n_304__36_, r_n_304__35_, r_n_304__34_, r_n_304__33_, r_n_304__32_, r_n_304__31_, r_n_304__30_, r_n_304__29_, r_n_304__28_, r_n_304__27_, r_n_304__26_, r_n_304__25_, r_n_304__24_, r_n_304__23_, r_n_304__22_, r_n_304__21_, r_n_304__20_, r_n_304__19_, r_n_304__18_, r_n_304__17_, r_n_304__16_, r_n_304__15_, r_n_304__14_, r_n_304__13_, r_n_304__12_, r_n_304__11_, r_n_304__10_, r_n_304__9_, r_n_304__8_, r_n_304__7_, r_n_304__6_, r_n_304__5_, r_n_304__4_, r_n_304__3_, r_n_304__2_, r_n_304__1_, r_n_304__0_ } = (N608)? { r_305__63_, r_305__62_, r_305__61_, r_305__60_, r_305__59_, r_305__58_, r_305__57_, r_305__56_, r_305__55_, r_305__54_, r_305__53_, r_305__52_, r_305__51_, r_305__50_, r_305__49_, r_305__48_, r_305__47_, r_305__46_, r_305__45_, r_305__44_, r_305__43_, r_305__42_, r_305__41_, r_305__40_, r_305__39_, r_305__38_, r_305__37_, r_305__36_, r_305__35_, r_305__34_, r_305__33_, r_305__32_, r_305__31_, r_305__30_, r_305__29_, r_305__28_, r_305__27_, r_305__26_, r_305__25_, r_305__24_, r_305__23_, r_305__22_, r_305__21_, r_305__20_, r_305__19_, r_305__18_, r_305__17_, r_305__16_, r_305__15_, r_305__14_, r_305__13_, r_305__12_, r_305__11_, r_305__10_, r_305__9_, r_305__8_, r_305__7_, r_305__6_, r_305__5_, r_305__4_, r_305__3_, r_305__2_, r_305__1_, r_305__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N609)? data_i : 1'b0;
  assign N608 = sel_i[608];
  assign N609 = N2548;
  assign { r_n_305__63_, r_n_305__62_, r_n_305__61_, r_n_305__60_, r_n_305__59_, r_n_305__58_, r_n_305__57_, r_n_305__56_, r_n_305__55_, r_n_305__54_, r_n_305__53_, r_n_305__52_, r_n_305__51_, r_n_305__50_, r_n_305__49_, r_n_305__48_, r_n_305__47_, r_n_305__46_, r_n_305__45_, r_n_305__44_, r_n_305__43_, r_n_305__42_, r_n_305__41_, r_n_305__40_, r_n_305__39_, r_n_305__38_, r_n_305__37_, r_n_305__36_, r_n_305__35_, r_n_305__34_, r_n_305__33_, r_n_305__32_, r_n_305__31_, r_n_305__30_, r_n_305__29_, r_n_305__28_, r_n_305__27_, r_n_305__26_, r_n_305__25_, r_n_305__24_, r_n_305__23_, r_n_305__22_, r_n_305__21_, r_n_305__20_, r_n_305__19_, r_n_305__18_, r_n_305__17_, r_n_305__16_, r_n_305__15_, r_n_305__14_, r_n_305__13_, r_n_305__12_, r_n_305__11_, r_n_305__10_, r_n_305__9_, r_n_305__8_, r_n_305__7_, r_n_305__6_, r_n_305__5_, r_n_305__4_, r_n_305__3_, r_n_305__2_, r_n_305__1_, r_n_305__0_ } = (N610)? { r_306__63_, r_306__62_, r_306__61_, r_306__60_, r_306__59_, r_306__58_, r_306__57_, r_306__56_, r_306__55_, r_306__54_, r_306__53_, r_306__52_, r_306__51_, r_306__50_, r_306__49_, r_306__48_, r_306__47_, r_306__46_, r_306__45_, r_306__44_, r_306__43_, r_306__42_, r_306__41_, r_306__40_, r_306__39_, r_306__38_, r_306__37_, r_306__36_, r_306__35_, r_306__34_, r_306__33_, r_306__32_, r_306__31_, r_306__30_, r_306__29_, r_306__28_, r_306__27_, r_306__26_, r_306__25_, r_306__24_, r_306__23_, r_306__22_, r_306__21_, r_306__20_, r_306__19_, r_306__18_, r_306__17_, r_306__16_, r_306__15_, r_306__14_, r_306__13_, r_306__12_, r_306__11_, r_306__10_, r_306__9_, r_306__8_, r_306__7_, r_306__6_, r_306__5_, r_306__4_, r_306__3_, r_306__2_, r_306__1_, r_306__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N611)? data_i : 1'b0;
  assign N610 = sel_i[610];
  assign N611 = N2553;
  assign { r_n_306__63_, r_n_306__62_, r_n_306__61_, r_n_306__60_, r_n_306__59_, r_n_306__58_, r_n_306__57_, r_n_306__56_, r_n_306__55_, r_n_306__54_, r_n_306__53_, r_n_306__52_, r_n_306__51_, r_n_306__50_, r_n_306__49_, r_n_306__48_, r_n_306__47_, r_n_306__46_, r_n_306__45_, r_n_306__44_, r_n_306__43_, r_n_306__42_, r_n_306__41_, r_n_306__40_, r_n_306__39_, r_n_306__38_, r_n_306__37_, r_n_306__36_, r_n_306__35_, r_n_306__34_, r_n_306__33_, r_n_306__32_, r_n_306__31_, r_n_306__30_, r_n_306__29_, r_n_306__28_, r_n_306__27_, r_n_306__26_, r_n_306__25_, r_n_306__24_, r_n_306__23_, r_n_306__22_, r_n_306__21_, r_n_306__20_, r_n_306__19_, r_n_306__18_, r_n_306__17_, r_n_306__16_, r_n_306__15_, r_n_306__14_, r_n_306__13_, r_n_306__12_, r_n_306__11_, r_n_306__10_, r_n_306__9_, r_n_306__8_, r_n_306__7_, r_n_306__6_, r_n_306__5_, r_n_306__4_, r_n_306__3_, r_n_306__2_, r_n_306__1_, r_n_306__0_ } = (N612)? { r_307__63_, r_307__62_, r_307__61_, r_307__60_, r_307__59_, r_307__58_, r_307__57_, r_307__56_, r_307__55_, r_307__54_, r_307__53_, r_307__52_, r_307__51_, r_307__50_, r_307__49_, r_307__48_, r_307__47_, r_307__46_, r_307__45_, r_307__44_, r_307__43_, r_307__42_, r_307__41_, r_307__40_, r_307__39_, r_307__38_, r_307__37_, r_307__36_, r_307__35_, r_307__34_, r_307__33_, r_307__32_, r_307__31_, r_307__30_, r_307__29_, r_307__28_, r_307__27_, r_307__26_, r_307__25_, r_307__24_, r_307__23_, r_307__22_, r_307__21_, r_307__20_, r_307__19_, r_307__18_, r_307__17_, r_307__16_, r_307__15_, r_307__14_, r_307__13_, r_307__12_, r_307__11_, r_307__10_, r_307__9_, r_307__8_, r_307__7_, r_307__6_, r_307__5_, r_307__4_, r_307__3_, r_307__2_, r_307__1_, r_307__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N613)? data_i : 1'b0;
  assign N612 = sel_i[612];
  assign N613 = N2558;
  assign { r_n_307__63_, r_n_307__62_, r_n_307__61_, r_n_307__60_, r_n_307__59_, r_n_307__58_, r_n_307__57_, r_n_307__56_, r_n_307__55_, r_n_307__54_, r_n_307__53_, r_n_307__52_, r_n_307__51_, r_n_307__50_, r_n_307__49_, r_n_307__48_, r_n_307__47_, r_n_307__46_, r_n_307__45_, r_n_307__44_, r_n_307__43_, r_n_307__42_, r_n_307__41_, r_n_307__40_, r_n_307__39_, r_n_307__38_, r_n_307__37_, r_n_307__36_, r_n_307__35_, r_n_307__34_, r_n_307__33_, r_n_307__32_, r_n_307__31_, r_n_307__30_, r_n_307__29_, r_n_307__28_, r_n_307__27_, r_n_307__26_, r_n_307__25_, r_n_307__24_, r_n_307__23_, r_n_307__22_, r_n_307__21_, r_n_307__20_, r_n_307__19_, r_n_307__18_, r_n_307__17_, r_n_307__16_, r_n_307__15_, r_n_307__14_, r_n_307__13_, r_n_307__12_, r_n_307__11_, r_n_307__10_, r_n_307__9_, r_n_307__8_, r_n_307__7_, r_n_307__6_, r_n_307__5_, r_n_307__4_, r_n_307__3_, r_n_307__2_, r_n_307__1_, r_n_307__0_ } = (N614)? { r_308__63_, r_308__62_, r_308__61_, r_308__60_, r_308__59_, r_308__58_, r_308__57_, r_308__56_, r_308__55_, r_308__54_, r_308__53_, r_308__52_, r_308__51_, r_308__50_, r_308__49_, r_308__48_, r_308__47_, r_308__46_, r_308__45_, r_308__44_, r_308__43_, r_308__42_, r_308__41_, r_308__40_, r_308__39_, r_308__38_, r_308__37_, r_308__36_, r_308__35_, r_308__34_, r_308__33_, r_308__32_, r_308__31_, r_308__30_, r_308__29_, r_308__28_, r_308__27_, r_308__26_, r_308__25_, r_308__24_, r_308__23_, r_308__22_, r_308__21_, r_308__20_, r_308__19_, r_308__18_, r_308__17_, r_308__16_, r_308__15_, r_308__14_, r_308__13_, r_308__12_, r_308__11_, r_308__10_, r_308__9_, r_308__8_, r_308__7_, r_308__6_, r_308__5_, r_308__4_, r_308__3_, r_308__2_, r_308__1_, r_308__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N615)? data_i : 1'b0;
  assign N614 = sel_i[614];
  assign N615 = N2563;
  assign { r_n_308__63_, r_n_308__62_, r_n_308__61_, r_n_308__60_, r_n_308__59_, r_n_308__58_, r_n_308__57_, r_n_308__56_, r_n_308__55_, r_n_308__54_, r_n_308__53_, r_n_308__52_, r_n_308__51_, r_n_308__50_, r_n_308__49_, r_n_308__48_, r_n_308__47_, r_n_308__46_, r_n_308__45_, r_n_308__44_, r_n_308__43_, r_n_308__42_, r_n_308__41_, r_n_308__40_, r_n_308__39_, r_n_308__38_, r_n_308__37_, r_n_308__36_, r_n_308__35_, r_n_308__34_, r_n_308__33_, r_n_308__32_, r_n_308__31_, r_n_308__30_, r_n_308__29_, r_n_308__28_, r_n_308__27_, r_n_308__26_, r_n_308__25_, r_n_308__24_, r_n_308__23_, r_n_308__22_, r_n_308__21_, r_n_308__20_, r_n_308__19_, r_n_308__18_, r_n_308__17_, r_n_308__16_, r_n_308__15_, r_n_308__14_, r_n_308__13_, r_n_308__12_, r_n_308__11_, r_n_308__10_, r_n_308__9_, r_n_308__8_, r_n_308__7_, r_n_308__6_, r_n_308__5_, r_n_308__4_, r_n_308__3_, r_n_308__2_, r_n_308__1_, r_n_308__0_ } = (N616)? { r_309__63_, r_309__62_, r_309__61_, r_309__60_, r_309__59_, r_309__58_, r_309__57_, r_309__56_, r_309__55_, r_309__54_, r_309__53_, r_309__52_, r_309__51_, r_309__50_, r_309__49_, r_309__48_, r_309__47_, r_309__46_, r_309__45_, r_309__44_, r_309__43_, r_309__42_, r_309__41_, r_309__40_, r_309__39_, r_309__38_, r_309__37_, r_309__36_, r_309__35_, r_309__34_, r_309__33_, r_309__32_, r_309__31_, r_309__30_, r_309__29_, r_309__28_, r_309__27_, r_309__26_, r_309__25_, r_309__24_, r_309__23_, r_309__22_, r_309__21_, r_309__20_, r_309__19_, r_309__18_, r_309__17_, r_309__16_, r_309__15_, r_309__14_, r_309__13_, r_309__12_, r_309__11_, r_309__10_, r_309__9_, r_309__8_, r_309__7_, r_309__6_, r_309__5_, r_309__4_, r_309__3_, r_309__2_, r_309__1_, r_309__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N617)? data_i : 1'b0;
  assign N616 = sel_i[616];
  assign N617 = N2568;
  assign { r_n_309__63_, r_n_309__62_, r_n_309__61_, r_n_309__60_, r_n_309__59_, r_n_309__58_, r_n_309__57_, r_n_309__56_, r_n_309__55_, r_n_309__54_, r_n_309__53_, r_n_309__52_, r_n_309__51_, r_n_309__50_, r_n_309__49_, r_n_309__48_, r_n_309__47_, r_n_309__46_, r_n_309__45_, r_n_309__44_, r_n_309__43_, r_n_309__42_, r_n_309__41_, r_n_309__40_, r_n_309__39_, r_n_309__38_, r_n_309__37_, r_n_309__36_, r_n_309__35_, r_n_309__34_, r_n_309__33_, r_n_309__32_, r_n_309__31_, r_n_309__30_, r_n_309__29_, r_n_309__28_, r_n_309__27_, r_n_309__26_, r_n_309__25_, r_n_309__24_, r_n_309__23_, r_n_309__22_, r_n_309__21_, r_n_309__20_, r_n_309__19_, r_n_309__18_, r_n_309__17_, r_n_309__16_, r_n_309__15_, r_n_309__14_, r_n_309__13_, r_n_309__12_, r_n_309__11_, r_n_309__10_, r_n_309__9_, r_n_309__8_, r_n_309__7_, r_n_309__6_, r_n_309__5_, r_n_309__4_, r_n_309__3_, r_n_309__2_, r_n_309__1_, r_n_309__0_ } = (N618)? { r_310__63_, r_310__62_, r_310__61_, r_310__60_, r_310__59_, r_310__58_, r_310__57_, r_310__56_, r_310__55_, r_310__54_, r_310__53_, r_310__52_, r_310__51_, r_310__50_, r_310__49_, r_310__48_, r_310__47_, r_310__46_, r_310__45_, r_310__44_, r_310__43_, r_310__42_, r_310__41_, r_310__40_, r_310__39_, r_310__38_, r_310__37_, r_310__36_, r_310__35_, r_310__34_, r_310__33_, r_310__32_, r_310__31_, r_310__30_, r_310__29_, r_310__28_, r_310__27_, r_310__26_, r_310__25_, r_310__24_, r_310__23_, r_310__22_, r_310__21_, r_310__20_, r_310__19_, r_310__18_, r_310__17_, r_310__16_, r_310__15_, r_310__14_, r_310__13_, r_310__12_, r_310__11_, r_310__10_, r_310__9_, r_310__8_, r_310__7_, r_310__6_, r_310__5_, r_310__4_, r_310__3_, r_310__2_, r_310__1_, r_310__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N619)? data_i : 1'b0;
  assign N618 = sel_i[618];
  assign N619 = N2573;
  assign { r_n_310__63_, r_n_310__62_, r_n_310__61_, r_n_310__60_, r_n_310__59_, r_n_310__58_, r_n_310__57_, r_n_310__56_, r_n_310__55_, r_n_310__54_, r_n_310__53_, r_n_310__52_, r_n_310__51_, r_n_310__50_, r_n_310__49_, r_n_310__48_, r_n_310__47_, r_n_310__46_, r_n_310__45_, r_n_310__44_, r_n_310__43_, r_n_310__42_, r_n_310__41_, r_n_310__40_, r_n_310__39_, r_n_310__38_, r_n_310__37_, r_n_310__36_, r_n_310__35_, r_n_310__34_, r_n_310__33_, r_n_310__32_, r_n_310__31_, r_n_310__30_, r_n_310__29_, r_n_310__28_, r_n_310__27_, r_n_310__26_, r_n_310__25_, r_n_310__24_, r_n_310__23_, r_n_310__22_, r_n_310__21_, r_n_310__20_, r_n_310__19_, r_n_310__18_, r_n_310__17_, r_n_310__16_, r_n_310__15_, r_n_310__14_, r_n_310__13_, r_n_310__12_, r_n_310__11_, r_n_310__10_, r_n_310__9_, r_n_310__8_, r_n_310__7_, r_n_310__6_, r_n_310__5_, r_n_310__4_, r_n_310__3_, r_n_310__2_, r_n_310__1_, r_n_310__0_ } = (N620)? { r_311__63_, r_311__62_, r_311__61_, r_311__60_, r_311__59_, r_311__58_, r_311__57_, r_311__56_, r_311__55_, r_311__54_, r_311__53_, r_311__52_, r_311__51_, r_311__50_, r_311__49_, r_311__48_, r_311__47_, r_311__46_, r_311__45_, r_311__44_, r_311__43_, r_311__42_, r_311__41_, r_311__40_, r_311__39_, r_311__38_, r_311__37_, r_311__36_, r_311__35_, r_311__34_, r_311__33_, r_311__32_, r_311__31_, r_311__30_, r_311__29_, r_311__28_, r_311__27_, r_311__26_, r_311__25_, r_311__24_, r_311__23_, r_311__22_, r_311__21_, r_311__20_, r_311__19_, r_311__18_, r_311__17_, r_311__16_, r_311__15_, r_311__14_, r_311__13_, r_311__12_, r_311__11_, r_311__10_, r_311__9_, r_311__8_, r_311__7_, r_311__6_, r_311__5_, r_311__4_, r_311__3_, r_311__2_, r_311__1_, r_311__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N621)? data_i : 1'b0;
  assign N620 = sel_i[620];
  assign N621 = N2578;
  assign { r_n_311__63_, r_n_311__62_, r_n_311__61_, r_n_311__60_, r_n_311__59_, r_n_311__58_, r_n_311__57_, r_n_311__56_, r_n_311__55_, r_n_311__54_, r_n_311__53_, r_n_311__52_, r_n_311__51_, r_n_311__50_, r_n_311__49_, r_n_311__48_, r_n_311__47_, r_n_311__46_, r_n_311__45_, r_n_311__44_, r_n_311__43_, r_n_311__42_, r_n_311__41_, r_n_311__40_, r_n_311__39_, r_n_311__38_, r_n_311__37_, r_n_311__36_, r_n_311__35_, r_n_311__34_, r_n_311__33_, r_n_311__32_, r_n_311__31_, r_n_311__30_, r_n_311__29_, r_n_311__28_, r_n_311__27_, r_n_311__26_, r_n_311__25_, r_n_311__24_, r_n_311__23_, r_n_311__22_, r_n_311__21_, r_n_311__20_, r_n_311__19_, r_n_311__18_, r_n_311__17_, r_n_311__16_, r_n_311__15_, r_n_311__14_, r_n_311__13_, r_n_311__12_, r_n_311__11_, r_n_311__10_, r_n_311__9_, r_n_311__8_, r_n_311__7_, r_n_311__6_, r_n_311__5_, r_n_311__4_, r_n_311__3_, r_n_311__2_, r_n_311__1_, r_n_311__0_ } = (N622)? { r_312__63_, r_312__62_, r_312__61_, r_312__60_, r_312__59_, r_312__58_, r_312__57_, r_312__56_, r_312__55_, r_312__54_, r_312__53_, r_312__52_, r_312__51_, r_312__50_, r_312__49_, r_312__48_, r_312__47_, r_312__46_, r_312__45_, r_312__44_, r_312__43_, r_312__42_, r_312__41_, r_312__40_, r_312__39_, r_312__38_, r_312__37_, r_312__36_, r_312__35_, r_312__34_, r_312__33_, r_312__32_, r_312__31_, r_312__30_, r_312__29_, r_312__28_, r_312__27_, r_312__26_, r_312__25_, r_312__24_, r_312__23_, r_312__22_, r_312__21_, r_312__20_, r_312__19_, r_312__18_, r_312__17_, r_312__16_, r_312__15_, r_312__14_, r_312__13_, r_312__12_, r_312__11_, r_312__10_, r_312__9_, r_312__8_, r_312__7_, r_312__6_, r_312__5_, r_312__4_, r_312__3_, r_312__2_, r_312__1_, r_312__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N623)? data_i : 1'b0;
  assign N622 = sel_i[622];
  assign N623 = N2583;
  assign { r_n_312__63_, r_n_312__62_, r_n_312__61_, r_n_312__60_, r_n_312__59_, r_n_312__58_, r_n_312__57_, r_n_312__56_, r_n_312__55_, r_n_312__54_, r_n_312__53_, r_n_312__52_, r_n_312__51_, r_n_312__50_, r_n_312__49_, r_n_312__48_, r_n_312__47_, r_n_312__46_, r_n_312__45_, r_n_312__44_, r_n_312__43_, r_n_312__42_, r_n_312__41_, r_n_312__40_, r_n_312__39_, r_n_312__38_, r_n_312__37_, r_n_312__36_, r_n_312__35_, r_n_312__34_, r_n_312__33_, r_n_312__32_, r_n_312__31_, r_n_312__30_, r_n_312__29_, r_n_312__28_, r_n_312__27_, r_n_312__26_, r_n_312__25_, r_n_312__24_, r_n_312__23_, r_n_312__22_, r_n_312__21_, r_n_312__20_, r_n_312__19_, r_n_312__18_, r_n_312__17_, r_n_312__16_, r_n_312__15_, r_n_312__14_, r_n_312__13_, r_n_312__12_, r_n_312__11_, r_n_312__10_, r_n_312__9_, r_n_312__8_, r_n_312__7_, r_n_312__6_, r_n_312__5_, r_n_312__4_, r_n_312__3_, r_n_312__2_, r_n_312__1_, r_n_312__0_ } = (N624)? { r_313__63_, r_313__62_, r_313__61_, r_313__60_, r_313__59_, r_313__58_, r_313__57_, r_313__56_, r_313__55_, r_313__54_, r_313__53_, r_313__52_, r_313__51_, r_313__50_, r_313__49_, r_313__48_, r_313__47_, r_313__46_, r_313__45_, r_313__44_, r_313__43_, r_313__42_, r_313__41_, r_313__40_, r_313__39_, r_313__38_, r_313__37_, r_313__36_, r_313__35_, r_313__34_, r_313__33_, r_313__32_, r_313__31_, r_313__30_, r_313__29_, r_313__28_, r_313__27_, r_313__26_, r_313__25_, r_313__24_, r_313__23_, r_313__22_, r_313__21_, r_313__20_, r_313__19_, r_313__18_, r_313__17_, r_313__16_, r_313__15_, r_313__14_, r_313__13_, r_313__12_, r_313__11_, r_313__10_, r_313__9_, r_313__8_, r_313__7_, r_313__6_, r_313__5_, r_313__4_, r_313__3_, r_313__2_, r_313__1_, r_313__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N625)? data_i : 1'b0;
  assign N624 = sel_i[624];
  assign N625 = N2588;
  assign { r_n_313__63_, r_n_313__62_, r_n_313__61_, r_n_313__60_, r_n_313__59_, r_n_313__58_, r_n_313__57_, r_n_313__56_, r_n_313__55_, r_n_313__54_, r_n_313__53_, r_n_313__52_, r_n_313__51_, r_n_313__50_, r_n_313__49_, r_n_313__48_, r_n_313__47_, r_n_313__46_, r_n_313__45_, r_n_313__44_, r_n_313__43_, r_n_313__42_, r_n_313__41_, r_n_313__40_, r_n_313__39_, r_n_313__38_, r_n_313__37_, r_n_313__36_, r_n_313__35_, r_n_313__34_, r_n_313__33_, r_n_313__32_, r_n_313__31_, r_n_313__30_, r_n_313__29_, r_n_313__28_, r_n_313__27_, r_n_313__26_, r_n_313__25_, r_n_313__24_, r_n_313__23_, r_n_313__22_, r_n_313__21_, r_n_313__20_, r_n_313__19_, r_n_313__18_, r_n_313__17_, r_n_313__16_, r_n_313__15_, r_n_313__14_, r_n_313__13_, r_n_313__12_, r_n_313__11_, r_n_313__10_, r_n_313__9_, r_n_313__8_, r_n_313__7_, r_n_313__6_, r_n_313__5_, r_n_313__4_, r_n_313__3_, r_n_313__2_, r_n_313__1_, r_n_313__0_ } = (N626)? { r_314__63_, r_314__62_, r_314__61_, r_314__60_, r_314__59_, r_314__58_, r_314__57_, r_314__56_, r_314__55_, r_314__54_, r_314__53_, r_314__52_, r_314__51_, r_314__50_, r_314__49_, r_314__48_, r_314__47_, r_314__46_, r_314__45_, r_314__44_, r_314__43_, r_314__42_, r_314__41_, r_314__40_, r_314__39_, r_314__38_, r_314__37_, r_314__36_, r_314__35_, r_314__34_, r_314__33_, r_314__32_, r_314__31_, r_314__30_, r_314__29_, r_314__28_, r_314__27_, r_314__26_, r_314__25_, r_314__24_, r_314__23_, r_314__22_, r_314__21_, r_314__20_, r_314__19_, r_314__18_, r_314__17_, r_314__16_, r_314__15_, r_314__14_, r_314__13_, r_314__12_, r_314__11_, r_314__10_, r_314__9_, r_314__8_, r_314__7_, r_314__6_, r_314__5_, r_314__4_, r_314__3_, r_314__2_, r_314__1_, r_314__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N627)? data_i : 1'b0;
  assign N626 = sel_i[626];
  assign N627 = N2593;
  assign { r_n_314__63_, r_n_314__62_, r_n_314__61_, r_n_314__60_, r_n_314__59_, r_n_314__58_, r_n_314__57_, r_n_314__56_, r_n_314__55_, r_n_314__54_, r_n_314__53_, r_n_314__52_, r_n_314__51_, r_n_314__50_, r_n_314__49_, r_n_314__48_, r_n_314__47_, r_n_314__46_, r_n_314__45_, r_n_314__44_, r_n_314__43_, r_n_314__42_, r_n_314__41_, r_n_314__40_, r_n_314__39_, r_n_314__38_, r_n_314__37_, r_n_314__36_, r_n_314__35_, r_n_314__34_, r_n_314__33_, r_n_314__32_, r_n_314__31_, r_n_314__30_, r_n_314__29_, r_n_314__28_, r_n_314__27_, r_n_314__26_, r_n_314__25_, r_n_314__24_, r_n_314__23_, r_n_314__22_, r_n_314__21_, r_n_314__20_, r_n_314__19_, r_n_314__18_, r_n_314__17_, r_n_314__16_, r_n_314__15_, r_n_314__14_, r_n_314__13_, r_n_314__12_, r_n_314__11_, r_n_314__10_, r_n_314__9_, r_n_314__8_, r_n_314__7_, r_n_314__6_, r_n_314__5_, r_n_314__4_, r_n_314__3_, r_n_314__2_, r_n_314__1_, r_n_314__0_ } = (N628)? { r_315__63_, r_315__62_, r_315__61_, r_315__60_, r_315__59_, r_315__58_, r_315__57_, r_315__56_, r_315__55_, r_315__54_, r_315__53_, r_315__52_, r_315__51_, r_315__50_, r_315__49_, r_315__48_, r_315__47_, r_315__46_, r_315__45_, r_315__44_, r_315__43_, r_315__42_, r_315__41_, r_315__40_, r_315__39_, r_315__38_, r_315__37_, r_315__36_, r_315__35_, r_315__34_, r_315__33_, r_315__32_, r_315__31_, r_315__30_, r_315__29_, r_315__28_, r_315__27_, r_315__26_, r_315__25_, r_315__24_, r_315__23_, r_315__22_, r_315__21_, r_315__20_, r_315__19_, r_315__18_, r_315__17_, r_315__16_, r_315__15_, r_315__14_, r_315__13_, r_315__12_, r_315__11_, r_315__10_, r_315__9_, r_315__8_, r_315__7_, r_315__6_, r_315__5_, r_315__4_, r_315__3_, r_315__2_, r_315__1_, r_315__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N629)? data_i : 1'b0;
  assign N628 = sel_i[628];
  assign N629 = N2598;
  assign { r_n_315__63_, r_n_315__62_, r_n_315__61_, r_n_315__60_, r_n_315__59_, r_n_315__58_, r_n_315__57_, r_n_315__56_, r_n_315__55_, r_n_315__54_, r_n_315__53_, r_n_315__52_, r_n_315__51_, r_n_315__50_, r_n_315__49_, r_n_315__48_, r_n_315__47_, r_n_315__46_, r_n_315__45_, r_n_315__44_, r_n_315__43_, r_n_315__42_, r_n_315__41_, r_n_315__40_, r_n_315__39_, r_n_315__38_, r_n_315__37_, r_n_315__36_, r_n_315__35_, r_n_315__34_, r_n_315__33_, r_n_315__32_, r_n_315__31_, r_n_315__30_, r_n_315__29_, r_n_315__28_, r_n_315__27_, r_n_315__26_, r_n_315__25_, r_n_315__24_, r_n_315__23_, r_n_315__22_, r_n_315__21_, r_n_315__20_, r_n_315__19_, r_n_315__18_, r_n_315__17_, r_n_315__16_, r_n_315__15_, r_n_315__14_, r_n_315__13_, r_n_315__12_, r_n_315__11_, r_n_315__10_, r_n_315__9_, r_n_315__8_, r_n_315__7_, r_n_315__6_, r_n_315__5_, r_n_315__4_, r_n_315__3_, r_n_315__2_, r_n_315__1_, r_n_315__0_ } = (N630)? { r_316__63_, r_316__62_, r_316__61_, r_316__60_, r_316__59_, r_316__58_, r_316__57_, r_316__56_, r_316__55_, r_316__54_, r_316__53_, r_316__52_, r_316__51_, r_316__50_, r_316__49_, r_316__48_, r_316__47_, r_316__46_, r_316__45_, r_316__44_, r_316__43_, r_316__42_, r_316__41_, r_316__40_, r_316__39_, r_316__38_, r_316__37_, r_316__36_, r_316__35_, r_316__34_, r_316__33_, r_316__32_, r_316__31_, r_316__30_, r_316__29_, r_316__28_, r_316__27_, r_316__26_, r_316__25_, r_316__24_, r_316__23_, r_316__22_, r_316__21_, r_316__20_, r_316__19_, r_316__18_, r_316__17_, r_316__16_, r_316__15_, r_316__14_, r_316__13_, r_316__12_, r_316__11_, r_316__10_, r_316__9_, r_316__8_, r_316__7_, r_316__6_, r_316__5_, r_316__4_, r_316__3_, r_316__2_, r_316__1_, r_316__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N631)? data_i : 1'b0;
  assign N630 = sel_i[630];
  assign N631 = N2603;
  assign { r_n_316__63_, r_n_316__62_, r_n_316__61_, r_n_316__60_, r_n_316__59_, r_n_316__58_, r_n_316__57_, r_n_316__56_, r_n_316__55_, r_n_316__54_, r_n_316__53_, r_n_316__52_, r_n_316__51_, r_n_316__50_, r_n_316__49_, r_n_316__48_, r_n_316__47_, r_n_316__46_, r_n_316__45_, r_n_316__44_, r_n_316__43_, r_n_316__42_, r_n_316__41_, r_n_316__40_, r_n_316__39_, r_n_316__38_, r_n_316__37_, r_n_316__36_, r_n_316__35_, r_n_316__34_, r_n_316__33_, r_n_316__32_, r_n_316__31_, r_n_316__30_, r_n_316__29_, r_n_316__28_, r_n_316__27_, r_n_316__26_, r_n_316__25_, r_n_316__24_, r_n_316__23_, r_n_316__22_, r_n_316__21_, r_n_316__20_, r_n_316__19_, r_n_316__18_, r_n_316__17_, r_n_316__16_, r_n_316__15_, r_n_316__14_, r_n_316__13_, r_n_316__12_, r_n_316__11_, r_n_316__10_, r_n_316__9_, r_n_316__8_, r_n_316__7_, r_n_316__6_, r_n_316__5_, r_n_316__4_, r_n_316__3_, r_n_316__2_, r_n_316__1_, r_n_316__0_ } = (N632)? { r_317__63_, r_317__62_, r_317__61_, r_317__60_, r_317__59_, r_317__58_, r_317__57_, r_317__56_, r_317__55_, r_317__54_, r_317__53_, r_317__52_, r_317__51_, r_317__50_, r_317__49_, r_317__48_, r_317__47_, r_317__46_, r_317__45_, r_317__44_, r_317__43_, r_317__42_, r_317__41_, r_317__40_, r_317__39_, r_317__38_, r_317__37_, r_317__36_, r_317__35_, r_317__34_, r_317__33_, r_317__32_, r_317__31_, r_317__30_, r_317__29_, r_317__28_, r_317__27_, r_317__26_, r_317__25_, r_317__24_, r_317__23_, r_317__22_, r_317__21_, r_317__20_, r_317__19_, r_317__18_, r_317__17_, r_317__16_, r_317__15_, r_317__14_, r_317__13_, r_317__12_, r_317__11_, r_317__10_, r_317__9_, r_317__8_, r_317__7_, r_317__6_, r_317__5_, r_317__4_, r_317__3_, r_317__2_, r_317__1_, r_317__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N633)? data_i : 1'b0;
  assign N632 = sel_i[632];
  assign N633 = N2608;
  assign { r_n_317__63_, r_n_317__62_, r_n_317__61_, r_n_317__60_, r_n_317__59_, r_n_317__58_, r_n_317__57_, r_n_317__56_, r_n_317__55_, r_n_317__54_, r_n_317__53_, r_n_317__52_, r_n_317__51_, r_n_317__50_, r_n_317__49_, r_n_317__48_, r_n_317__47_, r_n_317__46_, r_n_317__45_, r_n_317__44_, r_n_317__43_, r_n_317__42_, r_n_317__41_, r_n_317__40_, r_n_317__39_, r_n_317__38_, r_n_317__37_, r_n_317__36_, r_n_317__35_, r_n_317__34_, r_n_317__33_, r_n_317__32_, r_n_317__31_, r_n_317__30_, r_n_317__29_, r_n_317__28_, r_n_317__27_, r_n_317__26_, r_n_317__25_, r_n_317__24_, r_n_317__23_, r_n_317__22_, r_n_317__21_, r_n_317__20_, r_n_317__19_, r_n_317__18_, r_n_317__17_, r_n_317__16_, r_n_317__15_, r_n_317__14_, r_n_317__13_, r_n_317__12_, r_n_317__11_, r_n_317__10_, r_n_317__9_, r_n_317__8_, r_n_317__7_, r_n_317__6_, r_n_317__5_, r_n_317__4_, r_n_317__3_, r_n_317__2_, r_n_317__1_, r_n_317__0_ } = (N634)? { r_318__63_, r_318__62_, r_318__61_, r_318__60_, r_318__59_, r_318__58_, r_318__57_, r_318__56_, r_318__55_, r_318__54_, r_318__53_, r_318__52_, r_318__51_, r_318__50_, r_318__49_, r_318__48_, r_318__47_, r_318__46_, r_318__45_, r_318__44_, r_318__43_, r_318__42_, r_318__41_, r_318__40_, r_318__39_, r_318__38_, r_318__37_, r_318__36_, r_318__35_, r_318__34_, r_318__33_, r_318__32_, r_318__31_, r_318__30_, r_318__29_, r_318__28_, r_318__27_, r_318__26_, r_318__25_, r_318__24_, r_318__23_, r_318__22_, r_318__21_, r_318__20_, r_318__19_, r_318__18_, r_318__17_, r_318__16_, r_318__15_, r_318__14_, r_318__13_, r_318__12_, r_318__11_, r_318__10_, r_318__9_, r_318__8_, r_318__7_, r_318__6_, r_318__5_, r_318__4_, r_318__3_, r_318__2_, r_318__1_, r_318__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N635)? data_i : 1'b0;
  assign N634 = sel_i[634];
  assign N635 = N2613;
  assign { r_n_318__63_, r_n_318__62_, r_n_318__61_, r_n_318__60_, r_n_318__59_, r_n_318__58_, r_n_318__57_, r_n_318__56_, r_n_318__55_, r_n_318__54_, r_n_318__53_, r_n_318__52_, r_n_318__51_, r_n_318__50_, r_n_318__49_, r_n_318__48_, r_n_318__47_, r_n_318__46_, r_n_318__45_, r_n_318__44_, r_n_318__43_, r_n_318__42_, r_n_318__41_, r_n_318__40_, r_n_318__39_, r_n_318__38_, r_n_318__37_, r_n_318__36_, r_n_318__35_, r_n_318__34_, r_n_318__33_, r_n_318__32_, r_n_318__31_, r_n_318__30_, r_n_318__29_, r_n_318__28_, r_n_318__27_, r_n_318__26_, r_n_318__25_, r_n_318__24_, r_n_318__23_, r_n_318__22_, r_n_318__21_, r_n_318__20_, r_n_318__19_, r_n_318__18_, r_n_318__17_, r_n_318__16_, r_n_318__15_, r_n_318__14_, r_n_318__13_, r_n_318__12_, r_n_318__11_, r_n_318__10_, r_n_318__9_, r_n_318__8_, r_n_318__7_, r_n_318__6_, r_n_318__5_, r_n_318__4_, r_n_318__3_, r_n_318__2_, r_n_318__1_, r_n_318__0_ } = (N636)? { r_319__63_, r_319__62_, r_319__61_, r_319__60_, r_319__59_, r_319__58_, r_319__57_, r_319__56_, r_319__55_, r_319__54_, r_319__53_, r_319__52_, r_319__51_, r_319__50_, r_319__49_, r_319__48_, r_319__47_, r_319__46_, r_319__45_, r_319__44_, r_319__43_, r_319__42_, r_319__41_, r_319__40_, r_319__39_, r_319__38_, r_319__37_, r_319__36_, r_319__35_, r_319__34_, r_319__33_, r_319__32_, r_319__31_, r_319__30_, r_319__29_, r_319__28_, r_319__27_, r_319__26_, r_319__25_, r_319__24_, r_319__23_, r_319__22_, r_319__21_, r_319__20_, r_319__19_, r_319__18_, r_319__17_, r_319__16_, r_319__15_, r_319__14_, r_319__13_, r_319__12_, r_319__11_, r_319__10_, r_319__9_, r_319__8_, r_319__7_, r_319__6_, r_319__5_, r_319__4_, r_319__3_, r_319__2_, r_319__1_, r_319__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N637)? data_i : 1'b0;
  assign N636 = sel_i[636];
  assign N637 = N2618;
  assign { r_n_319__63_, r_n_319__62_, r_n_319__61_, r_n_319__60_, r_n_319__59_, r_n_319__58_, r_n_319__57_, r_n_319__56_, r_n_319__55_, r_n_319__54_, r_n_319__53_, r_n_319__52_, r_n_319__51_, r_n_319__50_, r_n_319__49_, r_n_319__48_, r_n_319__47_, r_n_319__46_, r_n_319__45_, r_n_319__44_, r_n_319__43_, r_n_319__42_, r_n_319__41_, r_n_319__40_, r_n_319__39_, r_n_319__38_, r_n_319__37_, r_n_319__36_, r_n_319__35_, r_n_319__34_, r_n_319__33_, r_n_319__32_, r_n_319__31_, r_n_319__30_, r_n_319__29_, r_n_319__28_, r_n_319__27_, r_n_319__26_, r_n_319__25_, r_n_319__24_, r_n_319__23_, r_n_319__22_, r_n_319__21_, r_n_319__20_, r_n_319__19_, r_n_319__18_, r_n_319__17_, r_n_319__16_, r_n_319__15_, r_n_319__14_, r_n_319__13_, r_n_319__12_, r_n_319__11_, r_n_319__10_, r_n_319__9_, r_n_319__8_, r_n_319__7_, r_n_319__6_, r_n_319__5_, r_n_319__4_, r_n_319__3_, r_n_319__2_, r_n_319__1_, r_n_319__0_ } = (N638)? { r_320__63_, r_320__62_, r_320__61_, r_320__60_, r_320__59_, r_320__58_, r_320__57_, r_320__56_, r_320__55_, r_320__54_, r_320__53_, r_320__52_, r_320__51_, r_320__50_, r_320__49_, r_320__48_, r_320__47_, r_320__46_, r_320__45_, r_320__44_, r_320__43_, r_320__42_, r_320__41_, r_320__40_, r_320__39_, r_320__38_, r_320__37_, r_320__36_, r_320__35_, r_320__34_, r_320__33_, r_320__32_, r_320__31_, r_320__30_, r_320__29_, r_320__28_, r_320__27_, r_320__26_, r_320__25_, r_320__24_, r_320__23_, r_320__22_, r_320__21_, r_320__20_, r_320__19_, r_320__18_, r_320__17_, r_320__16_, r_320__15_, r_320__14_, r_320__13_, r_320__12_, r_320__11_, r_320__10_, r_320__9_, r_320__8_, r_320__7_, r_320__6_, r_320__5_, r_320__4_, r_320__3_, r_320__2_, r_320__1_, r_320__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N639)? data_i : 1'b0;
  assign N638 = sel_i[638];
  assign N639 = N2623;
  assign { r_n_320__63_, r_n_320__62_, r_n_320__61_, r_n_320__60_, r_n_320__59_, r_n_320__58_, r_n_320__57_, r_n_320__56_, r_n_320__55_, r_n_320__54_, r_n_320__53_, r_n_320__52_, r_n_320__51_, r_n_320__50_, r_n_320__49_, r_n_320__48_, r_n_320__47_, r_n_320__46_, r_n_320__45_, r_n_320__44_, r_n_320__43_, r_n_320__42_, r_n_320__41_, r_n_320__40_, r_n_320__39_, r_n_320__38_, r_n_320__37_, r_n_320__36_, r_n_320__35_, r_n_320__34_, r_n_320__33_, r_n_320__32_, r_n_320__31_, r_n_320__30_, r_n_320__29_, r_n_320__28_, r_n_320__27_, r_n_320__26_, r_n_320__25_, r_n_320__24_, r_n_320__23_, r_n_320__22_, r_n_320__21_, r_n_320__20_, r_n_320__19_, r_n_320__18_, r_n_320__17_, r_n_320__16_, r_n_320__15_, r_n_320__14_, r_n_320__13_, r_n_320__12_, r_n_320__11_, r_n_320__10_, r_n_320__9_, r_n_320__8_, r_n_320__7_, r_n_320__6_, r_n_320__5_, r_n_320__4_, r_n_320__3_, r_n_320__2_, r_n_320__1_, r_n_320__0_ } = (N640)? { r_321__63_, r_321__62_, r_321__61_, r_321__60_, r_321__59_, r_321__58_, r_321__57_, r_321__56_, r_321__55_, r_321__54_, r_321__53_, r_321__52_, r_321__51_, r_321__50_, r_321__49_, r_321__48_, r_321__47_, r_321__46_, r_321__45_, r_321__44_, r_321__43_, r_321__42_, r_321__41_, r_321__40_, r_321__39_, r_321__38_, r_321__37_, r_321__36_, r_321__35_, r_321__34_, r_321__33_, r_321__32_, r_321__31_, r_321__30_, r_321__29_, r_321__28_, r_321__27_, r_321__26_, r_321__25_, r_321__24_, r_321__23_, r_321__22_, r_321__21_, r_321__20_, r_321__19_, r_321__18_, r_321__17_, r_321__16_, r_321__15_, r_321__14_, r_321__13_, r_321__12_, r_321__11_, r_321__10_, r_321__9_, r_321__8_, r_321__7_, r_321__6_, r_321__5_, r_321__4_, r_321__3_, r_321__2_, r_321__1_, r_321__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N641)? data_i : 1'b0;
  assign N640 = sel_i[640];
  assign N641 = N2628;
  assign { r_n_321__63_, r_n_321__62_, r_n_321__61_, r_n_321__60_, r_n_321__59_, r_n_321__58_, r_n_321__57_, r_n_321__56_, r_n_321__55_, r_n_321__54_, r_n_321__53_, r_n_321__52_, r_n_321__51_, r_n_321__50_, r_n_321__49_, r_n_321__48_, r_n_321__47_, r_n_321__46_, r_n_321__45_, r_n_321__44_, r_n_321__43_, r_n_321__42_, r_n_321__41_, r_n_321__40_, r_n_321__39_, r_n_321__38_, r_n_321__37_, r_n_321__36_, r_n_321__35_, r_n_321__34_, r_n_321__33_, r_n_321__32_, r_n_321__31_, r_n_321__30_, r_n_321__29_, r_n_321__28_, r_n_321__27_, r_n_321__26_, r_n_321__25_, r_n_321__24_, r_n_321__23_, r_n_321__22_, r_n_321__21_, r_n_321__20_, r_n_321__19_, r_n_321__18_, r_n_321__17_, r_n_321__16_, r_n_321__15_, r_n_321__14_, r_n_321__13_, r_n_321__12_, r_n_321__11_, r_n_321__10_, r_n_321__9_, r_n_321__8_, r_n_321__7_, r_n_321__6_, r_n_321__5_, r_n_321__4_, r_n_321__3_, r_n_321__2_, r_n_321__1_, r_n_321__0_ } = (N642)? { r_322__63_, r_322__62_, r_322__61_, r_322__60_, r_322__59_, r_322__58_, r_322__57_, r_322__56_, r_322__55_, r_322__54_, r_322__53_, r_322__52_, r_322__51_, r_322__50_, r_322__49_, r_322__48_, r_322__47_, r_322__46_, r_322__45_, r_322__44_, r_322__43_, r_322__42_, r_322__41_, r_322__40_, r_322__39_, r_322__38_, r_322__37_, r_322__36_, r_322__35_, r_322__34_, r_322__33_, r_322__32_, r_322__31_, r_322__30_, r_322__29_, r_322__28_, r_322__27_, r_322__26_, r_322__25_, r_322__24_, r_322__23_, r_322__22_, r_322__21_, r_322__20_, r_322__19_, r_322__18_, r_322__17_, r_322__16_, r_322__15_, r_322__14_, r_322__13_, r_322__12_, r_322__11_, r_322__10_, r_322__9_, r_322__8_, r_322__7_, r_322__6_, r_322__5_, r_322__4_, r_322__3_, r_322__2_, r_322__1_, r_322__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N643)? data_i : 1'b0;
  assign N642 = sel_i[642];
  assign N643 = N2633;
  assign { r_n_322__63_, r_n_322__62_, r_n_322__61_, r_n_322__60_, r_n_322__59_, r_n_322__58_, r_n_322__57_, r_n_322__56_, r_n_322__55_, r_n_322__54_, r_n_322__53_, r_n_322__52_, r_n_322__51_, r_n_322__50_, r_n_322__49_, r_n_322__48_, r_n_322__47_, r_n_322__46_, r_n_322__45_, r_n_322__44_, r_n_322__43_, r_n_322__42_, r_n_322__41_, r_n_322__40_, r_n_322__39_, r_n_322__38_, r_n_322__37_, r_n_322__36_, r_n_322__35_, r_n_322__34_, r_n_322__33_, r_n_322__32_, r_n_322__31_, r_n_322__30_, r_n_322__29_, r_n_322__28_, r_n_322__27_, r_n_322__26_, r_n_322__25_, r_n_322__24_, r_n_322__23_, r_n_322__22_, r_n_322__21_, r_n_322__20_, r_n_322__19_, r_n_322__18_, r_n_322__17_, r_n_322__16_, r_n_322__15_, r_n_322__14_, r_n_322__13_, r_n_322__12_, r_n_322__11_, r_n_322__10_, r_n_322__9_, r_n_322__8_, r_n_322__7_, r_n_322__6_, r_n_322__5_, r_n_322__4_, r_n_322__3_, r_n_322__2_, r_n_322__1_, r_n_322__0_ } = (N644)? { r_323__63_, r_323__62_, r_323__61_, r_323__60_, r_323__59_, r_323__58_, r_323__57_, r_323__56_, r_323__55_, r_323__54_, r_323__53_, r_323__52_, r_323__51_, r_323__50_, r_323__49_, r_323__48_, r_323__47_, r_323__46_, r_323__45_, r_323__44_, r_323__43_, r_323__42_, r_323__41_, r_323__40_, r_323__39_, r_323__38_, r_323__37_, r_323__36_, r_323__35_, r_323__34_, r_323__33_, r_323__32_, r_323__31_, r_323__30_, r_323__29_, r_323__28_, r_323__27_, r_323__26_, r_323__25_, r_323__24_, r_323__23_, r_323__22_, r_323__21_, r_323__20_, r_323__19_, r_323__18_, r_323__17_, r_323__16_, r_323__15_, r_323__14_, r_323__13_, r_323__12_, r_323__11_, r_323__10_, r_323__9_, r_323__8_, r_323__7_, r_323__6_, r_323__5_, r_323__4_, r_323__3_, r_323__2_, r_323__1_, r_323__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N645)? data_i : 1'b0;
  assign N644 = sel_i[644];
  assign N645 = N2638;
  assign { r_n_323__63_, r_n_323__62_, r_n_323__61_, r_n_323__60_, r_n_323__59_, r_n_323__58_, r_n_323__57_, r_n_323__56_, r_n_323__55_, r_n_323__54_, r_n_323__53_, r_n_323__52_, r_n_323__51_, r_n_323__50_, r_n_323__49_, r_n_323__48_, r_n_323__47_, r_n_323__46_, r_n_323__45_, r_n_323__44_, r_n_323__43_, r_n_323__42_, r_n_323__41_, r_n_323__40_, r_n_323__39_, r_n_323__38_, r_n_323__37_, r_n_323__36_, r_n_323__35_, r_n_323__34_, r_n_323__33_, r_n_323__32_, r_n_323__31_, r_n_323__30_, r_n_323__29_, r_n_323__28_, r_n_323__27_, r_n_323__26_, r_n_323__25_, r_n_323__24_, r_n_323__23_, r_n_323__22_, r_n_323__21_, r_n_323__20_, r_n_323__19_, r_n_323__18_, r_n_323__17_, r_n_323__16_, r_n_323__15_, r_n_323__14_, r_n_323__13_, r_n_323__12_, r_n_323__11_, r_n_323__10_, r_n_323__9_, r_n_323__8_, r_n_323__7_, r_n_323__6_, r_n_323__5_, r_n_323__4_, r_n_323__3_, r_n_323__2_, r_n_323__1_, r_n_323__0_ } = (N646)? { r_324__63_, r_324__62_, r_324__61_, r_324__60_, r_324__59_, r_324__58_, r_324__57_, r_324__56_, r_324__55_, r_324__54_, r_324__53_, r_324__52_, r_324__51_, r_324__50_, r_324__49_, r_324__48_, r_324__47_, r_324__46_, r_324__45_, r_324__44_, r_324__43_, r_324__42_, r_324__41_, r_324__40_, r_324__39_, r_324__38_, r_324__37_, r_324__36_, r_324__35_, r_324__34_, r_324__33_, r_324__32_, r_324__31_, r_324__30_, r_324__29_, r_324__28_, r_324__27_, r_324__26_, r_324__25_, r_324__24_, r_324__23_, r_324__22_, r_324__21_, r_324__20_, r_324__19_, r_324__18_, r_324__17_, r_324__16_, r_324__15_, r_324__14_, r_324__13_, r_324__12_, r_324__11_, r_324__10_, r_324__9_, r_324__8_, r_324__7_, r_324__6_, r_324__5_, r_324__4_, r_324__3_, r_324__2_, r_324__1_, r_324__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N647)? data_i : 1'b0;
  assign N646 = sel_i[646];
  assign N647 = N2643;
  assign { r_n_324__63_, r_n_324__62_, r_n_324__61_, r_n_324__60_, r_n_324__59_, r_n_324__58_, r_n_324__57_, r_n_324__56_, r_n_324__55_, r_n_324__54_, r_n_324__53_, r_n_324__52_, r_n_324__51_, r_n_324__50_, r_n_324__49_, r_n_324__48_, r_n_324__47_, r_n_324__46_, r_n_324__45_, r_n_324__44_, r_n_324__43_, r_n_324__42_, r_n_324__41_, r_n_324__40_, r_n_324__39_, r_n_324__38_, r_n_324__37_, r_n_324__36_, r_n_324__35_, r_n_324__34_, r_n_324__33_, r_n_324__32_, r_n_324__31_, r_n_324__30_, r_n_324__29_, r_n_324__28_, r_n_324__27_, r_n_324__26_, r_n_324__25_, r_n_324__24_, r_n_324__23_, r_n_324__22_, r_n_324__21_, r_n_324__20_, r_n_324__19_, r_n_324__18_, r_n_324__17_, r_n_324__16_, r_n_324__15_, r_n_324__14_, r_n_324__13_, r_n_324__12_, r_n_324__11_, r_n_324__10_, r_n_324__9_, r_n_324__8_, r_n_324__7_, r_n_324__6_, r_n_324__5_, r_n_324__4_, r_n_324__3_, r_n_324__2_, r_n_324__1_, r_n_324__0_ } = (N648)? { r_325__63_, r_325__62_, r_325__61_, r_325__60_, r_325__59_, r_325__58_, r_325__57_, r_325__56_, r_325__55_, r_325__54_, r_325__53_, r_325__52_, r_325__51_, r_325__50_, r_325__49_, r_325__48_, r_325__47_, r_325__46_, r_325__45_, r_325__44_, r_325__43_, r_325__42_, r_325__41_, r_325__40_, r_325__39_, r_325__38_, r_325__37_, r_325__36_, r_325__35_, r_325__34_, r_325__33_, r_325__32_, r_325__31_, r_325__30_, r_325__29_, r_325__28_, r_325__27_, r_325__26_, r_325__25_, r_325__24_, r_325__23_, r_325__22_, r_325__21_, r_325__20_, r_325__19_, r_325__18_, r_325__17_, r_325__16_, r_325__15_, r_325__14_, r_325__13_, r_325__12_, r_325__11_, r_325__10_, r_325__9_, r_325__8_, r_325__7_, r_325__6_, r_325__5_, r_325__4_, r_325__3_, r_325__2_, r_325__1_, r_325__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N649)? data_i : 1'b0;
  assign N648 = sel_i[648];
  assign N649 = N2648;
  assign { r_n_325__63_, r_n_325__62_, r_n_325__61_, r_n_325__60_, r_n_325__59_, r_n_325__58_, r_n_325__57_, r_n_325__56_, r_n_325__55_, r_n_325__54_, r_n_325__53_, r_n_325__52_, r_n_325__51_, r_n_325__50_, r_n_325__49_, r_n_325__48_, r_n_325__47_, r_n_325__46_, r_n_325__45_, r_n_325__44_, r_n_325__43_, r_n_325__42_, r_n_325__41_, r_n_325__40_, r_n_325__39_, r_n_325__38_, r_n_325__37_, r_n_325__36_, r_n_325__35_, r_n_325__34_, r_n_325__33_, r_n_325__32_, r_n_325__31_, r_n_325__30_, r_n_325__29_, r_n_325__28_, r_n_325__27_, r_n_325__26_, r_n_325__25_, r_n_325__24_, r_n_325__23_, r_n_325__22_, r_n_325__21_, r_n_325__20_, r_n_325__19_, r_n_325__18_, r_n_325__17_, r_n_325__16_, r_n_325__15_, r_n_325__14_, r_n_325__13_, r_n_325__12_, r_n_325__11_, r_n_325__10_, r_n_325__9_, r_n_325__8_, r_n_325__7_, r_n_325__6_, r_n_325__5_, r_n_325__4_, r_n_325__3_, r_n_325__2_, r_n_325__1_, r_n_325__0_ } = (N650)? { r_326__63_, r_326__62_, r_326__61_, r_326__60_, r_326__59_, r_326__58_, r_326__57_, r_326__56_, r_326__55_, r_326__54_, r_326__53_, r_326__52_, r_326__51_, r_326__50_, r_326__49_, r_326__48_, r_326__47_, r_326__46_, r_326__45_, r_326__44_, r_326__43_, r_326__42_, r_326__41_, r_326__40_, r_326__39_, r_326__38_, r_326__37_, r_326__36_, r_326__35_, r_326__34_, r_326__33_, r_326__32_, r_326__31_, r_326__30_, r_326__29_, r_326__28_, r_326__27_, r_326__26_, r_326__25_, r_326__24_, r_326__23_, r_326__22_, r_326__21_, r_326__20_, r_326__19_, r_326__18_, r_326__17_, r_326__16_, r_326__15_, r_326__14_, r_326__13_, r_326__12_, r_326__11_, r_326__10_, r_326__9_, r_326__8_, r_326__7_, r_326__6_, r_326__5_, r_326__4_, r_326__3_, r_326__2_, r_326__1_, r_326__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N651)? data_i : 1'b0;
  assign N650 = sel_i[650];
  assign N651 = N2653;
  assign { r_n_326__63_, r_n_326__62_, r_n_326__61_, r_n_326__60_, r_n_326__59_, r_n_326__58_, r_n_326__57_, r_n_326__56_, r_n_326__55_, r_n_326__54_, r_n_326__53_, r_n_326__52_, r_n_326__51_, r_n_326__50_, r_n_326__49_, r_n_326__48_, r_n_326__47_, r_n_326__46_, r_n_326__45_, r_n_326__44_, r_n_326__43_, r_n_326__42_, r_n_326__41_, r_n_326__40_, r_n_326__39_, r_n_326__38_, r_n_326__37_, r_n_326__36_, r_n_326__35_, r_n_326__34_, r_n_326__33_, r_n_326__32_, r_n_326__31_, r_n_326__30_, r_n_326__29_, r_n_326__28_, r_n_326__27_, r_n_326__26_, r_n_326__25_, r_n_326__24_, r_n_326__23_, r_n_326__22_, r_n_326__21_, r_n_326__20_, r_n_326__19_, r_n_326__18_, r_n_326__17_, r_n_326__16_, r_n_326__15_, r_n_326__14_, r_n_326__13_, r_n_326__12_, r_n_326__11_, r_n_326__10_, r_n_326__9_, r_n_326__8_, r_n_326__7_, r_n_326__6_, r_n_326__5_, r_n_326__4_, r_n_326__3_, r_n_326__2_, r_n_326__1_, r_n_326__0_ } = (N652)? { r_327__63_, r_327__62_, r_327__61_, r_327__60_, r_327__59_, r_327__58_, r_327__57_, r_327__56_, r_327__55_, r_327__54_, r_327__53_, r_327__52_, r_327__51_, r_327__50_, r_327__49_, r_327__48_, r_327__47_, r_327__46_, r_327__45_, r_327__44_, r_327__43_, r_327__42_, r_327__41_, r_327__40_, r_327__39_, r_327__38_, r_327__37_, r_327__36_, r_327__35_, r_327__34_, r_327__33_, r_327__32_, r_327__31_, r_327__30_, r_327__29_, r_327__28_, r_327__27_, r_327__26_, r_327__25_, r_327__24_, r_327__23_, r_327__22_, r_327__21_, r_327__20_, r_327__19_, r_327__18_, r_327__17_, r_327__16_, r_327__15_, r_327__14_, r_327__13_, r_327__12_, r_327__11_, r_327__10_, r_327__9_, r_327__8_, r_327__7_, r_327__6_, r_327__5_, r_327__4_, r_327__3_, r_327__2_, r_327__1_, r_327__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N653)? data_i : 1'b0;
  assign N652 = sel_i[652];
  assign N653 = N2658;
  assign { r_n_327__63_, r_n_327__62_, r_n_327__61_, r_n_327__60_, r_n_327__59_, r_n_327__58_, r_n_327__57_, r_n_327__56_, r_n_327__55_, r_n_327__54_, r_n_327__53_, r_n_327__52_, r_n_327__51_, r_n_327__50_, r_n_327__49_, r_n_327__48_, r_n_327__47_, r_n_327__46_, r_n_327__45_, r_n_327__44_, r_n_327__43_, r_n_327__42_, r_n_327__41_, r_n_327__40_, r_n_327__39_, r_n_327__38_, r_n_327__37_, r_n_327__36_, r_n_327__35_, r_n_327__34_, r_n_327__33_, r_n_327__32_, r_n_327__31_, r_n_327__30_, r_n_327__29_, r_n_327__28_, r_n_327__27_, r_n_327__26_, r_n_327__25_, r_n_327__24_, r_n_327__23_, r_n_327__22_, r_n_327__21_, r_n_327__20_, r_n_327__19_, r_n_327__18_, r_n_327__17_, r_n_327__16_, r_n_327__15_, r_n_327__14_, r_n_327__13_, r_n_327__12_, r_n_327__11_, r_n_327__10_, r_n_327__9_, r_n_327__8_, r_n_327__7_, r_n_327__6_, r_n_327__5_, r_n_327__4_, r_n_327__3_, r_n_327__2_, r_n_327__1_, r_n_327__0_ } = (N654)? { r_328__63_, r_328__62_, r_328__61_, r_328__60_, r_328__59_, r_328__58_, r_328__57_, r_328__56_, r_328__55_, r_328__54_, r_328__53_, r_328__52_, r_328__51_, r_328__50_, r_328__49_, r_328__48_, r_328__47_, r_328__46_, r_328__45_, r_328__44_, r_328__43_, r_328__42_, r_328__41_, r_328__40_, r_328__39_, r_328__38_, r_328__37_, r_328__36_, r_328__35_, r_328__34_, r_328__33_, r_328__32_, r_328__31_, r_328__30_, r_328__29_, r_328__28_, r_328__27_, r_328__26_, r_328__25_, r_328__24_, r_328__23_, r_328__22_, r_328__21_, r_328__20_, r_328__19_, r_328__18_, r_328__17_, r_328__16_, r_328__15_, r_328__14_, r_328__13_, r_328__12_, r_328__11_, r_328__10_, r_328__9_, r_328__8_, r_328__7_, r_328__6_, r_328__5_, r_328__4_, r_328__3_, r_328__2_, r_328__1_, r_328__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N655)? data_i : 1'b0;
  assign N654 = sel_i[654];
  assign N655 = N2663;
  assign { r_n_328__63_, r_n_328__62_, r_n_328__61_, r_n_328__60_, r_n_328__59_, r_n_328__58_, r_n_328__57_, r_n_328__56_, r_n_328__55_, r_n_328__54_, r_n_328__53_, r_n_328__52_, r_n_328__51_, r_n_328__50_, r_n_328__49_, r_n_328__48_, r_n_328__47_, r_n_328__46_, r_n_328__45_, r_n_328__44_, r_n_328__43_, r_n_328__42_, r_n_328__41_, r_n_328__40_, r_n_328__39_, r_n_328__38_, r_n_328__37_, r_n_328__36_, r_n_328__35_, r_n_328__34_, r_n_328__33_, r_n_328__32_, r_n_328__31_, r_n_328__30_, r_n_328__29_, r_n_328__28_, r_n_328__27_, r_n_328__26_, r_n_328__25_, r_n_328__24_, r_n_328__23_, r_n_328__22_, r_n_328__21_, r_n_328__20_, r_n_328__19_, r_n_328__18_, r_n_328__17_, r_n_328__16_, r_n_328__15_, r_n_328__14_, r_n_328__13_, r_n_328__12_, r_n_328__11_, r_n_328__10_, r_n_328__9_, r_n_328__8_, r_n_328__7_, r_n_328__6_, r_n_328__5_, r_n_328__4_, r_n_328__3_, r_n_328__2_, r_n_328__1_, r_n_328__0_ } = (N656)? { r_329__63_, r_329__62_, r_329__61_, r_329__60_, r_329__59_, r_329__58_, r_329__57_, r_329__56_, r_329__55_, r_329__54_, r_329__53_, r_329__52_, r_329__51_, r_329__50_, r_329__49_, r_329__48_, r_329__47_, r_329__46_, r_329__45_, r_329__44_, r_329__43_, r_329__42_, r_329__41_, r_329__40_, r_329__39_, r_329__38_, r_329__37_, r_329__36_, r_329__35_, r_329__34_, r_329__33_, r_329__32_, r_329__31_, r_329__30_, r_329__29_, r_329__28_, r_329__27_, r_329__26_, r_329__25_, r_329__24_, r_329__23_, r_329__22_, r_329__21_, r_329__20_, r_329__19_, r_329__18_, r_329__17_, r_329__16_, r_329__15_, r_329__14_, r_329__13_, r_329__12_, r_329__11_, r_329__10_, r_329__9_, r_329__8_, r_329__7_, r_329__6_, r_329__5_, r_329__4_, r_329__3_, r_329__2_, r_329__1_, r_329__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N657)? data_i : 1'b0;
  assign N656 = sel_i[656];
  assign N657 = N2668;
  assign { r_n_329__63_, r_n_329__62_, r_n_329__61_, r_n_329__60_, r_n_329__59_, r_n_329__58_, r_n_329__57_, r_n_329__56_, r_n_329__55_, r_n_329__54_, r_n_329__53_, r_n_329__52_, r_n_329__51_, r_n_329__50_, r_n_329__49_, r_n_329__48_, r_n_329__47_, r_n_329__46_, r_n_329__45_, r_n_329__44_, r_n_329__43_, r_n_329__42_, r_n_329__41_, r_n_329__40_, r_n_329__39_, r_n_329__38_, r_n_329__37_, r_n_329__36_, r_n_329__35_, r_n_329__34_, r_n_329__33_, r_n_329__32_, r_n_329__31_, r_n_329__30_, r_n_329__29_, r_n_329__28_, r_n_329__27_, r_n_329__26_, r_n_329__25_, r_n_329__24_, r_n_329__23_, r_n_329__22_, r_n_329__21_, r_n_329__20_, r_n_329__19_, r_n_329__18_, r_n_329__17_, r_n_329__16_, r_n_329__15_, r_n_329__14_, r_n_329__13_, r_n_329__12_, r_n_329__11_, r_n_329__10_, r_n_329__9_, r_n_329__8_, r_n_329__7_, r_n_329__6_, r_n_329__5_, r_n_329__4_, r_n_329__3_, r_n_329__2_, r_n_329__1_, r_n_329__0_ } = (N658)? { r_330__63_, r_330__62_, r_330__61_, r_330__60_, r_330__59_, r_330__58_, r_330__57_, r_330__56_, r_330__55_, r_330__54_, r_330__53_, r_330__52_, r_330__51_, r_330__50_, r_330__49_, r_330__48_, r_330__47_, r_330__46_, r_330__45_, r_330__44_, r_330__43_, r_330__42_, r_330__41_, r_330__40_, r_330__39_, r_330__38_, r_330__37_, r_330__36_, r_330__35_, r_330__34_, r_330__33_, r_330__32_, r_330__31_, r_330__30_, r_330__29_, r_330__28_, r_330__27_, r_330__26_, r_330__25_, r_330__24_, r_330__23_, r_330__22_, r_330__21_, r_330__20_, r_330__19_, r_330__18_, r_330__17_, r_330__16_, r_330__15_, r_330__14_, r_330__13_, r_330__12_, r_330__11_, r_330__10_, r_330__9_, r_330__8_, r_330__7_, r_330__6_, r_330__5_, r_330__4_, r_330__3_, r_330__2_, r_330__1_, r_330__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N659)? data_i : 1'b0;
  assign N658 = sel_i[658];
  assign N659 = N2673;
  assign { r_n_330__63_, r_n_330__62_, r_n_330__61_, r_n_330__60_, r_n_330__59_, r_n_330__58_, r_n_330__57_, r_n_330__56_, r_n_330__55_, r_n_330__54_, r_n_330__53_, r_n_330__52_, r_n_330__51_, r_n_330__50_, r_n_330__49_, r_n_330__48_, r_n_330__47_, r_n_330__46_, r_n_330__45_, r_n_330__44_, r_n_330__43_, r_n_330__42_, r_n_330__41_, r_n_330__40_, r_n_330__39_, r_n_330__38_, r_n_330__37_, r_n_330__36_, r_n_330__35_, r_n_330__34_, r_n_330__33_, r_n_330__32_, r_n_330__31_, r_n_330__30_, r_n_330__29_, r_n_330__28_, r_n_330__27_, r_n_330__26_, r_n_330__25_, r_n_330__24_, r_n_330__23_, r_n_330__22_, r_n_330__21_, r_n_330__20_, r_n_330__19_, r_n_330__18_, r_n_330__17_, r_n_330__16_, r_n_330__15_, r_n_330__14_, r_n_330__13_, r_n_330__12_, r_n_330__11_, r_n_330__10_, r_n_330__9_, r_n_330__8_, r_n_330__7_, r_n_330__6_, r_n_330__5_, r_n_330__4_, r_n_330__3_, r_n_330__2_, r_n_330__1_, r_n_330__0_ } = (N660)? { r_331__63_, r_331__62_, r_331__61_, r_331__60_, r_331__59_, r_331__58_, r_331__57_, r_331__56_, r_331__55_, r_331__54_, r_331__53_, r_331__52_, r_331__51_, r_331__50_, r_331__49_, r_331__48_, r_331__47_, r_331__46_, r_331__45_, r_331__44_, r_331__43_, r_331__42_, r_331__41_, r_331__40_, r_331__39_, r_331__38_, r_331__37_, r_331__36_, r_331__35_, r_331__34_, r_331__33_, r_331__32_, r_331__31_, r_331__30_, r_331__29_, r_331__28_, r_331__27_, r_331__26_, r_331__25_, r_331__24_, r_331__23_, r_331__22_, r_331__21_, r_331__20_, r_331__19_, r_331__18_, r_331__17_, r_331__16_, r_331__15_, r_331__14_, r_331__13_, r_331__12_, r_331__11_, r_331__10_, r_331__9_, r_331__8_, r_331__7_, r_331__6_, r_331__5_, r_331__4_, r_331__3_, r_331__2_, r_331__1_, r_331__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N661)? data_i : 1'b0;
  assign N660 = sel_i[660];
  assign N661 = N2678;
  assign { r_n_331__63_, r_n_331__62_, r_n_331__61_, r_n_331__60_, r_n_331__59_, r_n_331__58_, r_n_331__57_, r_n_331__56_, r_n_331__55_, r_n_331__54_, r_n_331__53_, r_n_331__52_, r_n_331__51_, r_n_331__50_, r_n_331__49_, r_n_331__48_, r_n_331__47_, r_n_331__46_, r_n_331__45_, r_n_331__44_, r_n_331__43_, r_n_331__42_, r_n_331__41_, r_n_331__40_, r_n_331__39_, r_n_331__38_, r_n_331__37_, r_n_331__36_, r_n_331__35_, r_n_331__34_, r_n_331__33_, r_n_331__32_, r_n_331__31_, r_n_331__30_, r_n_331__29_, r_n_331__28_, r_n_331__27_, r_n_331__26_, r_n_331__25_, r_n_331__24_, r_n_331__23_, r_n_331__22_, r_n_331__21_, r_n_331__20_, r_n_331__19_, r_n_331__18_, r_n_331__17_, r_n_331__16_, r_n_331__15_, r_n_331__14_, r_n_331__13_, r_n_331__12_, r_n_331__11_, r_n_331__10_, r_n_331__9_, r_n_331__8_, r_n_331__7_, r_n_331__6_, r_n_331__5_, r_n_331__4_, r_n_331__3_, r_n_331__2_, r_n_331__1_, r_n_331__0_ } = (N662)? { r_332__63_, r_332__62_, r_332__61_, r_332__60_, r_332__59_, r_332__58_, r_332__57_, r_332__56_, r_332__55_, r_332__54_, r_332__53_, r_332__52_, r_332__51_, r_332__50_, r_332__49_, r_332__48_, r_332__47_, r_332__46_, r_332__45_, r_332__44_, r_332__43_, r_332__42_, r_332__41_, r_332__40_, r_332__39_, r_332__38_, r_332__37_, r_332__36_, r_332__35_, r_332__34_, r_332__33_, r_332__32_, r_332__31_, r_332__30_, r_332__29_, r_332__28_, r_332__27_, r_332__26_, r_332__25_, r_332__24_, r_332__23_, r_332__22_, r_332__21_, r_332__20_, r_332__19_, r_332__18_, r_332__17_, r_332__16_, r_332__15_, r_332__14_, r_332__13_, r_332__12_, r_332__11_, r_332__10_, r_332__9_, r_332__8_, r_332__7_, r_332__6_, r_332__5_, r_332__4_, r_332__3_, r_332__2_, r_332__1_, r_332__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N663)? data_i : 1'b0;
  assign N662 = sel_i[662];
  assign N663 = N2683;
  assign { r_n_332__63_, r_n_332__62_, r_n_332__61_, r_n_332__60_, r_n_332__59_, r_n_332__58_, r_n_332__57_, r_n_332__56_, r_n_332__55_, r_n_332__54_, r_n_332__53_, r_n_332__52_, r_n_332__51_, r_n_332__50_, r_n_332__49_, r_n_332__48_, r_n_332__47_, r_n_332__46_, r_n_332__45_, r_n_332__44_, r_n_332__43_, r_n_332__42_, r_n_332__41_, r_n_332__40_, r_n_332__39_, r_n_332__38_, r_n_332__37_, r_n_332__36_, r_n_332__35_, r_n_332__34_, r_n_332__33_, r_n_332__32_, r_n_332__31_, r_n_332__30_, r_n_332__29_, r_n_332__28_, r_n_332__27_, r_n_332__26_, r_n_332__25_, r_n_332__24_, r_n_332__23_, r_n_332__22_, r_n_332__21_, r_n_332__20_, r_n_332__19_, r_n_332__18_, r_n_332__17_, r_n_332__16_, r_n_332__15_, r_n_332__14_, r_n_332__13_, r_n_332__12_, r_n_332__11_, r_n_332__10_, r_n_332__9_, r_n_332__8_, r_n_332__7_, r_n_332__6_, r_n_332__5_, r_n_332__4_, r_n_332__3_, r_n_332__2_, r_n_332__1_, r_n_332__0_ } = (N664)? { r_333__63_, r_333__62_, r_333__61_, r_333__60_, r_333__59_, r_333__58_, r_333__57_, r_333__56_, r_333__55_, r_333__54_, r_333__53_, r_333__52_, r_333__51_, r_333__50_, r_333__49_, r_333__48_, r_333__47_, r_333__46_, r_333__45_, r_333__44_, r_333__43_, r_333__42_, r_333__41_, r_333__40_, r_333__39_, r_333__38_, r_333__37_, r_333__36_, r_333__35_, r_333__34_, r_333__33_, r_333__32_, r_333__31_, r_333__30_, r_333__29_, r_333__28_, r_333__27_, r_333__26_, r_333__25_, r_333__24_, r_333__23_, r_333__22_, r_333__21_, r_333__20_, r_333__19_, r_333__18_, r_333__17_, r_333__16_, r_333__15_, r_333__14_, r_333__13_, r_333__12_, r_333__11_, r_333__10_, r_333__9_, r_333__8_, r_333__7_, r_333__6_, r_333__5_, r_333__4_, r_333__3_, r_333__2_, r_333__1_, r_333__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N665)? data_i : 1'b0;
  assign N664 = sel_i[664];
  assign N665 = N2688;
  assign { r_n_333__63_, r_n_333__62_, r_n_333__61_, r_n_333__60_, r_n_333__59_, r_n_333__58_, r_n_333__57_, r_n_333__56_, r_n_333__55_, r_n_333__54_, r_n_333__53_, r_n_333__52_, r_n_333__51_, r_n_333__50_, r_n_333__49_, r_n_333__48_, r_n_333__47_, r_n_333__46_, r_n_333__45_, r_n_333__44_, r_n_333__43_, r_n_333__42_, r_n_333__41_, r_n_333__40_, r_n_333__39_, r_n_333__38_, r_n_333__37_, r_n_333__36_, r_n_333__35_, r_n_333__34_, r_n_333__33_, r_n_333__32_, r_n_333__31_, r_n_333__30_, r_n_333__29_, r_n_333__28_, r_n_333__27_, r_n_333__26_, r_n_333__25_, r_n_333__24_, r_n_333__23_, r_n_333__22_, r_n_333__21_, r_n_333__20_, r_n_333__19_, r_n_333__18_, r_n_333__17_, r_n_333__16_, r_n_333__15_, r_n_333__14_, r_n_333__13_, r_n_333__12_, r_n_333__11_, r_n_333__10_, r_n_333__9_, r_n_333__8_, r_n_333__7_, r_n_333__6_, r_n_333__5_, r_n_333__4_, r_n_333__3_, r_n_333__2_, r_n_333__1_, r_n_333__0_ } = (N666)? { r_334__63_, r_334__62_, r_334__61_, r_334__60_, r_334__59_, r_334__58_, r_334__57_, r_334__56_, r_334__55_, r_334__54_, r_334__53_, r_334__52_, r_334__51_, r_334__50_, r_334__49_, r_334__48_, r_334__47_, r_334__46_, r_334__45_, r_334__44_, r_334__43_, r_334__42_, r_334__41_, r_334__40_, r_334__39_, r_334__38_, r_334__37_, r_334__36_, r_334__35_, r_334__34_, r_334__33_, r_334__32_, r_334__31_, r_334__30_, r_334__29_, r_334__28_, r_334__27_, r_334__26_, r_334__25_, r_334__24_, r_334__23_, r_334__22_, r_334__21_, r_334__20_, r_334__19_, r_334__18_, r_334__17_, r_334__16_, r_334__15_, r_334__14_, r_334__13_, r_334__12_, r_334__11_, r_334__10_, r_334__9_, r_334__8_, r_334__7_, r_334__6_, r_334__5_, r_334__4_, r_334__3_, r_334__2_, r_334__1_, r_334__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N667)? data_i : 1'b0;
  assign N666 = sel_i[666];
  assign N667 = N2693;
  assign { r_n_334__63_, r_n_334__62_, r_n_334__61_, r_n_334__60_, r_n_334__59_, r_n_334__58_, r_n_334__57_, r_n_334__56_, r_n_334__55_, r_n_334__54_, r_n_334__53_, r_n_334__52_, r_n_334__51_, r_n_334__50_, r_n_334__49_, r_n_334__48_, r_n_334__47_, r_n_334__46_, r_n_334__45_, r_n_334__44_, r_n_334__43_, r_n_334__42_, r_n_334__41_, r_n_334__40_, r_n_334__39_, r_n_334__38_, r_n_334__37_, r_n_334__36_, r_n_334__35_, r_n_334__34_, r_n_334__33_, r_n_334__32_, r_n_334__31_, r_n_334__30_, r_n_334__29_, r_n_334__28_, r_n_334__27_, r_n_334__26_, r_n_334__25_, r_n_334__24_, r_n_334__23_, r_n_334__22_, r_n_334__21_, r_n_334__20_, r_n_334__19_, r_n_334__18_, r_n_334__17_, r_n_334__16_, r_n_334__15_, r_n_334__14_, r_n_334__13_, r_n_334__12_, r_n_334__11_, r_n_334__10_, r_n_334__9_, r_n_334__8_, r_n_334__7_, r_n_334__6_, r_n_334__5_, r_n_334__4_, r_n_334__3_, r_n_334__2_, r_n_334__1_, r_n_334__0_ } = (N668)? { r_335__63_, r_335__62_, r_335__61_, r_335__60_, r_335__59_, r_335__58_, r_335__57_, r_335__56_, r_335__55_, r_335__54_, r_335__53_, r_335__52_, r_335__51_, r_335__50_, r_335__49_, r_335__48_, r_335__47_, r_335__46_, r_335__45_, r_335__44_, r_335__43_, r_335__42_, r_335__41_, r_335__40_, r_335__39_, r_335__38_, r_335__37_, r_335__36_, r_335__35_, r_335__34_, r_335__33_, r_335__32_, r_335__31_, r_335__30_, r_335__29_, r_335__28_, r_335__27_, r_335__26_, r_335__25_, r_335__24_, r_335__23_, r_335__22_, r_335__21_, r_335__20_, r_335__19_, r_335__18_, r_335__17_, r_335__16_, r_335__15_, r_335__14_, r_335__13_, r_335__12_, r_335__11_, r_335__10_, r_335__9_, r_335__8_, r_335__7_, r_335__6_, r_335__5_, r_335__4_, r_335__3_, r_335__2_, r_335__1_, r_335__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N669)? data_i : 1'b0;
  assign N668 = sel_i[668];
  assign N669 = N2698;
  assign { r_n_335__63_, r_n_335__62_, r_n_335__61_, r_n_335__60_, r_n_335__59_, r_n_335__58_, r_n_335__57_, r_n_335__56_, r_n_335__55_, r_n_335__54_, r_n_335__53_, r_n_335__52_, r_n_335__51_, r_n_335__50_, r_n_335__49_, r_n_335__48_, r_n_335__47_, r_n_335__46_, r_n_335__45_, r_n_335__44_, r_n_335__43_, r_n_335__42_, r_n_335__41_, r_n_335__40_, r_n_335__39_, r_n_335__38_, r_n_335__37_, r_n_335__36_, r_n_335__35_, r_n_335__34_, r_n_335__33_, r_n_335__32_, r_n_335__31_, r_n_335__30_, r_n_335__29_, r_n_335__28_, r_n_335__27_, r_n_335__26_, r_n_335__25_, r_n_335__24_, r_n_335__23_, r_n_335__22_, r_n_335__21_, r_n_335__20_, r_n_335__19_, r_n_335__18_, r_n_335__17_, r_n_335__16_, r_n_335__15_, r_n_335__14_, r_n_335__13_, r_n_335__12_, r_n_335__11_, r_n_335__10_, r_n_335__9_, r_n_335__8_, r_n_335__7_, r_n_335__6_, r_n_335__5_, r_n_335__4_, r_n_335__3_, r_n_335__2_, r_n_335__1_, r_n_335__0_ } = (N670)? { r_336__63_, r_336__62_, r_336__61_, r_336__60_, r_336__59_, r_336__58_, r_336__57_, r_336__56_, r_336__55_, r_336__54_, r_336__53_, r_336__52_, r_336__51_, r_336__50_, r_336__49_, r_336__48_, r_336__47_, r_336__46_, r_336__45_, r_336__44_, r_336__43_, r_336__42_, r_336__41_, r_336__40_, r_336__39_, r_336__38_, r_336__37_, r_336__36_, r_336__35_, r_336__34_, r_336__33_, r_336__32_, r_336__31_, r_336__30_, r_336__29_, r_336__28_, r_336__27_, r_336__26_, r_336__25_, r_336__24_, r_336__23_, r_336__22_, r_336__21_, r_336__20_, r_336__19_, r_336__18_, r_336__17_, r_336__16_, r_336__15_, r_336__14_, r_336__13_, r_336__12_, r_336__11_, r_336__10_, r_336__9_, r_336__8_, r_336__7_, r_336__6_, r_336__5_, r_336__4_, r_336__3_, r_336__2_, r_336__1_, r_336__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N671)? data_i : 1'b0;
  assign N670 = sel_i[670];
  assign N671 = N2703;
  assign { r_n_336__63_, r_n_336__62_, r_n_336__61_, r_n_336__60_, r_n_336__59_, r_n_336__58_, r_n_336__57_, r_n_336__56_, r_n_336__55_, r_n_336__54_, r_n_336__53_, r_n_336__52_, r_n_336__51_, r_n_336__50_, r_n_336__49_, r_n_336__48_, r_n_336__47_, r_n_336__46_, r_n_336__45_, r_n_336__44_, r_n_336__43_, r_n_336__42_, r_n_336__41_, r_n_336__40_, r_n_336__39_, r_n_336__38_, r_n_336__37_, r_n_336__36_, r_n_336__35_, r_n_336__34_, r_n_336__33_, r_n_336__32_, r_n_336__31_, r_n_336__30_, r_n_336__29_, r_n_336__28_, r_n_336__27_, r_n_336__26_, r_n_336__25_, r_n_336__24_, r_n_336__23_, r_n_336__22_, r_n_336__21_, r_n_336__20_, r_n_336__19_, r_n_336__18_, r_n_336__17_, r_n_336__16_, r_n_336__15_, r_n_336__14_, r_n_336__13_, r_n_336__12_, r_n_336__11_, r_n_336__10_, r_n_336__9_, r_n_336__8_, r_n_336__7_, r_n_336__6_, r_n_336__5_, r_n_336__4_, r_n_336__3_, r_n_336__2_, r_n_336__1_, r_n_336__0_ } = (N672)? { r_337__63_, r_337__62_, r_337__61_, r_337__60_, r_337__59_, r_337__58_, r_337__57_, r_337__56_, r_337__55_, r_337__54_, r_337__53_, r_337__52_, r_337__51_, r_337__50_, r_337__49_, r_337__48_, r_337__47_, r_337__46_, r_337__45_, r_337__44_, r_337__43_, r_337__42_, r_337__41_, r_337__40_, r_337__39_, r_337__38_, r_337__37_, r_337__36_, r_337__35_, r_337__34_, r_337__33_, r_337__32_, r_337__31_, r_337__30_, r_337__29_, r_337__28_, r_337__27_, r_337__26_, r_337__25_, r_337__24_, r_337__23_, r_337__22_, r_337__21_, r_337__20_, r_337__19_, r_337__18_, r_337__17_, r_337__16_, r_337__15_, r_337__14_, r_337__13_, r_337__12_, r_337__11_, r_337__10_, r_337__9_, r_337__8_, r_337__7_, r_337__6_, r_337__5_, r_337__4_, r_337__3_, r_337__2_, r_337__1_, r_337__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N673)? data_i : 1'b0;
  assign N672 = sel_i[672];
  assign N673 = N2708;
  assign { r_n_337__63_, r_n_337__62_, r_n_337__61_, r_n_337__60_, r_n_337__59_, r_n_337__58_, r_n_337__57_, r_n_337__56_, r_n_337__55_, r_n_337__54_, r_n_337__53_, r_n_337__52_, r_n_337__51_, r_n_337__50_, r_n_337__49_, r_n_337__48_, r_n_337__47_, r_n_337__46_, r_n_337__45_, r_n_337__44_, r_n_337__43_, r_n_337__42_, r_n_337__41_, r_n_337__40_, r_n_337__39_, r_n_337__38_, r_n_337__37_, r_n_337__36_, r_n_337__35_, r_n_337__34_, r_n_337__33_, r_n_337__32_, r_n_337__31_, r_n_337__30_, r_n_337__29_, r_n_337__28_, r_n_337__27_, r_n_337__26_, r_n_337__25_, r_n_337__24_, r_n_337__23_, r_n_337__22_, r_n_337__21_, r_n_337__20_, r_n_337__19_, r_n_337__18_, r_n_337__17_, r_n_337__16_, r_n_337__15_, r_n_337__14_, r_n_337__13_, r_n_337__12_, r_n_337__11_, r_n_337__10_, r_n_337__9_, r_n_337__8_, r_n_337__7_, r_n_337__6_, r_n_337__5_, r_n_337__4_, r_n_337__3_, r_n_337__2_, r_n_337__1_, r_n_337__0_ } = (N674)? { r_338__63_, r_338__62_, r_338__61_, r_338__60_, r_338__59_, r_338__58_, r_338__57_, r_338__56_, r_338__55_, r_338__54_, r_338__53_, r_338__52_, r_338__51_, r_338__50_, r_338__49_, r_338__48_, r_338__47_, r_338__46_, r_338__45_, r_338__44_, r_338__43_, r_338__42_, r_338__41_, r_338__40_, r_338__39_, r_338__38_, r_338__37_, r_338__36_, r_338__35_, r_338__34_, r_338__33_, r_338__32_, r_338__31_, r_338__30_, r_338__29_, r_338__28_, r_338__27_, r_338__26_, r_338__25_, r_338__24_, r_338__23_, r_338__22_, r_338__21_, r_338__20_, r_338__19_, r_338__18_, r_338__17_, r_338__16_, r_338__15_, r_338__14_, r_338__13_, r_338__12_, r_338__11_, r_338__10_, r_338__9_, r_338__8_, r_338__7_, r_338__6_, r_338__5_, r_338__4_, r_338__3_, r_338__2_, r_338__1_, r_338__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N675)? data_i : 1'b0;
  assign N674 = sel_i[674];
  assign N675 = N2713;
  assign { r_n_338__63_, r_n_338__62_, r_n_338__61_, r_n_338__60_, r_n_338__59_, r_n_338__58_, r_n_338__57_, r_n_338__56_, r_n_338__55_, r_n_338__54_, r_n_338__53_, r_n_338__52_, r_n_338__51_, r_n_338__50_, r_n_338__49_, r_n_338__48_, r_n_338__47_, r_n_338__46_, r_n_338__45_, r_n_338__44_, r_n_338__43_, r_n_338__42_, r_n_338__41_, r_n_338__40_, r_n_338__39_, r_n_338__38_, r_n_338__37_, r_n_338__36_, r_n_338__35_, r_n_338__34_, r_n_338__33_, r_n_338__32_, r_n_338__31_, r_n_338__30_, r_n_338__29_, r_n_338__28_, r_n_338__27_, r_n_338__26_, r_n_338__25_, r_n_338__24_, r_n_338__23_, r_n_338__22_, r_n_338__21_, r_n_338__20_, r_n_338__19_, r_n_338__18_, r_n_338__17_, r_n_338__16_, r_n_338__15_, r_n_338__14_, r_n_338__13_, r_n_338__12_, r_n_338__11_, r_n_338__10_, r_n_338__9_, r_n_338__8_, r_n_338__7_, r_n_338__6_, r_n_338__5_, r_n_338__4_, r_n_338__3_, r_n_338__2_, r_n_338__1_, r_n_338__0_ } = (N676)? { r_339__63_, r_339__62_, r_339__61_, r_339__60_, r_339__59_, r_339__58_, r_339__57_, r_339__56_, r_339__55_, r_339__54_, r_339__53_, r_339__52_, r_339__51_, r_339__50_, r_339__49_, r_339__48_, r_339__47_, r_339__46_, r_339__45_, r_339__44_, r_339__43_, r_339__42_, r_339__41_, r_339__40_, r_339__39_, r_339__38_, r_339__37_, r_339__36_, r_339__35_, r_339__34_, r_339__33_, r_339__32_, r_339__31_, r_339__30_, r_339__29_, r_339__28_, r_339__27_, r_339__26_, r_339__25_, r_339__24_, r_339__23_, r_339__22_, r_339__21_, r_339__20_, r_339__19_, r_339__18_, r_339__17_, r_339__16_, r_339__15_, r_339__14_, r_339__13_, r_339__12_, r_339__11_, r_339__10_, r_339__9_, r_339__8_, r_339__7_, r_339__6_, r_339__5_, r_339__4_, r_339__3_, r_339__2_, r_339__1_, r_339__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N677)? data_i : 1'b0;
  assign N676 = sel_i[676];
  assign N677 = N2718;
  assign { r_n_339__63_, r_n_339__62_, r_n_339__61_, r_n_339__60_, r_n_339__59_, r_n_339__58_, r_n_339__57_, r_n_339__56_, r_n_339__55_, r_n_339__54_, r_n_339__53_, r_n_339__52_, r_n_339__51_, r_n_339__50_, r_n_339__49_, r_n_339__48_, r_n_339__47_, r_n_339__46_, r_n_339__45_, r_n_339__44_, r_n_339__43_, r_n_339__42_, r_n_339__41_, r_n_339__40_, r_n_339__39_, r_n_339__38_, r_n_339__37_, r_n_339__36_, r_n_339__35_, r_n_339__34_, r_n_339__33_, r_n_339__32_, r_n_339__31_, r_n_339__30_, r_n_339__29_, r_n_339__28_, r_n_339__27_, r_n_339__26_, r_n_339__25_, r_n_339__24_, r_n_339__23_, r_n_339__22_, r_n_339__21_, r_n_339__20_, r_n_339__19_, r_n_339__18_, r_n_339__17_, r_n_339__16_, r_n_339__15_, r_n_339__14_, r_n_339__13_, r_n_339__12_, r_n_339__11_, r_n_339__10_, r_n_339__9_, r_n_339__8_, r_n_339__7_, r_n_339__6_, r_n_339__5_, r_n_339__4_, r_n_339__3_, r_n_339__2_, r_n_339__1_, r_n_339__0_ } = (N678)? { r_340__63_, r_340__62_, r_340__61_, r_340__60_, r_340__59_, r_340__58_, r_340__57_, r_340__56_, r_340__55_, r_340__54_, r_340__53_, r_340__52_, r_340__51_, r_340__50_, r_340__49_, r_340__48_, r_340__47_, r_340__46_, r_340__45_, r_340__44_, r_340__43_, r_340__42_, r_340__41_, r_340__40_, r_340__39_, r_340__38_, r_340__37_, r_340__36_, r_340__35_, r_340__34_, r_340__33_, r_340__32_, r_340__31_, r_340__30_, r_340__29_, r_340__28_, r_340__27_, r_340__26_, r_340__25_, r_340__24_, r_340__23_, r_340__22_, r_340__21_, r_340__20_, r_340__19_, r_340__18_, r_340__17_, r_340__16_, r_340__15_, r_340__14_, r_340__13_, r_340__12_, r_340__11_, r_340__10_, r_340__9_, r_340__8_, r_340__7_, r_340__6_, r_340__5_, r_340__4_, r_340__3_, r_340__2_, r_340__1_, r_340__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N679)? data_i : 1'b0;
  assign N678 = sel_i[678];
  assign N679 = N2723;
  assign { r_n_340__63_, r_n_340__62_, r_n_340__61_, r_n_340__60_, r_n_340__59_, r_n_340__58_, r_n_340__57_, r_n_340__56_, r_n_340__55_, r_n_340__54_, r_n_340__53_, r_n_340__52_, r_n_340__51_, r_n_340__50_, r_n_340__49_, r_n_340__48_, r_n_340__47_, r_n_340__46_, r_n_340__45_, r_n_340__44_, r_n_340__43_, r_n_340__42_, r_n_340__41_, r_n_340__40_, r_n_340__39_, r_n_340__38_, r_n_340__37_, r_n_340__36_, r_n_340__35_, r_n_340__34_, r_n_340__33_, r_n_340__32_, r_n_340__31_, r_n_340__30_, r_n_340__29_, r_n_340__28_, r_n_340__27_, r_n_340__26_, r_n_340__25_, r_n_340__24_, r_n_340__23_, r_n_340__22_, r_n_340__21_, r_n_340__20_, r_n_340__19_, r_n_340__18_, r_n_340__17_, r_n_340__16_, r_n_340__15_, r_n_340__14_, r_n_340__13_, r_n_340__12_, r_n_340__11_, r_n_340__10_, r_n_340__9_, r_n_340__8_, r_n_340__7_, r_n_340__6_, r_n_340__5_, r_n_340__4_, r_n_340__3_, r_n_340__2_, r_n_340__1_, r_n_340__0_ } = (N680)? { r_341__63_, r_341__62_, r_341__61_, r_341__60_, r_341__59_, r_341__58_, r_341__57_, r_341__56_, r_341__55_, r_341__54_, r_341__53_, r_341__52_, r_341__51_, r_341__50_, r_341__49_, r_341__48_, r_341__47_, r_341__46_, r_341__45_, r_341__44_, r_341__43_, r_341__42_, r_341__41_, r_341__40_, r_341__39_, r_341__38_, r_341__37_, r_341__36_, r_341__35_, r_341__34_, r_341__33_, r_341__32_, r_341__31_, r_341__30_, r_341__29_, r_341__28_, r_341__27_, r_341__26_, r_341__25_, r_341__24_, r_341__23_, r_341__22_, r_341__21_, r_341__20_, r_341__19_, r_341__18_, r_341__17_, r_341__16_, r_341__15_, r_341__14_, r_341__13_, r_341__12_, r_341__11_, r_341__10_, r_341__9_, r_341__8_, r_341__7_, r_341__6_, r_341__5_, r_341__4_, r_341__3_, r_341__2_, r_341__1_, r_341__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N681)? data_i : 1'b0;
  assign N680 = sel_i[680];
  assign N681 = N2728;
  assign { r_n_341__63_, r_n_341__62_, r_n_341__61_, r_n_341__60_, r_n_341__59_, r_n_341__58_, r_n_341__57_, r_n_341__56_, r_n_341__55_, r_n_341__54_, r_n_341__53_, r_n_341__52_, r_n_341__51_, r_n_341__50_, r_n_341__49_, r_n_341__48_, r_n_341__47_, r_n_341__46_, r_n_341__45_, r_n_341__44_, r_n_341__43_, r_n_341__42_, r_n_341__41_, r_n_341__40_, r_n_341__39_, r_n_341__38_, r_n_341__37_, r_n_341__36_, r_n_341__35_, r_n_341__34_, r_n_341__33_, r_n_341__32_, r_n_341__31_, r_n_341__30_, r_n_341__29_, r_n_341__28_, r_n_341__27_, r_n_341__26_, r_n_341__25_, r_n_341__24_, r_n_341__23_, r_n_341__22_, r_n_341__21_, r_n_341__20_, r_n_341__19_, r_n_341__18_, r_n_341__17_, r_n_341__16_, r_n_341__15_, r_n_341__14_, r_n_341__13_, r_n_341__12_, r_n_341__11_, r_n_341__10_, r_n_341__9_, r_n_341__8_, r_n_341__7_, r_n_341__6_, r_n_341__5_, r_n_341__4_, r_n_341__3_, r_n_341__2_, r_n_341__1_, r_n_341__0_ } = (N682)? { r_342__63_, r_342__62_, r_342__61_, r_342__60_, r_342__59_, r_342__58_, r_342__57_, r_342__56_, r_342__55_, r_342__54_, r_342__53_, r_342__52_, r_342__51_, r_342__50_, r_342__49_, r_342__48_, r_342__47_, r_342__46_, r_342__45_, r_342__44_, r_342__43_, r_342__42_, r_342__41_, r_342__40_, r_342__39_, r_342__38_, r_342__37_, r_342__36_, r_342__35_, r_342__34_, r_342__33_, r_342__32_, r_342__31_, r_342__30_, r_342__29_, r_342__28_, r_342__27_, r_342__26_, r_342__25_, r_342__24_, r_342__23_, r_342__22_, r_342__21_, r_342__20_, r_342__19_, r_342__18_, r_342__17_, r_342__16_, r_342__15_, r_342__14_, r_342__13_, r_342__12_, r_342__11_, r_342__10_, r_342__9_, r_342__8_, r_342__7_, r_342__6_, r_342__5_, r_342__4_, r_342__3_, r_342__2_, r_342__1_, r_342__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N683)? data_i : 1'b0;
  assign N682 = sel_i[682];
  assign N683 = N2733;
  assign { r_n_342__63_, r_n_342__62_, r_n_342__61_, r_n_342__60_, r_n_342__59_, r_n_342__58_, r_n_342__57_, r_n_342__56_, r_n_342__55_, r_n_342__54_, r_n_342__53_, r_n_342__52_, r_n_342__51_, r_n_342__50_, r_n_342__49_, r_n_342__48_, r_n_342__47_, r_n_342__46_, r_n_342__45_, r_n_342__44_, r_n_342__43_, r_n_342__42_, r_n_342__41_, r_n_342__40_, r_n_342__39_, r_n_342__38_, r_n_342__37_, r_n_342__36_, r_n_342__35_, r_n_342__34_, r_n_342__33_, r_n_342__32_, r_n_342__31_, r_n_342__30_, r_n_342__29_, r_n_342__28_, r_n_342__27_, r_n_342__26_, r_n_342__25_, r_n_342__24_, r_n_342__23_, r_n_342__22_, r_n_342__21_, r_n_342__20_, r_n_342__19_, r_n_342__18_, r_n_342__17_, r_n_342__16_, r_n_342__15_, r_n_342__14_, r_n_342__13_, r_n_342__12_, r_n_342__11_, r_n_342__10_, r_n_342__9_, r_n_342__8_, r_n_342__7_, r_n_342__6_, r_n_342__5_, r_n_342__4_, r_n_342__3_, r_n_342__2_, r_n_342__1_, r_n_342__0_ } = (N684)? { r_343__63_, r_343__62_, r_343__61_, r_343__60_, r_343__59_, r_343__58_, r_343__57_, r_343__56_, r_343__55_, r_343__54_, r_343__53_, r_343__52_, r_343__51_, r_343__50_, r_343__49_, r_343__48_, r_343__47_, r_343__46_, r_343__45_, r_343__44_, r_343__43_, r_343__42_, r_343__41_, r_343__40_, r_343__39_, r_343__38_, r_343__37_, r_343__36_, r_343__35_, r_343__34_, r_343__33_, r_343__32_, r_343__31_, r_343__30_, r_343__29_, r_343__28_, r_343__27_, r_343__26_, r_343__25_, r_343__24_, r_343__23_, r_343__22_, r_343__21_, r_343__20_, r_343__19_, r_343__18_, r_343__17_, r_343__16_, r_343__15_, r_343__14_, r_343__13_, r_343__12_, r_343__11_, r_343__10_, r_343__9_, r_343__8_, r_343__7_, r_343__6_, r_343__5_, r_343__4_, r_343__3_, r_343__2_, r_343__1_, r_343__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N685)? data_i : 1'b0;
  assign N684 = sel_i[684];
  assign N685 = N2738;
  assign { r_n_343__63_, r_n_343__62_, r_n_343__61_, r_n_343__60_, r_n_343__59_, r_n_343__58_, r_n_343__57_, r_n_343__56_, r_n_343__55_, r_n_343__54_, r_n_343__53_, r_n_343__52_, r_n_343__51_, r_n_343__50_, r_n_343__49_, r_n_343__48_, r_n_343__47_, r_n_343__46_, r_n_343__45_, r_n_343__44_, r_n_343__43_, r_n_343__42_, r_n_343__41_, r_n_343__40_, r_n_343__39_, r_n_343__38_, r_n_343__37_, r_n_343__36_, r_n_343__35_, r_n_343__34_, r_n_343__33_, r_n_343__32_, r_n_343__31_, r_n_343__30_, r_n_343__29_, r_n_343__28_, r_n_343__27_, r_n_343__26_, r_n_343__25_, r_n_343__24_, r_n_343__23_, r_n_343__22_, r_n_343__21_, r_n_343__20_, r_n_343__19_, r_n_343__18_, r_n_343__17_, r_n_343__16_, r_n_343__15_, r_n_343__14_, r_n_343__13_, r_n_343__12_, r_n_343__11_, r_n_343__10_, r_n_343__9_, r_n_343__8_, r_n_343__7_, r_n_343__6_, r_n_343__5_, r_n_343__4_, r_n_343__3_, r_n_343__2_, r_n_343__1_, r_n_343__0_ } = (N686)? { r_344__63_, r_344__62_, r_344__61_, r_344__60_, r_344__59_, r_344__58_, r_344__57_, r_344__56_, r_344__55_, r_344__54_, r_344__53_, r_344__52_, r_344__51_, r_344__50_, r_344__49_, r_344__48_, r_344__47_, r_344__46_, r_344__45_, r_344__44_, r_344__43_, r_344__42_, r_344__41_, r_344__40_, r_344__39_, r_344__38_, r_344__37_, r_344__36_, r_344__35_, r_344__34_, r_344__33_, r_344__32_, r_344__31_, r_344__30_, r_344__29_, r_344__28_, r_344__27_, r_344__26_, r_344__25_, r_344__24_, r_344__23_, r_344__22_, r_344__21_, r_344__20_, r_344__19_, r_344__18_, r_344__17_, r_344__16_, r_344__15_, r_344__14_, r_344__13_, r_344__12_, r_344__11_, r_344__10_, r_344__9_, r_344__8_, r_344__7_, r_344__6_, r_344__5_, r_344__4_, r_344__3_, r_344__2_, r_344__1_, r_344__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N687)? data_i : 1'b0;
  assign N686 = sel_i[686];
  assign N687 = N2743;
  assign { r_n_344__63_, r_n_344__62_, r_n_344__61_, r_n_344__60_, r_n_344__59_, r_n_344__58_, r_n_344__57_, r_n_344__56_, r_n_344__55_, r_n_344__54_, r_n_344__53_, r_n_344__52_, r_n_344__51_, r_n_344__50_, r_n_344__49_, r_n_344__48_, r_n_344__47_, r_n_344__46_, r_n_344__45_, r_n_344__44_, r_n_344__43_, r_n_344__42_, r_n_344__41_, r_n_344__40_, r_n_344__39_, r_n_344__38_, r_n_344__37_, r_n_344__36_, r_n_344__35_, r_n_344__34_, r_n_344__33_, r_n_344__32_, r_n_344__31_, r_n_344__30_, r_n_344__29_, r_n_344__28_, r_n_344__27_, r_n_344__26_, r_n_344__25_, r_n_344__24_, r_n_344__23_, r_n_344__22_, r_n_344__21_, r_n_344__20_, r_n_344__19_, r_n_344__18_, r_n_344__17_, r_n_344__16_, r_n_344__15_, r_n_344__14_, r_n_344__13_, r_n_344__12_, r_n_344__11_, r_n_344__10_, r_n_344__9_, r_n_344__8_, r_n_344__7_, r_n_344__6_, r_n_344__5_, r_n_344__4_, r_n_344__3_, r_n_344__2_, r_n_344__1_, r_n_344__0_ } = (N688)? { r_345__63_, r_345__62_, r_345__61_, r_345__60_, r_345__59_, r_345__58_, r_345__57_, r_345__56_, r_345__55_, r_345__54_, r_345__53_, r_345__52_, r_345__51_, r_345__50_, r_345__49_, r_345__48_, r_345__47_, r_345__46_, r_345__45_, r_345__44_, r_345__43_, r_345__42_, r_345__41_, r_345__40_, r_345__39_, r_345__38_, r_345__37_, r_345__36_, r_345__35_, r_345__34_, r_345__33_, r_345__32_, r_345__31_, r_345__30_, r_345__29_, r_345__28_, r_345__27_, r_345__26_, r_345__25_, r_345__24_, r_345__23_, r_345__22_, r_345__21_, r_345__20_, r_345__19_, r_345__18_, r_345__17_, r_345__16_, r_345__15_, r_345__14_, r_345__13_, r_345__12_, r_345__11_, r_345__10_, r_345__9_, r_345__8_, r_345__7_, r_345__6_, r_345__5_, r_345__4_, r_345__3_, r_345__2_, r_345__1_, r_345__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N689)? data_i : 1'b0;
  assign N688 = sel_i[688];
  assign N689 = N2748;
  assign { r_n_345__63_, r_n_345__62_, r_n_345__61_, r_n_345__60_, r_n_345__59_, r_n_345__58_, r_n_345__57_, r_n_345__56_, r_n_345__55_, r_n_345__54_, r_n_345__53_, r_n_345__52_, r_n_345__51_, r_n_345__50_, r_n_345__49_, r_n_345__48_, r_n_345__47_, r_n_345__46_, r_n_345__45_, r_n_345__44_, r_n_345__43_, r_n_345__42_, r_n_345__41_, r_n_345__40_, r_n_345__39_, r_n_345__38_, r_n_345__37_, r_n_345__36_, r_n_345__35_, r_n_345__34_, r_n_345__33_, r_n_345__32_, r_n_345__31_, r_n_345__30_, r_n_345__29_, r_n_345__28_, r_n_345__27_, r_n_345__26_, r_n_345__25_, r_n_345__24_, r_n_345__23_, r_n_345__22_, r_n_345__21_, r_n_345__20_, r_n_345__19_, r_n_345__18_, r_n_345__17_, r_n_345__16_, r_n_345__15_, r_n_345__14_, r_n_345__13_, r_n_345__12_, r_n_345__11_, r_n_345__10_, r_n_345__9_, r_n_345__8_, r_n_345__7_, r_n_345__6_, r_n_345__5_, r_n_345__4_, r_n_345__3_, r_n_345__2_, r_n_345__1_, r_n_345__0_ } = (N690)? { r_346__63_, r_346__62_, r_346__61_, r_346__60_, r_346__59_, r_346__58_, r_346__57_, r_346__56_, r_346__55_, r_346__54_, r_346__53_, r_346__52_, r_346__51_, r_346__50_, r_346__49_, r_346__48_, r_346__47_, r_346__46_, r_346__45_, r_346__44_, r_346__43_, r_346__42_, r_346__41_, r_346__40_, r_346__39_, r_346__38_, r_346__37_, r_346__36_, r_346__35_, r_346__34_, r_346__33_, r_346__32_, r_346__31_, r_346__30_, r_346__29_, r_346__28_, r_346__27_, r_346__26_, r_346__25_, r_346__24_, r_346__23_, r_346__22_, r_346__21_, r_346__20_, r_346__19_, r_346__18_, r_346__17_, r_346__16_, r_346__15_, r_346__14_, r_346__13_, r_346__12_, r_346__11_, r_346__10_, r_346__9_, r_346__8_, r_346__7_, r_346__6_, r_346__5_, r_346__4_, r_346__3_, r_346__2_, r_346__1_, r_346__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N691)? data_i : 1'b0;
  assign N690 = sel_i[690];
  assign N691 = N2753;
  assign { r_n_346__63_, r_n_346__62_, r_n_346__61_, r_n_346__60_, r_n_346__59_, r_n_346__58_, r_n_346__57_, r_n_346__56_, r_n_346__55_, r_n_346__54_, r_n_346__53_, r_n_346__52_, r_n_346__51_, r_n_346__50_, r_n_346__49_, r_n_346__48_, r_n_346__47_, r_n_346__46_, r_n_346__45_, r_n_346__44_, r_n_346__43_, r_n_346__42_, r_n_346__41_, r_n_346__40_, r_n_346__39_, r_n_346__38_, r_n_346__37_, r_n_346__36_, r_n_346__35_, r_n_346__34_, r_n_346__33_, r_n_346__32_, r_n_346__31_, r_n_346__30_, r_n_346__29_, r_n_346__28_, r_n_346__27_, r_n_346__26_, r_n_346__25_, r_n_346__24_, r_n_346__23_, r_n_346__22_, r_n_346__21_, r_n_346__20_, r_n_346__19_, r_n_346__18_, r_n_346__17_, r_n_346__16_, r_n_346__15_, r_n_346__14_, r_n_346__13_, r_n_346__12_, r_n_346__11_, r_n_346__10_, r_n_346__9_, r_n_346__8_, r_n_346__7_, r_n_346__6_, r_n_346__5_, r_n_346__4_, r_n_346__3_, r_n_346__2_, r_n_346__1_, r_n_346__0_ } = (N692)? { r_347__63_, r_347__62_, r_347__61_, r_347__60_, r_347__59_, r_347__58_, r_347__57_, r_347__56_, r_347__55_, r_347__54_, r_347__53_, r_347__52_, r_347__51_, r_347__50_, r_347__49_, r_347__48_, r_347__47_, r_347__46_, r_347__45_, r_347__44_, r_347__43_, r_347__42_, r_347__41_, r_347__40_, r_347__39_, r_347__38_, r_347__37_, r_347__36_, r_347__35_, r_347__34_, r_347__33_, r_347__32_, r_347__31_, r_347__30_, r_347__29_, r_347__28_, r_347__27_, r_347__26_, r_347__25_, r_347__24_, r_347__23_, r_347__22_, r_347__21_, r_347__20_, r_347__19_, r_347__18_, r_347__17_, r_347__16_, r_347__15_, r_347__14_, r_347__13_, r_347__12_, r_347__11_, r_347__10_, r_347__9_, r_347__8_, r_347__7_, r_347__6_, r_347__5_, r_347__4_, r_347__3_, r_347__2_, r_347__1_, r_347__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N693)? data_i : 1'b0;
  assign N692 = sel_i[692];
  assign N693 = N2758;
  assign { r_n_347__63_, r_n_347__62_, r_n_347__61_, r_n_347__60_, r_n_347__59_, r_n_347__58_, r_n_347__57_, r_n_347__56_, r_n_347__55_, r_n_347__54_, r_n_347__53_, r_n_347__52_, r_n_347__51_, r_n_347__50_, r_n_347__49_, r_n_347__48_, r_n_347__47_, r_n_347__46_, r_n_347__45_, r_n_347__44_, r_n_347__43_, r_n_347__42_, r_n_347__41_, r_n_347__40_, r_n_347__39_, r_n_347__38_, r_n_347__37_, r_n_347__36_, r_n_347__35_, r_n_347__34_, r_n_347__33_, r_n_347__32_, r_n_347__31_, r_n_347__30_, r_n_347__29_, r_n_347__28_, r_n_347__27_, r_n_347__26_, r_n_347__25_, r_n_347__24_, r_n_347__23_, r_n_347__22_, r_n_347__21_, r_n_347__20_, r_n_347__19_, r_n_347__18_, r_n_347__17_, r_n_347__16_, r_n_347__15_, r_n_347__14_, r_n_347__13_, r_n_347__12_, r_n_347__11_, r_n_347__10_, r_n_347__9_, r_n_347__8_, r_n_347__7_, r_n_347__6_, r_n_347__5_, r_n_347__4_, r_n_347__3_, r_n_347__2_, r_n_347__1_, r_n_347__0_ } = (N694)? { r_348__63_, r_348__62_, r_348__61_, r_348__60_, r_348__59_, r_348__58_, r_348__57_, r_348__56_, r_348__55_, r_348__54_, r_348__53_, r_348__52_, r_348__51_, r_348__50_, r_348__49_, r_348__48_, r_348__47_, r_348__46_, r_348__45_, r_348__44_, r_348__43_, r_348__42_, r_348__41_, r_348__40_, r_348__39_, r_348__38_, r_348__37_, r_348__36_, r_348__35_, r_348__34_, r_348__33_, r_348__32_, r_348__31_, r_348__30_, r_348__29_, r_348__28_, r_348__27_, r_348__26_, r_348__25_, r_348__24_, r_348__23_, r_348__22_, r_348__21_, r_348__20_, r_348__19_, r_348__18_, r_348__17_, r_348__16_, r_348__15_, r_348__14_, r_348__13_, r_348__12_, r_348__11_, r_348__10_, r_348__9_, r_348__8_, r_348__7_, r_348__6_, r_348__5_, r_348__4_, r_348__3_, r_348__2_, r_348__1_, r_348__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N695)? data_i : 1'b0;
  assign N694 = sel_i[694];
  assign N695 = N2763;
  assign { r_n_348__63_, r_n_348__62_, r_n_348__61_, r_n_348__60_, r_n_348__59_, r_n_348__58_, r_n_348__57_, r_n_348__56_, r_n_348__55_, r_n_348__54_, r_n_348__53_, r_n_348__52_, r_n_348__51_, r_n_348__50_, r_n_348__49_, r_n_348__48_, r_n_348__47_, r_n_348__46_, r_n_348__45_, r_n_348__44_, r_n_348__43_, r_n_348__42_, r_n_348__41_, r_n_348__40_, r_n_348__39_, r_n_348__38_, r_n_348__37_, r_n_348__36_, r_n_348__35_, r_n_348__34_, r_n_348__33_, r_n_348__32_, r_n_348__31_, r_n_348__30_, r_n_348__29_, r_n_348__28_, r_n_348__27_, r_n_348__26_, r_n_348__25_, r_n_348__24_, r_n_348__23_, r_n_348__22_, r_n_348__21_, r_n_348__20_, r_n_348__19_, r_n_348__18_, r_n_348__17_, r_n_348__16_, r_n_348__15_, r_n_348__14_, r_n_348__13_, r_n_348__12_, r_n_348__11_, r_n_348__10_, r_n_348__9_, r_n_348__8_, r_n_348__7_, r_n_348__6_, r_n_348__5_, r_n_348__4_, r_n_348__3_, r_n_348__2_, r_n_348__1_, r_n_348__0_ } = (N696)? { r_349__63_, r_349__62_, r_349__61_, r_349__60_, r_349__59_, r_349__58_, r_349__57_, r_349__56_, r_349__55_, r_349__54_, r_349__53_, r_349__52_, r_349__51_, r_349__50_, r_349__49_, r_349__48_, r_349__47_, r_349__46_, r_349__45_, r_349__44_, r_349__43_, r_349__42_, r_349__41_, r_349__40_, r_349__39_, r_349__38_, r_349__37_, r_349__36_, r_349__35_, r_349__34_, r_349__33_, r_349__32_, r_349__31_, r_349__30_, r_349__29_, r_349__28_, r_349__27_, r_349__26_, r_349__25_, r_349__24_, r_349__23_, r_349__22_, r_349__21_, r_349__20_, r_349__19_, r_349__18_, r_349__17_, r_349__16_, r_349__15_, r_349__14_, r_349__13_, r_349__12_, r_349__11_, r_349__10_, r_349__9_, r_349__8_, r_349__7_, r_349__6_, r_349__5_, r_349__4_, r_349__3_, r_349__2_, r_349__1_, r_349__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N697)? data_i : 1'b0;
  assign N696 = sel_i[696];
  assign N697 = N2768;
  assign { r_n_349__63_, r_n_349__62_, r_n_349__61_, r_n_349__60_, r_n_349__59_, r_n_349__58_, r_n_349__57_, r_n_349__56_, r_n_349__55_, r_n_349__54_, r_n_349__53_, r_n_349__52_, r_n_349__51_, r_n_349__50_, r_n_349__49_, r_n_349__48_, r_n_349__47_, r_n_349__46_, r_n_349__45_, r_n_349__44_, r_n_349__43_, r_n_349__42_, r_n_349__41_, r_n_349__40_, r_n_349__39_, r_n_349__38_, r_n_349__37_, r_n_349__36_, r_n_349__35_, r_n_349__34_, r_n_349__33_, r_n_349__32_, r_n_349__31_, r_n_349__30_, r_n_349__29_, r_n_349__28_, r_n_349__27_, r_n_349__26_, r_n_349__25_, r_n_349__24_, r_n_349__23_, r_n_349__22_, r_n_349__21_, r_n_349__20_, r_n_349__19_, r_n_349__18_, r_n_349__17_, r_n_349__16_, r_n_349__15_, r_n_349__14_, r_n_349__13_, r_n_349__12_, r_n_349__11_, r_n_349__10_, r_n_349__9_, r_n_349__8_, r_n_349__7_, r_n_349__6_, r_n_349__5_, r_n_349__4_, r_n_349__3_, r_n_349__2_, r_n_349__1_, r_n_349__0_ } = (N698)? { r_350__63_, r_350__62_, r_350__61_, r_350__60_, r_350__59_, r_350__58_, r_350__57_, r_350__56_, r_350__55_, r_350__54_, r_350__53_, r_350__52_, r_350__51_, r_350__50_, r_350__49_, r_350__48_, r_350__47_, r_350__46_, r_350__45_, r_350__44_, r_350__43_, r_350__42_, r_350__41_, r_350__40_, r_350__39_, r_350__38_, r_350__37_, r_350__36_, r_350__35_, r_350__34_, r_350__33_, r_350__32_, r_350__31_, r_350__30_, r_350__29_, r_350__28_, r_350__27_, r_350__26_, r_350__25_, r_350__24_, r_350__23_, r_350__22_, r_350__21_, r_350__20_, r_350__19_, r_350__18_, r_350__17_, r_350__16_, r_350__15_, r_350__14_, r_350__13_, r_350__12_, r_350__11_, r_350__10_, r_350__9_, r_350__8_, r_350__7_, r_350__6_, r_350__5_, r_350__4_, r_350__3_, r_350__2_, r_350__1_, r_350__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N699)? data_i : 1'b0;
  assign N698 = sel_i[698];
  assign N699 = N2773;
  assign { r_n_350__63_, r_n_350__62_, r_n_350__61_, r_n_350__60_, r_n_350__59_, r_n_350__58_, r_n_350__57_, r_n_350__56_, r_n_350__55_, r_n_350__54_, r_n_350__53_, r_n_350__52_, r_n_350__51_, r_n_350__50_, r_n_350__49_, r_n_350__48_, r_n_350__47_, r_n_350__46_, r_n_350__45_, r_n_350__44_, r_n_350__43_, r_n_350__42_, r_n_350__41_, r_n_350__40_, r_n_350__39_, r_n_350__38_, r_n_350__37_, r_n_350__36_, r_n_350__35_, r_n_350__34_, r_n_350__33_, r_n_350__32_, r_n_350__31_, r_n_350__30_, r_n_350__29_, r_n_350__28_, r_n_350__27_, r_n_350__26_, r_n_350__25_, r_n_350__24_, r_n_350__23_, r_n_350__22_, r_n_350__21_, r_n_350__20_, r_n_350__19_, r_n_350__18_, r_n_350__17_, r_n_350__16_, r_n_350__15_, r_n_350__14_, r_n_350__13_, r_n_350__12_, r_n_350__11_, r_n_350__10_, r_n_350__9_, r_n_350__8_, r_n_350__7_, r_n_350__6_, r_n_350__5_, r_n_350__4_, r_n_350__3_, r_n_350__2_, r_n_350__1_, r_n_350__0_ } = (N700)? { r_351__63_, r_351__62_, r_351__61_, r_351__60_, r_351__59_, r_351__58_, r_351__57_, r_351__56_, r_351__55_, r_351__54_, r_351__53_, r_351__52_, r_351__51_, r_351__50_, r_351__49_, r_351__48_, r_351__47_, r_351__46_, r_351__45_, r_351__44_, r_351__43_, r_351__42_, r_351__41_, r_351__40_, r_351__39_, r_351__38_, r_351__37_, r_351__36_, r_351__35_, r_351__34_, r_351__33_, r_351__32_, r_351__31_, r_351__30_, r_351__29_, r_351__28_, r_351__27_, r_351__26_, r_351__25_, r_351__24_, r_351__23_, r_351__22_, r_351__21_, r_351__20_, r_351__19_, r_351__18_, r_351__17_, r_351__16_, r_351__15_, r_351__14_, r_351__13_, r_351__12_, r_351__11_, r_351__10_, r_351__9_, r_351__8_, r_351__7_, r_351__6_, r_351__5_, r_351__4_, r_351__3_, r_351__2_, r_351__1_, r_351__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N701)? data_i : 1'b0;
  assign N700 = sel_i[700];
  assign N701 = N2778;
  assign { r_n_351__63_, r_n_351__62_, r_n_351__61_, r_n_351__60_, r_n_351__59_, r_n_351__58_, r_n_351__57_, r_n_351__56_, r_n_351__55_, r_n_351__54_, r_n_351__53_, r_n_351__52_, r_n_351__51_, r_n_351__50_, r_n_351__49_, r_n_351__48_, r_n_351__47_, r_n_351__46_, r_n_351__45_, r_n_351__44_, r_n_351__43_, r_n_351__42_, r_n_351__41_, r_n_351__40_, r_n_351__39_, r_n_351__38_, r_n_351__37_, r_n_351__36_, r_n_351__35_, r_n_351__34_, r_n_351__33_, r_n_351__32_, r_n_351__31_, r_n_351__30_, r_n_351__29_, r_n_351__28_, r_n_351__27_, r_n_351__26_, r_n_351__25_, r_n_351__24_, r_n_351__23_, r_n_351__22_, r_n_351__21_, r_n_351__20_, r_n_351__19_, r_n_351__18_, r_n_351__17_, r_n_351__16_, r_n_351__15_, r_n_351__14_, r_n_351__13_, r_n_351__12_, r_n_351__11_, r_n_351__10_, r_n_351__9_, r_n_351__8_, r_n_351__7_, r_n_351__6_, r_n_351__5_, r_n_351__4_, r_n_351__3_, r_n_351__2_, r_n_351__1_, r_n_351__0_ } = (N702)? { r_352__63_, r_352__62_, r_352__61_, r_352__60_, r_352__59_, r_352__58_, r_352__57_, r_352__56_, r_352__55_, r_352__54_, r_352__53_, r_352__52_, r_352__51_, r_352__50_, r_352__49_, r_352__48_, r_352__47_, r_352__46_, r_352__45_, r_352__44_, r_352__43_, r_352__42_, r_352__41_, r_352__40_, r_352__39_, r_352__38_, r_352__37_, r_352__36_, r_352__35_, r_352__34_, r_352__33_, r_352__32_, r_352__31_, r_352__30_, r_352__29_, r_352__28_, r_352__27_, r_352__26_, r_352__25_, r_352__24_, r_352__23_, r_352__22_, r_352__21_, r_352__20_, r_352__19_, r_352__18_, r_352__17_, r_352__16_, r_352__15_, r_352__14_, r_352__13_, r_352__12_, r_352__11_, r_352__10_, r_352__9_, r_352__8_, r_352__7_, r_352__6_, r_352__5_, r_352__4_, r_352__3_, r_352__2_, r_352__1_, r_352__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N703)? data_i : 1'b0;
  assign N702 = sel_i[702];
  assign N703 = N2783;
  assign { r_n_352__63_, r_n_352__62_, r_n_352__61_, r_n_352__60_, r_n_352__59_, r_n_352__58_, r_n_352__57_, r_n_352__56_, r_n_352__55_, r_n_352__54_, r_n_352__53_, r_n_352__52_, r_n_352__51_, r_n_352__50_, r_n_352__49_, r_n_352__48_, r_n_352__47_, r_n_352__46_, r_n_352__45_, r_n_352__44_, r_n_352__43_, r_n_352__42_, r_n_352__41_, r_n_352__40_, r_n_352__39_, r_n_352__38_, r_n_352__37_, r_n_352__36_, r_n_352__35_, r_n_352__34_, r_n_352__33_, r_n_352__32_, r_n_352__31_, r_n_352__30_, r_n_352__29_, r_n_352__28_, r_n_352__27_, r_n_352__26_, r_n_352__25_, r_n_352__24_, r_n_352__23_, r_n_352__22_, r_n_352__21_, r_n_352__20_, r_n_352__19_, r_n_352__18_, r_n_352__17_, r_n_352__16_, r_n_352__15_, r_n_352__14_, r_n_352__13_, r_n_352__12_, r_n_352__11_, r_n_352__10_, r_n_352__9_, r_n_352__8_, r_n_352__7_, r_n_352__6_, r_n_352__5_, r_n_352__4_, r_n_352__3_, r_n_352__2_, r_n_352__1_, r_n_352__0_ } = (N704)? { r_353__63_, r_353__62_, r_353__61_, r_353__60_, r_353__59_, r_353__58_, r_353__57_, r_353__56_, r_353__55_, r_353__54_, r_353__53_, r_353__52_, r_353__51_, r_353__50_, r_353__49_, r_353__48_, r_353__47_, r_353__46_, r_353__45_, r_353__44_, r_353__43_, r_353__42_, r_353__41_, r_353__40_, r_353__39_, r_353__38_, r_353__37_, r_353__36_, r_353__35_, r_353__34_, r_353__33_, r_353__32_, r_353__31_, r_353__30_, r_353__29_, r_353__28_, r_353__27_, r_353__26_, r_353__25_, r_353__24_, r_353__23_, r_353__22_, r_353__21_, r_353__20_, r_353__19_, r_353__18_, r_353__17_, r_353__16_, r_353__15_, r_353__14_, r_353__13_, r_353__12_, r_353__11_, r_353__10_, r_353__9_, r_353__8_, r_353__7_, r_353__6_, r_353__5_, r_353__4_, r_353__3_, r_353__2_, r_353__1_, r_353__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N705)? data_i : 1'b0;
  assign N704 = sel_i[704];
  assign N705 = N2788;
  assign { r_n_353__63_, r_n_353__62_, r_n_353__61_, r_n_353__60_, r_n_353__59_, r_n_353__58_, r_n_353__57_, r_n_353__56_, r_n_353__55_, r_n_353__54_, r_n_353__53_, r_n_353__52_, r_n_353__51_, r_n_353__50_, r_n_353__49_, r_n_353__48_, r_n_353__47_, r_n_353__46_, r_n_353__45_, r_n_353__44_, r_n_353__43_, r_n_353__42_, r_n_353__41_, r_n_353__40_, r_n_353__39_, r_n_353__38_, r_n_353__37_, r_n_353__36_, r_n_353__35_, r_n_353__34_, r_n_353__33_, r_n_353__32_, r_n_353__31_, r_n_353__30_, r_n_353__29_, r_n_353__28_, r_n_353__27_, r_n_353__26_, r_n_353__25_, r_n_353__24_, r_n_353__23_, r_n_353__22_, r_n_353__21_, r_n_353__20_, r_n_353__19_, r_n_353__18_, r_n_353__17_, r_n_353__16_, r_n_353__15_, r_n_353__14_, r_n_353__13_, r_n_353__12_, r_n_353__11_, r_n_353__10_, r_n_353__9_, r_n_353__8_, r_n_353__7_, r_n_353__6_, r_n_353__5_, r_n_353__4_, r_n_353__3_, r_n_353__2_, r_n_353__1_, r_n_353__0_ } = (N706)? { r_354__63_, r_354__62_, r_354__61_, r_354__60_, r_354__59_, r_354__58_, r_354__57_, r_354__56_, r_354__55_, r_354__54_, r_354__53_, r_354__52_, r_354__51_, r_354__50_, r_354__49_, r_354__48_, r_354__47_, r_354__46_, r_354__45_, r_354__44_, r_354__43_, r_354__42_, r_354__41_, r_354__40_, r_354__39_, r_354__38_, r_354__37_, r_354__36_, r_354__35_, r_354__34_, r_354__33_, r_354__32_, r_354__31_, r_354__30_, r_354__29_, r_354__28_, r_354__27_, r_354__26_, r_354__25_, r_354__24_, r_354__23_, r_354__22_, r_354__21_, r_354__20_, r_354__19_, r_354__18_, r_354__17_, r_354__16_, r_354__15_, r_354__14_, r_354__13_, r_354__12_, r_354__11_, r_354__10_, r_354__9_, r_354__8_, r_354__7_, r_354__6_, r_354__5_, r_354__4_, r_354__3_, r_354__2_, r_354__1_, r_354__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N707)? data_i : 1'b0;
  assign N706 = sel_i[706];
  assign N707 = N2793;
  assign { r_n_354__63_, r_n_354__62_, r_n_354__61_, r_n_354__60_, r_n_354__59_, r_n_354__58_, r_n_354__57_, r_n_354__56_, r_n_354__55_, r_n_354__54_, r_n_354__53_, r_n_354__52_, r_n_354__51_, r_n_354__50_, r_n_354__49_, r_n_354__48_, r_n_354__47_, r_n_354__46_, r_n_354__45_, r_n_354__44_, r_n_354__43_, r_n_354__42_, r_n_354__41_, r_n_354__40_, r_n_354__39_, r_n_354__38_, r_n_354__37_, r_n_354__36_, r_n_354__35_, r_n_354__34_, r_n_354__33_, r_n_354__32_, r_n_354__31_, r_n_354__30_, r_n_354__29_, r_n_354__28_, r_n_354__27_, r_n_354__26_, r_n_354__25_, r_n_354__24_, r_n_354__23_, r_n_354__22_, r_n_354__21_, r_n_354__20_, r_n_354__19_, r_n_354__18_, r_n_354__17_, r_n_354__16_, r_n_354__15_, r_n_354__14_, r_n_354__13_, r_n_354__12_, r_n_354__11_, r_n_354__10_, r_n_354__9_, r_n_354__8_, r_n_354__7_, r_n_354__6_, r_n_354__5_, r_n_354__4_, r_n_354__3_, r_n_354__2_, r_n_354__1_, r_n_354__0_ } = (N708)? { r_355__63_, r_355__62_, r_355__61_, r_355__60_, r_355__59_, r_355__58_, r_355__57_, r_355__56_, r_355__55_, r_355__54_, r_355__53_, r_355__52_, r_355__51_, r_355__50_, r_355__49_, r_355__48_, r_355__47_, r_355__46_, r_355__45_, r_355__44_, r_355__43_, r_355__42_, r_355__41_, r_355__40_, r_355__39_, r_355__38_, r_355__37_, r_355__36_, r_355__35_, r_355__34_, r_355__33_, r_355__32_, r_355__31_, r_355__30_, r_355__29_, r_355__28_, r_355__27_, r_355__26_, r_355__25_, r_355__24_, r_355__23_, r_355__22_, r_355__21_, r_355__20_, r_355__19_, r_355__18_, r_355__17_, r_355__16_, r_355__15_, r_355__14_, r_355__13_, r_355__12_, r_355__11_, r_355__10_, r_355__9_, r_355__8_, r_355__7_, r_355__6_, r_355__5_, r_355__4_, r_355__3_, r_355__2_, r_355__1_, r_355__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N709)? data_i : 1'b0;
  assign N708 = sel_i[708];
  assign N709 = N2798;
  assign { r_n_355__63_, r_n_355__62_, r_n_355__61_, r_n_355__60_, r_n_355__59_, r_n_355__58_, r_n_355__57_, r_n_355__56_, r_n_355__55_, r_n_355__54_, r_n_355__53_, r_n_355__52_, r_n_355__51_, r_n_355__50_, r_n_355__49_, r_n_355__48_, r_n_355__47_, r_n_355__46_, r_n_355__45_, r_n_355__44_, r_n_355__43_, r_n_355__42_, r_n_355__41_, r_n_355__40_, r_n_355__39_, r_n_355__38_, r_n_355__37_, r_n_355__36_, r_n_355__35_, r_n_355__34_, r_n_355__33_, r_n_355__32_, r_n_355__31_, r_n_355__30_, r_n_355__29_, r_n_355__28_, r_n_355__27_, r_n_355__26_, r_n_355__25_, r_n_355__24_, r_n_355__23_, r_n_355__22_, r_n_355__21_, r_n_355__20_, r_n_355__19_, r_n_355__18_, r_n_355__17_, r_n_355__16_, r_n_355__15_, r_n_355__14_, r_n_355__13_, r_n_355__12_, r_n_355__11_, r_n_355__10_, r_n_355__9_, r_n_355__8_, r_n_355__7_, r_n_355__6_, r_n_355__5_, r_n_355__4_, r_n_355__3_, r_n_355__2_, r_n_355__1_, r_n_355__0_ } = (N710)? { r_356__63_, r_356__62_, r_356__61_, r_356__60_, r_356__59_, r_356__58_, r_356__57_, r_356__56_, r_356__55_, r_356__54_, r_356__53_, r_356__52_, r_356__51_, r_356__50_, r_356__49_, r_356__48_, r_356__47_, r_356__46_, r_356__45_, r_356__44_, r_356__43_, r_356__42_, r_356__41_, r_356__40_, r_356__39_, r_356__38_, r_356__37_, r_356__36_, r_356__35_, r_356__34_, r_356__33_, r_356__32_, r_356__31_, r_356__30_, r_356__29_, r_356__28_, r_356__27_, r_356__26_, r_356__25_, r_356__24_, r_356__23_, r_356__22_, r_356__21_, r_356__20_, r_356__19_, r_356__18_, r_356__17_, r_356__16_, r_356__15_, r_356__14_, r_356__13_, r_356__12_, r_356__11_, r_356__10_, r_356__9_, r_356__8_, r_356__7_, r_356__6_, r_356__5_, r_356__4_, r_356__3_, r_356__2_, r_356__1_, r_356__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N711)? data_i : 1'b0;
  assign N710 = sel_i[710];
  assign N711 = N2803;
  assign { r_n_356__63_, r_n_356__62_, r_n_356__61_, r_n_356__60_, r_n_356__59_, r_n_356__58_, r_n_356__57_, r_n_356__56_, r_n_356__55_, r_n_356__54_, r_n_356__53_, r_n_356__52_, r_n_356__51_, r_n_356__50_, r_n_356__49_, r_n_356__48_, r_n_356__47_, r_n_356__46_, r_n_356__45_, r_n_356__44_, r_n_356__43_, r_n_356__42_, r_n_356__41_, r_n_356__40_, r_n_356__39_, r_n_356__38_, r_n_356__37_, r_n_356__36_, r_n_356__35_, r_n_356__34_, r_n_356__33_, r_n_356__32_, r_n_356__31_, r_n_356__30_, r_n_356__29_, r_n_356__28_, r_n_356__27_, r_n_356__26_, r_n_356__25_, r_n_356__24_, r_n_356__23_, r_n_356__22_, r_n_356__21_, r_n_356__20_, r_n_356__19_, r_n_356__18_, r_n_356__17_, r_n_356__16_, r_n_356__15_, r_n_356__14_, r_n_356__13_, r_n_356__12_, r_n_356__11_, r_n_356__10_, r_n_356__9_, r_n_356__8_, r_n_356__7_, r_n_356__6_, r_n_356__5_, r_n_356__4_, r_n_356__3_, r_n_356__2_, r_n_356__1_, r_n_356__0_ } = (N712)? { r_357__63_, r_357__62_, r_357__61_, r_357__60_, r_357__59_, r_357__58_, r_357__57_, r_357__56_, r_357__55_, r_357__54_, r_357__53_, r_357__52_, r_357__51_, r_357__50_, r_357__49_, r_357__48_, r_357__47_, r_357__46_, r_357__45_, r_357__44_, r_357__43_, r_357__42_, r_357__41_, r_357__40_, r_357__39_, r_357__38_, r_357__37_, r_357__36_, r_357__35_, r_357__34_, r_357__33_, r_357__32_, r_357__31_, r_357__30_, r_357__29_, r_357__28_, r_357__27_, r_357__26_, r_357__25_, r_357__24_, r_357__23_, r_357__22_, r_357__21_, r_357__20_, r_357__19_, r_357__18_, r_357__17_, r_357__16_, r_357__15_, r_357__14_, r_357__13_, r_357__12_, r_357__11_, r_357__10_, r_357__9_, r_357__8_, r_357__7_, r_357__6_, r_357__5_, r_357__4_, r_357__3_, r_357__2_, r_357__1_, r_357__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N713)? data_i : 1'b0;
  assign N712 = sel_i[712];
  assign N713 = N2808;
  assign { r_n_357__63_, r_n_357__62_, r_n_357__61_, r_n_357__60_, r_n_357__59_, r_n_357__58_, r_n_357__57_, r_n_357__56_, r_n_357__55_, r_n_357__54_, r_n_357__53_, r_n_357__52_, r_n_357__51_, r_n_357__50_, r_n_357__49_, r_n_357__48_, r_n_357__47_, r_n_357__46_, r_n_357__45_, r_n_357__44_, r_n_357__43_, r_n_357__42_, r_n_357__41_, r_n_357__40_, r_n_357__39_, r_n_357__38_, r_n_357__37_, r_n_357__36_, r_n_357__35_, r_n_357__34_, r_n_357__33_, r_n_357__32_, r_n_357__31_, r_n_357__30_, r_n_357__29_, r_n_357__28_, r_n_357__27_, r_n_357__26_, r_n_357__25_, r_n_357__24_, r_n_357__23_, r_n_357__22_, r_n_357__21_, r_n_357__20_, r_n_357__19_, r_n_357__18_, r_n_357__17_, r_n_357__16_, r_n_357__15_, r_n_357__14_, r_n_357__13_, r_n_357__12_, r_n_357__11_, r_n_357__10_, r_n_357__9_, r_n_357__8_, r_n_357__7_, r_n_357__6_, r_n_357__5_, r_n_357__4_, r_n_357__3_, r_n_357__2_, r_n_357__1_, r_n_357__0_ } = (N714)? { r_358__63_, r_358__62_, r_358__61_, r_358__60_, r_358__59_, r_358__58_, r_358__57_, r_358__56_, r_358__55_, r_358__54_, r_358__53_, r_358__52_, r_358__51_, r_358__50_, r_358__49_, r_358__48_, r_358__47_, r_358__46_, r_358__45_, r_358__44_, r_358__43_, r_358__42_, r_358__41_, r_358__40_, r_358__39_, r_358__38_, r_358__37_, r_358__36_, r_358__35_, r_358__34_, r_358__33_, r_358__32_, r_358__31_, r_358__30_, r_358__29_, r_358__28_, r_358__27_, r_358__26_, r_358__25_, r_358__24_, r_358__23_, r_358__22_, r_358__21_, r_358__20_, r_358__19_, r_358__18_, r_358__17_, r_358__16_, r_358__15_, r_358__14_, r_358__13_, r_358__12_, r_358__11_, r_358__10_, r_358__9_, r_358__8_, r_358__7_, r_358__6_, r_358__5_, r_358__4_, r_358__3_, r_358__2_, r_358__1_, r_358__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N715)? data_i : 1'b0;
  assign N714 = sel_i[714];
  assign N715 = N2813;
  assign { r_n_358__63_, r_n_358__62_, r_n_358__61_, r_n_358__60_, r_n_358__59_, r_n_358__58_, r_n_358__57_, r_n_358__56_, r_n_358__55_, r_n_358__54_, r_n_358__53_, r_n_358__52_, r_n_358__51_, r_n_358__50_, r_n_358__49_, r_n_358__48_, r_n_358__47_, r_n_358__46_, r_n_358__45_, r_n_358__44_, r_n_358__43_, r_n_358__42_, r_n_358__41_, r_n_358__40_, r_n_358__39_, r_n_358__38_, r_n_358__37_, r_n_358__36_, r_n_358__35_, r_n_358__34_, r_n_358__33_, r_n_358__32_, r_n_358__31_, r_n_358__30_, r_n_358__29_, r_n_358__28_, r_n_358__27_, r_n_358__26_, r_n_358__25_, r_n_358__24_, r_n_358__23_, r_n_358__22_, r_n_358__21_, r_n_358__20_, r_n_358__19_, r_n_358__18_, r_n_358__17_, r_n_358__16_, r_n_358__15_, r_n_358__14_, r_n_358__13_, r_n_358__12_, r_n_358__11_, r_n_358__10_, r_n_358__9_, r_n_358__8_, r_n_358__7_, r_n_358__6_, r_n_358__5_, r_n_358__4_, r_n_358__3_, r_n_358__2_, r_n_358__1_, r_n_358__0_ } = (N716)? { r_359__63_, r_359__62_, r_359__61_, r_359__60_, r_359__59_, r_359__58_, r_359__57_, r_359__56_, r_359__55_, r_359__54_, r_359__53_, r_359__52_, r_359__51_, r_359__50_, r_359__49_, r_359__48_, r_359__47_, r_359__46_, r_359__45_, r_359__44_, r_359__43_, r_359__42_, r_359__41_, r_359__40_, r_359__39_, r_359__38_, r_359__37_, r_359__36_, r_359__35_, r_359__34_, r_359__33_, r_359__32_, r_359__31_, r_359__30_, r_359__29_, r_359__28_, r_359__27_, r_359__26_, r_359__25_, r_359__24_, r_359__23_, r_359__22_, r_359__21_, r_359__20_, r_359__19_, r_359__18_, r_359__17_, r_359__16_, r_359__15_, r_359__14_, r_359__13_, r_359__12_, r_359__11_, r_359__10_, r_359__9_, r_359__8_, r_359__7_, r_359__6_, r_359__5_, r_359__4_, r_359__3_, r_359__2_, r_359__1_, r_359__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N717)? data_i : 1'b0;
  assign N716 = sel_i[716];
  assign N717 = N2818;
  assign { r_n_359__63_, r_n_359__62_, r_n_359__61_, r_n_359__60_, r_n_359__59_, r_n_359__58_, r_n_359__57_, r_n_359__56_, r_n_359__55_, r_n_359__54_, r_n_359__53_, r_n_359__52_, r_n_359__51_, r_n_359__50_, r_n_359__49_, r_n_359__48_, r_n_359__47_, r_n_359__46_, r_n_359__45_, r_n_359__44_, r_n_359__43_, r_n_359__42_, r_n_359__41_, r_n_359__40_, r_n_359__39_, r_n_359__38_, r_n_359__37_, r_n_359__36_, r_n_359__35_, r_n_359__34_, r_n_359__33_, r_n_359__32_, r_n_359__31_, r_n_359__30_, r_n_359__29_, r_n_359__28_, r_n_359__27_, r_n_359__26_, r_n_359__25_, r_n_359__24_, r_n_359__23_, r_n_359__22_, r_n_359__21_, r_n_359__20_, r_n_359__19_, r_n_359__18_, r_n_359__17_, r_n_359__16_, r_n_359__15_, r_n_359__14_, r_n_359__13_, r_n_359__12_, r_n_359__11_, r_n_359__10_, r_n_359__9_, r_n_359__8_, r_n_359__7_, r_n_359__6_, r_n_359__5_, r_n_359__4_, r_n_359__3_, r_n_359__2_, r_n_359__1_, r_n_359__0_ } = (N718)? { r_360__63_, r_360__62_, r_360__61_, r_360__60_, r_360__59_, r_360__58_, r_360__57_, r_360__56_, r_360__55_, r_360__54_, r_360__53_, r_360__52_, r_360__51_, r_360__50_, r_360__49_, r_360__48_, r_360__47_, r_360__46_, r_360__45_, r_360__44_, r_360__43_, r_360__42_, r_360__41_, r_360__40_, r_360__39_, r_360__38_, r_360__37_, r_360__36_, r_360__35_, r_360__34_, r_360__33_, r_360__32_, r_360__31_, r_360__30_, r_360__29_, r_360__28_, r_360__27_, r_360__26_, r_360__25_, r_360__24_, r_360__23_, r_360__22_, r_360__21_, r_360__20_, r_360__19_, r_360__18_, r_360__17_, r_360__16_, r_360__15_, r_360__14_, r_360__13_, r_360__12_, r_360__11_, r_360__10_, r_360__9_, r_360__8_, r_360__7_, r_360__6_, r_360__5_, r_360__4_, r_360__3_, r_360__2_, r_360__1_, r_360__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N719)? data_i : 1'b0;
  assign N718 = sel_i[718];
  assign N719 = N2823;
  assign { r_n_360__63_, r_n_360__62_, r_n_360__61_, r_n_360__60_, r_n_360__59_, r_n_360__58_, r_n_360__57_, r_n_360__56_, r_n_360__55_, r_n_360__54_, r_n_360__53_, r_n_360__52_, r_n_360__51_, r_n_360__50_, r_n_360__49_, r_n_360__48_, r_n_360__47_, r_n_360__46_, r_n_360__45_, r_n_360__44_, r_n_360__43_, r_n_360__42_, r_n_360__41_, r_n_360__40_, r_n_360__39_, r_n_360__38_, r_n_360__37_, r_n_360__36_, r_n_360__35_, r_n_360__34_, r_n_360__33_, r_n_360__32_, r_n_360__31_, r_n_360__30_, r_n_360__29_, r_n_360__28_, r_n_360__27_, r_n_360__26_, r_n_360__25_, r_n_360__24_, r_n_360__23_, r_n_360__22_, r_n_360__21_, r_n_360__20_, r_n_360__19_, r_n_360__18_, r_n_360__17_, r_n_360__16_, r_n_360__15_, r_n_360__14_, r_n_360__13_, r_n_360__12_, r_n_360__11_, r_n_360__10_, r_n_360__9_, r_n_360__8_, r_n_360__7_, r_n_360__6_, r_n_360__5_, r_n_360__4_, r_n_360__3_, r_n_360__2_, r_n_360__1_, r_n_360__0_ } = (N720)? { r_361__63_, r_361__62_, r_361__61_, r_361__60_, r_361__59_, r_361__58_, r_361__57_, r_361__56_, r_361__55_, r_361__54_, r_361__53_, r_361__52_, r_361__51_, r_361__50_, r_361__49_, r_361__48_, r_361__47_, r_361__46_, r_361__45_, r_361__44_, r_361__43_, r_361__42_, r_361__41_, r_361__40_, r_361__39_, r_361__38_, r_361__37_, r_361__36_, r_361__35_, r_361__34_, r_361__33_, r_361__32_, r_361__31_, r_361__30_, r_361__29_, r_361__28_, r_361__27_, r_361__26_, r_361__25_, r_361__24_, r_361__23_, r_361__22_, r_361__21_, r_361__20_, r_361__19_, r_361__18_, r_361__17_, r_361__16_, r_361__15_, r_361__14_, r_361__13_, r_361__12_, r_361__11_, r_361__10_, r_361__9_, r_361__8_, r_361__7_, r_361__6_, r_361__5_, r_361__4_, r_361__3_, r_361__2_, r_361__1_, r_361__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N721)? data_i : 1'b0;
  assign N720 = sel_i[720];
  assign N721 = N2828;
  assign { r_n_361__63_, r_n_361__62_, r_n_361__61_, r_n_361__60_, r_n_361__59_, r_n_361__58_, r_n_361__57_, r_n_361__56_, r_n_361__55_, r_n_361__54_, r_n_361__53_, r_n_361__52_, r_n_361__51_, r_n_361__50_, r_n_361__49_, r_n_361__48_, r_n_361__47_, r_n_361__46_, r_n_361__45_, r_n_361__44_, r_n_361__43_, r_n_361__42_, r_n_361__41_, r_n_361__40_, r_n_361__39_, r_n_361__38_, r_n_361__37_, r_n_361__36_, r_n_361__35_, r_n_361__34_, r_n_361__33_, r_n_361__32_, r_n_361__31_, r_n_361__30_, r_n_361__29_, r_n_361__28_, r_n_361__27_, r_n_361__26_, r_n_361__25_, r_n_361__24_, r_n_361__23_, r_n_361__22_, r_n_361__21_, r_n_361__20_, r_n_361__19_, r_n_361__18_, r_n_361__17_, r_n_361__16_, r_n_361__15_, r_n_361__14_, r_n_361__13_, r_n_361__12_, r_n_361__11_, r_n_361__10_, r_n_361__9_, r_n_361__8_, r_n_361__7_, r_n_361__6_, r_n_361__5_, r_n_361__4_, r_n_361__3_, r_n_361__2_, r_n_361__1_, r_n_361__0_ } = (N722)? { r_362__63_, r_362__62_, r_362__61_, r_362__60_, r_362__59_, r_362__58_, r_362__57_, r_362__56_, r_362__55_, r_362__54_, r_362__53_, r_362__52_, r_362__51_, r_362__50_, r_362__49_, r_362__48_, r_362__47_, r_362__46_, r_362__45_, r_362__44_, r_362__43_, r_362__42_, r_362__41_, r_362__40_, r_362__39_, r_362__38_, r_362__37_, r_362__36_, r_362__35_, r_362__34_, r_362__33_, r_362__32_, r_362__31_, r_362__30_, r_362__29_, r_362__28_, r_362__27_, r_362__26_, r_362__25_, r_362__24_, r_362__23_, r_362__22_, r_362__21_, r_362__20_, r_362__19_, r_362__18_, r_362__17_, r_362__16_, r_362__15_, r_362__14_, r_362__13_, r_362__12_, r_362__11_, r_362__10_, r_362__9_, r_362__8_, r_362__7_, r_362__6_, r_362__5_, r_362__4_, r_362__3_, r_362__2_, r_362__1_, r_362__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N723)? data_i : 1'b0;
  assign N722 = sel_i[722];
  assign N723 = N2833;
  assign { r_n_362__63_, r_n_362__62_, r_n_362__61_, r_n_362__60_, r_n_362__59_, r_n_362__58_, r_n_362__57_, r_n_362__56_, r_n_362__55_, r_n_362__54_, r_n_362__53_, r_n_362__52_, r_n_362__51_, r_n_362__50_, r_n_362__49_, r_n_362__48_, r_n_362__47_, r_n_362__46_, r_n_362__45_, r_n_362__44_, r_n_362__43_, r_n_362__42_, r_n_362__41_, r_n_362__40_, r_n_362__39_, r_n_362__38_, r_n_362__37_, r_n_362__36_, r_n_362__35_, r_n_362__34_, r_n_362__33_, r_n_362__32_, r_n_362__31_, r_n_362__30_, r_n_362__29_, r_n_362__28_, r_n_362__27_, r_n_362__26_, r_n_362__25_, r_n_362__24_, r_n_362__23_, r_n_362__22_, r_n_362__21_, r_n_362__20_, r_n_362__19_, r_n_362__18_, r_n_362__17_, r_n_362__16_, r_n_362__15_, r_n_362__14_, r_n_362__13_, r_n_362__12_, r_n_362__11_, r_n_362__10_, r_n_362__9_, r_n_362__8_, r_n_362__7_, r_n_362__6_, r_n_362__5_, r_n_362__4_, r_n_362__3_, r_n_362__2_, r_n_362__1_, r_n_362__0_ } = (N724)? { r_363__63_, r_363__62_, r_363__61_, r_363__60_, r_363__59_, r_363__58_, r_363__57_, r_363__56_, r_363__55_, r_363__54_, r_363__53_, r_363__52_, r_363__51_, r_363__50_, r_363__49_, r_363__48_, r_363__47_, r_363__46_, r_363__45_, r_363__44_, r_363__43_, r_363__42_, r_363__41_, r_363__40_, r_363__39_, r_363__38_, r_363__37_, r_363__36_, r_363__35_, r_363__34_, r_363__33_, r_363__32_, r_363__31_, r_363__30_, r_363__29_, r_363__28_, r_363__27_, r_363__26_, r_363__25_, r_363__24_, r_363__23_, r_363__22_, r_363__21_, r_363__20_, r_363__19_, r_363__18_, r_363__17_, r_363__16_, r_363__15_, r_363__14_, r_363__13_, r_363__12_, r_363__11_, r_363__10_, r_363__9_, r_363__8_, r_363__7_, r_363__6_, r_363__5_, r_363__4_, r_363__3_, r_363__2_, r_363__1_, r_363__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N725)? data_i : 1'b0;
  assign N724 = sel_i[724];
  assign N725 = N2838;
  assign { r_n_363__63_, r_n_363__62_, r_n_363__61_, r_n_363__60_, r_n_363__59_, r_n_363__58_, r_n_363__57_, r_n_363__56_, r_n_363__55_, r_n_363__54_, r_n_363__53_, r_n_363__52_, r_n_363__51_, r_n_363__50_, r_n_363__49_, r_n_363__48_, r_n_363__47_, r_n_363__46_, r_n_363__45_, r_n_363__44_, r_n_363__43_, r_n_363__42_, r_n_363__41_, r_n_363__40_, r_n_363__39_, r_n_363__38_, r_n_363__37_, r_n_363__36_, r_n_363__35_, r_n_363__34_, r_n_363__33_, r_n_363__32_, r_n_363__31_, r_n_363__30_, r_n_363__29_, r_n_363__28_, r_n_363__27_, r_n_363__26_, r_n_363__25_, r_n_363__24_, r_n_363__23_, r_n_363__22_, r_n_363__21_, r_n_363__20_, r_n_363__19_, r_n_363__18_, r_n_363__17_, r_n_363__16_, r_n_363__15_, r_n_363__14_, r_n_363__13_, r_n_363__12_, r_n_363__11_, r_n_363__10_, r_n_363__9_, r_n_363__8_, r_n_363__7_, r_n_363__6_, r_n_363__5_, r_n_363__4_, r_n_363__3_, r_n_363__2_, r_n_363__1_, r_n_363__0_ } = (N726)? { r_364__63_, r_364__62_, r_364__61_, r_364__60_, r_364__59_, r_364__58_, r_364__57_, r_364__56_, r_364__55_, r_364__54_, r_364__53_, r_364__52_, r_364__51_, r_364__50_, r_364__49_, r_364__48_, r_364__47_, r_364__46_, r_364__45_, r_364__44_, r_364__43_, r_364__42_, r_364__41_, r_364__40_, r_364__39_, r_364__38_, r_364__37_, r_364__36_, r_364__35_, r_364__34_, r_364__33_, r_364__32_, r_364__31_, r_364__30_, r_364__29_, r_364__28_, r_364__27_, r_364__26_, r_364__25_, r_364__24_, r_364__23_, r_364__22_, r_364__21_, r_364__20_, r_364__19_, r_364__18_, r_364__17_, r_364__16_, r_364__15_, r_364__14_, r_364__13_, r_364__12_, r_364__11_, r_364__10_, r_364__9_, r_364__8_, r_364__7_, r_364__6_, r_364__5_, r_364__4_, r_364__3_, r_364__2_, r_364__1_, r_364__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N727)? data_i : 1'b0;
  assign N726 = sel_i[726];
  assign N727 = N2843;
  assign { r_n_364__63_, r_n_364__62_, r_n_364__61_, r_n_364__60_, r_n_364__59_, r_n_364__58_, r_n_364__57_, r_n_364__56_, r_n_364__55_, r_n_364__54_, r_n_364__53_, r_n_364__52_, r_n_364__51_, r_n_364__50_, r_n_364__49_, r_n_364__48_, r_n_364__47_, r_n_364__46_, r_n_364__45_, r_n_364__44_, r_n_364__43_, r_n_364__42_, r_n_364__41_, r_n_364__40_, r_n_364__39_, r_n_364__38_, r_n_364__37_, r_n_364__36_, r_n_364__35_, r_n_364__34_, r_n_364__33_, r_n_364__32_, r_n_364__31_, r_n_364__30_, r_n_364__29_, r_n_364__28_, r_n_364__27_, r_n_364__26_, r_n_364__25_, r_n_364__24_, r_n_364__23_, r_n_364__22_, r_n_364__21_, r_n_364__20_, r_n_364__19_, r_n_364__18_, r_n_364__17_, r_n_364__16_, r_n_364__15_, r_n_364__14_, r_n_364__13_, r_n_364__12_, r_n_364__11_, r_n_364__10_, r_n_364__9_, r_n_364__8_, r_n_364__7_, r_n_364__6_, r_n_364__5_, r_n_364__4_, r_n_364__3_, r_n_364__2_, r_n_364__1_, r_n_364__0_ } = (N728)? { r_365__63_, r_365__62_, r_365__61_, r_365__60_, r_365__59_, r_365__58_, r_365__57_, r_365__56_, r_365__55_, r_365__54_, r_365__53_, r_365__52_, r_365__51_, r_365__50_, r_365__49_, r_365__48_, r_365__47_, r_365__46_, r_365__45_, r_365__44_, r_365__43_, r_365__42_, r_365__41_, r_365__40_, r_365__39_, r_365__38_, r_365__37_, r_365__36_, r_365__35_, r_365__34_, r_365__33_, r_365__32_, r_365__31_, r_365__30_, r_365__29_, r_365__28_, r_365__27_, r_365__26_, r_365__25_, r_365__24_, r_365__23_, r_365__22_, r_365__21_, r_365__20_, r_365__19_, r_365__18_, r_365__17_, r_365__16_, r_365__15_, r_365__14_, r_365__13_, r_365__12_, r_365__11_, r_365__10_, r_365__9_, r_365__8_, r_365__7_, r_365__6_, r_365__5_, r_365__4_, r_365__3_, r_365__2_, r_365__1_, r_365__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N729)? data_i : 1'b0;
  assign N728 = sel_i[728];
  assign N729 = N2848;
  assign { r_n_365__63_, r_n_365__62_, r_n_365__61_, r_n_365__60_, r_n_365__59_, r_n_365__58_, r_n_365__57_, r_n_365__56_, r_n_365__55_, r_n_365__54_, r_n_365__53_, r_n_365__52_, r_n_365__51_, r_n_365__50_, r_n_365__49_, r_n_365__48_, r_n_365__47_, r_n_365__46_, r_n_365__45_, r_n_365__44_, r_n_365__43_, r_n_365__42_, r_n_365__41_, r_n_365__40_, r_n_365__39_, r_n_365__38_, r_n_365__37_, r_n_365__36_, r_n_365__35_, r_n_365__34_, r_n_365__33_, r_n_365__32_, r_n_365__31_, r_n_365__30_, r_n_365__29_, r_n_365__28_, r_n_365__27_, r_n_365__26_, r_n_365__25_, r_n_365__24_, r_n_365__23_, r_n_365__22_, r_n_365__21_, r_n_365__20_, r_n_365__19_, r_n_365__18_, r_n_365__17_, r_n_365__16_, r_n_365__15_, r_n_365__14_, r_n_365__13_, r_n_365__12_, r_n_365__11_, r_n_365__10_, r_n_365__9_, r_n_365__8_, r_n_365__7_, r_n_365__6_, r_n_365__5_, r_n_365__4_, r_n_365__3_, r_n_365__2_, r_n_365__1_, r_n_365__0_ } = (N730)? { r_366__63_, r_366__62_, r_366__61_, r_366__60_, r_366__59_, r_366__58_, r_366__57_, r_366__56_, r_366__55_, r_366__54_, r_366__53_, r_366__52_, r_366__51_, r_366__50_, r_366__49_, r_366__48_, r_366__47_, r_366__46_, r_366__45_, r_366__44_, r_366__43_, r_366__42_, r_366__41_, r_366__40_, r_366__39_, r_366__38_, r_366__37_, r_366__36_, r_366__35_, r_366__34_, r_366__33_, r_366__32_, r_366__31_, r_366__30_, r_366__29_, r_366__28_, r_366__27_, r_366__26_, r_366__25_, r_366__24_, r_366__23_, r_366__22_, r_366__21_, r_366__20_, r_366__19_, r_366__18_, r_366__17_, r_366__16_, r_366__15_, r_366__14_, r_366__13_, r_366__12_, r_366__11_, r_366__10_, r_366__9_, r_366__8_, r_366__7_, r_366__6_, r_366__5_, r_366__4_, r_366__3_, r_366__2_, r_366__1_, r_366__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N731)? data_i : 1'b0;
  assign N730 = sel_i[730];
  assign N731 = N2853;
  assign { r_n_366__63_, r_n_366__62_, r_n_366__61_, r_n_366__60_, r_n_366__59_, r_n_366__58_, r_n_366__57_, r_n_366__56_, r_n_366__55_, r_n_366__54_, r_n_366__53_, r_n_366__52_, r_n_366__51_, r_n_366__50_, r_n_366__49_, r_n_366__48_, r_n_366__47_, r_n_366__46_, r_n_366__45_, r_n_366__44_, r_n_366__43_, r_n_366__42_, r_n_366__41_, r_n_366__40_, r_n_366__39_, r_n_366__38_, r_n_366__37_, r_n_366__36_, r_n_366__35_, r_n_366__34_, r_n_366__33_, r_n_366__32_, r_n_366__31_, r_n_366__30_, r_n_366__29_, r_n_366__28_, r_n_366__27_, r_n_366__26_, r_n_366__25_, r_n_366__24_, r_n_366__23_, r_n_366__22_, r_n_366__21_, r_n_366__20_, r_n_366__19_, r_n_366__18_, r_n_366__17_, r_n_366__16_, r_n_366__15_, r_n_366__14_, r_n_366__13_, r_n_366__12_, r_n_366__11_, r_n_366__10_, r_n_366__9_, r_n_366__8_, r_n_366__7_, r_n_366__6_, r_n_366__5_, r_n_366__4_, r_n_366__3_, r_n_366__2_, r_n_366__1_, r_n_366__0_ } = (N732)? { r_367__63_, r_367__62_, r_367__61_, r_367__60_, r_367__59_, r_367__58_, r_367__57_, r_367__56_, r_367__55_, r_367__54_, r_367__53_, r_367__52_, r_367__51_, r_367__50_, r_367__49_, r_367__48_, r_367__47_, r_367__46_, r_367__45_, r_367__44_, r_367__43_, r_367__42_, r_367__41_, r_367__40_, r_367__39_, r_367__38_, r_367__37_, r_367__36_, r_367__35_, r_367__34_, r_367__33_, r_367__32_, r_367__31_, r_367__30_, r_367__29_, r_367__28_, r_367__27_, r_367__26_, r_367__25_, r_367__24_, r_367__23_, r_367__22_, r_367__21_, r_367__20_, r_367__19_, r_367__18_, r_367__17_, r_367__16_, r_367__15_, r_367__14_, r_367__13_, r_367__12_, r_367__11_, r_367__10_, r_367__9_, r_367__8_, r_367__7_, r_367__6_, r_367__5_, r_367__4_, r_367__3_, r_367__2_, r_367__1_, r_367__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N733)? data_i : 1'b0;
  assign N732 = sel_i[732];
  assign N733 = N2858;
  assign { r_n_367__63_, r_n_367__62_, r_n_367__61_, r_n_367__60_, r_n_367__59_, r_n_367__58_, r_n_367__57_, r_n_367__56_, r_n_367__55_, r_n_367__54_, r_n_367__53_, r_n_367__52_, r_n_367__51_, r_n_367__50_, r_n_367__49_, r_n_367__48_, r_n_367__47_, r_n_367__46_, r_n_367__45_, r_n_367__44_, r_n_367__43_, r_n_367__42_, r_n_367__41_, r_n_367__40_, r_n_367__39_, r_n_367__38_, r_n_367__37_, r_n_367__36_, r_n_367__35_, r_n_367__34_, r_n_367__33_, r_n_367__32_, r_n_367__31_, r_n_367__30_, r_n_367__29_, r_n_367__28_, r_n_367__27_, r_n_367__26_, r_n_367__25_, r_n_367__24_, r_n_367__23_, r_n_367__22_, r_n_367__21_, r_n_367__20_, r_n_367__19_, r_n_367__18_, r_n_367__17_, r_n_367__16_, r_n_367__15_, r_n_367__14_, r_n_367__13_, r_n_367__12_, r_n_367__11_, r_n_367__10_, r_n_367__9_, r_n_367__8_, r_n_367__7_, r_n_367__6_, r_n_367__5_, r_n_367__4_, r_n_367__3_, r_n_367__2_, r_n_367__1_, r_n_367__0_ } = (N734)? { r_368__63_, r_368__62_, r_368__61_, r_368__60_, r_368__59_, r_368__58_, r_368__57_, r_368__56_, r_368__55_, r_368__54_, r_368__53_, r_368__52_, r_368__51_, r_368__50_, r_368__49_, r_368__48_, r_368__47_, r_368__46_, r_368__45_, r_368__44_, r_368__43_, r_368__42_, r_368__41_, r_368__40_, r_368__39_, r_368__38_, r_368__37_, r_368__36_, r_368__35_, r_368__34_, r_368__33_, r_368__32_, r_368__31_, r_368__30_, r_368__29_, r_368__28_, r_368__27_, r_368__26_, r_368__25_, r_368__24_, r_368__23_, r_368__22_, r_368__21_, r_368__20_, r_368__19_, r_368__18_, r_368__17_, r_368__16_, r_368__15_, r_368__14_, r_368__13_, r_368__12_, r_368__11_, r_368__10_, r_368__9_, r_368__8_, r_368__7_, r_368__6_, r_368__5_, r_368__4_, r_368__3_, r_368__2_, r_368__1_, r_368__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N735)? data_i : 1'b0;
  assign N734 = sel_i[734];
  assign N735 = N2863;
  assign { r_n_368__63_, r_n_368__62_, r_n_368__61_, r_n_368__60_, r_n_368__59_, r_n_368__58_, r_n_368__57_, r_n_368__56_, r_n_368__55_, r_n_368__54_, r_n_368__53_, r_n_368__52_, r_n_368__51_, r_n_368__50_, r_n_368__49_, r_n_368__48_, r_n_368__47_, r_n_368__46_, r_n_368__45_, r_n_368__44_, r_n_368__43_, r_n_368__42_, r_n_368__41_, r_n_368__40_, r_n_368__39_, r_n_368__38_, r_n_368__37_, r_n_368__36_, r_n_368__35_, r_n_368__34_, r_n_368__33_, r_n_368__32_, r_n_368__31_, r_n_368__30_, r_n_368__29_, r_n_368__28_, r_n_368__27_, r_n_368__26_, r_n_368__25_, r_n_368__24_, r_n_368__23_, r_n_368__22_, r_n_368__21_, r_n_368__20_, r_n_368__19_, r_n_368__18_, r_n_368__17_, r_n_368__16_, r_n_368__15_, r_n_368__14_, r_n_368__13_, r_n_368__12_, r_n_368__11_, r_n_368__10_, r_n_368__9_, r_n_368__8_, r_n_368__7_, r_n_368__6_, r_n_368__5_, r_n_368__4_, r_n_368__3_, r_n_368__2_, r_n_368__1_, r_n_368__0_ } = (N736)? { r_369__63_, r_369__62_, r_369__61_, r_369__60_, r_369__59_, r_369__58_, r_369__57_, r_369__56_, r_369__55_, r_369__54_, r_369__53_, r_369__52_, r_369__51_, r_369__50_, r_369__49_, r_369__48_, r_369__47_, r_369__46_, r_369__45_, r_369__44_, r_369__43_, r_369__42_, r_369__41_, r_369__40_, r_369__39_, r_369__38_, r_369__37_, r_369__36_, r_369__35_, r_369__34_, r_369__33_, r_369__32_, r_369__31_, r_369__30_, r_369__29_, r_369__28_, r_369__27_, r_369__26_, r_369__25_, r_369__24_, r_369__23_, r_369__22_, r_369__21_, r_369__20_, r_369__19_, r_369__18_, r_369__17_, r_369__16_, r_369__15_, r_369__14_, r_369__13_, r_369__12_, r_369__11_, r_369__10_, r_369__9_, r_369__8_, r_369__7_, r_369__6_, r_369__5_, r_369__4_, r_369__3_, r_369__2_, r_369__1_, r_369__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N737)? data_i : 1'b0;
  assign N736 = sel_i[736];
  assign N737 = N2868;
  assign { r_n_369__63_, r_n_369__62_, r_n_369__61_, r_n_369__60_, r_n_369__59_, r_n_369__58_, r_n_369__57_, r_n_369__56_, r_n_369__55_, r_n_369__54_, r_n_369__53_, r_n_369__52_, r_n_369__51_, r_n_369__50_, r_n_369__49_, r_n_369__48_, r_n_369__47_, r_n_369__46_, r_n_369__45_, r_n_369__44_, r_n_369__43_, r_n_369__42_, r_n_369__41_, r_n_369__40_, r_n_369__39_, r_n_369__38_, r_n_369__37_, r_n_369__36_, r_n_369__35_, r_n_369__34_, r_n_369__33_, r_n_369__32_, r_n_369__31_, r_n_369__30_, r_n_369__29_, r_n_369__28_, r_n_369__27_, r_n_369__26_, r_n_369__25_, r_n_369__24_, r_n_369__23_, r_n_369__22_, r_n_369__21_, r_n_369__20_, r_n_369__19_, r_n_369__18_, r_n_369__17_, r_n_369__16_, r_n_369__15_, r_n_369__14_, r_n_369__13_, r_n_369__12_, r_n_369__11_, r_n_369__10_, r_n_369__9_, r_n_369__8_, r_n_369__7_, r_n_369__6_, r_n_369__5_, r_n_369__4_, r_n_369__3_, r_n_369__2_, r_n_369__1_, r_n_369__0_ } = (N738)? { r_370__63_, r_370__62_, r_370__61_, r_370__60_, r_370__59_, r_370__58_, r_370__57_, r_370__56_, r_370__55_, r_370__54_, r_370__53_, r_370__52_, r_370__51_, r_370__50_, r_370__49_, r_370__48_, r_370__47_, r_370__46_, r_370__45_, r_370__44_, r_370__43_, r_370__42_, r_370__41_, r_370__40_, r_370__39_, r_370__38_, r_370__37_, r_370__36_, r_370__35_, r_370__34_, r_370__33_, r_370__32_, r_370__31_, r_370__30_, r_370__29_, r_370__28_, r_370__27_, r_370__26_, r_370__25_, r_370__24_, r_370__23_, r_370__22_, r_370__21_, r_370__20_, r_370__19_, r_370__18_, r_370__17_, r_370__16_, r_370__15_, r_370__14_, r_370__13_, r_370__12_, r_370__11_, r_370__10_, r_370__9_, r_370__8_, r_370__7_, r_370__6_, r_370__5_, r_370__4_, r_370__3_, r_370__2_, r_370__1_, r_370__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N739)? data_i : 1'b0;
  assign N738 = sel_i[738];
  assign N739 = N2873;
  assign { r_n_370__63_, r_n_370__62_, r_n_370__61_, r_n_370__60_, r_n_370__59_, r_n_370__58_, r_n_370__57_, r_n_370__56_, r_n_370__55_, r_n_370__54_, r_n_370__53_, r_n_370__52_, r_n_370__51_, r_n_370__50_, r_n_370__49_, r_n_370__48_, r_n_370__47_, r_n_370__46_, r_n_370__45_, r_n_370__44_, r_n_370__43_, r_n_370__42_, r_n_370__41_, r_n_370__40_, r_n_370__39_, r_n_370__38_, r_n_370__37_, r_n_370__36_, r_n_370__35_, r_n_370__34_, r_n_370__33_, r_n_370__32_, r_n_370__31_, r_n_370__30_, r_n_370__29_, r_n_370__28_, r_n_370__27_, r_n_370__26_, r_n_370__25_, r_n_370__24_, r_n_370__23_, r_n_370__22_, r_n_370__21_, r_n_370__20_, r_n_370__19_, r_n_370__18_, r_n_370__17_, r_n_370__16_, r_n_370__15_, r_n_370__14_, r_n_370__13_, r_n_370__12_, r_n_370__11_, r_n_370__10_, r_n_370__9_, r_n_370__8_, r_n_370__7_, r_n_370__6_, r_n_370__5_, r_n_370__4_, r_n_370__3_, r_n_370__2_, r_n_370__1_, r_n_370__0_ } = (N740)? { r_371__63_, r_371__62_, r_371__61_, r_371__60_, r_371__59_, r_371__58_, r_371__57_, r_371__56_, r_371__55_, r_371__54_, r_371__53_, r_371__52_, r_371__51_, r_371__50_, r_371__49_, r_371__48_, r_371__47_, r_371__46_, r_371__45_, r_371__44_, r_371__43_, r_371__42_, r_371__41_, r_371__40_, r_371__39_, r_371__38_, r_371__37_, r_371__36_, r_371__35_, r_371__34_, r_371__33_, r_371__32_, r_371__31_, r_371__30_, r_371__29_, r_371__28_, r_371__27_, r_371__26_, r_371__25_, r_371__24_, r_371__23_, r_371__22_, r_371__21_, r_371__20_, r_371__19_, r_371__18_, r_371__17_, r_371__16_, r_371__15_, r_371__14_, r_371__13_, r_371__12_, r_371__11_, r_371__10_, r_371__9_, r_371__8_, r_371__7_, r_371__6_, r_371__5_, r_371__4_, r_371__3_, r_371__2_, r_371__1_, r_371__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N741)? data_i : 1'b0;
  assign N740 = sel_i[740];
  assign N741 = N2878;
  assign { r_n_371__63_, r_n_371__62_, r_n_371__61_, r_n_371__60_, r_n_371__59_, r_n_371__58_, r_n_371__57_, r_n_371__56_, r_n_371__55_, r_n_371__54_, r_n_371__53_, r_n_371__52_, r_n_371__51_, r_n_371__50_, r_n_371__49_, r_n_371__48_, r_n_371__47_, r_n_371__46_, r_n_371__45_, r_n_371__44_, r_n_371__43_, r_n_371__42_, r_n_371__41_, r_n_371__40_, r_n_371__39_, r_n_371__38_, r_n_371__37_, r_n_371__36_, r_n_371__35_, r_n_371__34_, r_n_371__33_, r_n_371__32_, r_n_371__31_, r_n_371__30_, r_n_371__29_, r_n_371__28_, r_n_371__27_, r_n_371__26_, r_n_371__25_, r_n_371__24_, r_n_371__23_, r_n_371__22_, r_n_371__21_, r_n_371__20_, r_n_371__19_, r_n_371__18_, r_n_371__17_, r_n_371__16_, r_n_371__15_, r_n_371__14_, r_n_371__13_, r_n_371__12_, r_n_371__11_, r_n_371__10_, r_n_371__9_, r_n_371__8_, r_n_371__7_, r_n_371__6_, r_n_371__5_, r_n_371__4_, r_n_371__3_, r_n_371__2_, r_n_371__1_, r_n_371__0_ } = (N742)? { r_372__63_, r_372__62_, r_372__61_, r_372__60_, r_372__59_, r_372__58_, r_372__57_, r_372__56_, r_372__55_, r_372__54_, r_372__53_, r_372__52_, r_372__51_, r_372__50_, r_372__49_, r_372__48_, r_372__47_, r_372__46_, r_372__45_, r_372__44_, r_372__43_, r_372__42_, r_372__41_, r_372__40_, r_372__39_, r_372__38_, r_372__37_, r_372__36_, r_372__35_, r_372__34_, r_372__33_, r_372__32_, r_372__31_, r_372__30_, r_372__29_, r_372__28_, r_372__27_, r_372__26_, r_372__25_, r_372__24_, r_372__23_, r_372__22_, r_372__21_, r_372__20_, r_372__19_, r_372__18_, r_372__17_, r_372__16_, r_372__15_, r_372__14_, r_372__13_, r_372__12_, r_372__11_, r_372__10_, r_372__9_, r_372__8_, r_372__7_, r_372__6_, r_372__5_, r_372__4_, r_372__3_, r_372__2_, r_372__1_, r_372__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N743)? data_i : 1'b0;
  assign N742 = sel_i[742];
  assign N743 = N2883;
  assign { r_n_372__63_, r_n_372__62_, r_n_372__61_, r_n_372__60_, r_n_372__59_, r_n_372__58_, r_n_372__57_, r_n_372__56_, r_n_372__55_, r_n_372__54_, r_n_372__53_, r_n_372__52_, r_n_372__51_, r_n_372__50_, r_n_372__49_, r_n_372__48_, r_n_372__47_, r_n_372__46_, r_n_372__45_, r_n_372__44_, r_n_372__43_, r_n_372__42_, r_n_372__41_, r_n_372__40_, r_n_372__39_, r_n_372__38_, r_n_372__37_, r_n_372__36_, r_n_372__35_, r_n_372__34_, r_n_372__33_, r_n_372__32_, r_n_372__31_, r_n_372__30_, r_n_372__29_, r_n_372__28_, r_n_372__27_, r_n_372__26_, r_n_372__25_, r_n_372__24_, r_n_372__23_, r_n_372__22_, r_n_372__21_, r_n_372__20_, r_n_372__19_, r_n_372__18_, r_n_372__17_, r_n_372__16_, r_n_372__15_, r_n_372__14_, r_n_372__13_, r_n_372__12_, r_n_372__11_, r_n_372__10_, r_n_372__9_, r_n_372__8_, r_n_372__7_, r_n_372__6_, r_n_372__5_, r_n_372__4_, r_n_372__3_, r_n_372__2_, r_n_372__1_, r_n_372__0_ } = (N744)? { r_373__63_, r_373__62_, r_373__61_, r_373__60_, r_373__59_, r_373__58_, r_373__57_, r_373__56_, r_373__55_, r_373__54_, r_373__53_, r_373__52_, r_373__51_, r_373__50_, r_373__49_, r_373__48_, r_373__47_, r_373__46_, r_373__45_, r_373__44_, r_373__43_, r_373__42_, r_373__41_, r_373__40_, r_373__39_, r_373__38_, r_373__37_, r_373__36_, r_373__35_, r_373__34_, r_373__33_, r_373__32_, r_373__31_, r_373__30_, r_373__29_, r_373__28_, r_373__27_, r_373__26_, r_373__25_, r_373__24_, r_373__23_, r_373__22_, r_373__21_, r_373__20_, r_373__19_, r_373__18_, r_373__17_, r_373__16_, r_373__15_, r_373__14_, r_373__13_, r_373__12_, r_373__11_, r_373__10_, r_373__9_, r_373__8_, r_373__7_, r_373__6_, r_373__5_, r_373__4_, r_373__3_, r_373__2_, r_373__1_, r_373__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N745)? data_i : 1'b0;
  assign N744 = sel_i[744];
  assign N745 = N2888;
  assign { r_n_373__63_, r_n_373__62_, r_n_373__61_, r_n_373__60_, r_n_373__59_, r_n_373__58_, r_n_373__57_, r_n_373__56_, r_n_373__55_, r_n_373__54_, r_n_373__53_, r_n_373__52_, r_n_373__51_, r_n_373__50_, r_n_373__49_, r_n_373__48_, r_n_373__47_, r_n_373__46_, r_n_373__45_, r_n_373__44_, r_n_373__43_, r_n_373__42_, r_n_373__41_, r_n_373__40_, r_n_373__39_, r_n_373__38_, r_n_373__37_, r_n_373__36_, r_n_373__35_, r_n_373__34_, r_n_373__33_, r_n_373__32_, r_n_373__31_, r_n_373__30_, r_n_373__29_, r_n_373__28_, r_n_373__27_, r_n_373__26_, r_n_373__25_, r_n_373__24_, r_n_373__23_, r_n_373__22_, r_n_373__21_, r_n_373__20_, r_n_373__19_, r_n_373__18_, r_n_373__17_, r_n_373__16_, r_n_373__15_, r_n_373__14_, r_n_373__13_, r_n_373__12_, r_n_373__11_, r_n_373__10_, r_n_373__9_, r_n_373__8_, r_n_373__7_, r_n_373__6_, r_n_373__5_, r_n_373__4_, r_n_373__3_, r_n_373__2_, r_n_373__1_, r_n_373__0_ } = (N746)? { r_374__63_, r_374__62_, r_374__61_, r_374__60_, r_374__59_, r_374__58_, r_374__57_, r_374__56_, r_374__55_, r_374__54_, r_374__53_, r_374__52_, r_374__51_, r_374__50_, r_374__49_, r_374__48_, r_374__47_, r_374__46_, r_374__45_, r_374__44_, r_374__43_, r_374__42_, r_374__41_, r_374__40_, r_374__39_, r_374__38_, r_374__37_, r_374__36_, r_374__35_, r_374__34_, r_374__33_, r_374__32_, r_374__31_, r_374__30_, r_374__29_, r_374__28_, r_374__27_, r_374__26_, r_374__25_, r_374__24_, r_374__23_, r_374__22_, r_374__21_, r_374__20_, r_374__19_, r_374__18_, r_374__17_, r_374__16_, r_374__15_, r_374__14_, r_374__13_, r_374__12_, r_374__11_, r_374__10_, r_374__9_, r_374__8_, r_374__7_, r_374__6_, r_374__5_, r_374__4_, r_374__3_, r_374__2_, r_374__1_, r_374__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N747)? data_i : 1'b0;
  assign N746 = sel_i[746];
  assign N747 = N2893;
  assign { r_n_374__63_, r_n_374__62_, r_n_374__61_, r_n_374__60_, r_n_374__59_, r_n_374__58_, r_n_374__57_, r_n_374__56_, r_n_374__55_, r_n_374__54_, r_n_374__53_, r_n_374__52_, r_n_374__51_, r_n_374__50_, r_n_374__49_, r_n_374__48_, r_n_374__47_, r_n_374__46_, r_n_374__45_, r_n_374__44_, r_n_374__43_, r_n_374__42_, r_n_374__41_, r_n_374__40_, r_n_374__39_, r_n_374__38_, r_n_374__37_, r_n_374__36_, r_n_374__35_, r_n_374__34_, r_n_374__33_, r_n_374__32_, r_n_374__31_, r_n_374__30_, r_n_374__29_, r_n_374__28_, r_n_374__27_, r_n_374__26_, r_n_374__25_, r_n_374__24_, r_n_374__23_, r_n_374__22_, r_n_374__21_, r_n_374__20_, r_n_374__19_, r_n_374__18_, r_n_374__17_, r_n_374__16_, r_n_374__15_, r_n_374__14_, r_n_374__13_, r_n_374__12_, r_n_374__11_, r_n_374__10_, r_n_374__9_, r_n_374__8_, r_n_374__7_, r_n_374__6_, r_n_374__5_, r_n_374__4_, r_n_374__3_, r_n_374__2_, r_n_374__1_, r_n_374__0_ } = (N748)? { r_375__63_, r_375__62_, r_375__61_, r_375__60_, r_375__59_, r_375__58_, r_375__57_, r_375__56_, r_375__55_, r_375__54_, r_375__53_, r_375__52_, r_375__51_, r_375__50_, r_375__49_, r_375__48_, r_375__47_, r_375__46_, r_375__45_, r_375__44_, r_375__43_, r_375__42_, r_375__41_, r_375__40_, r_375__39_, r_375__38_, r_375__37_, r_375__36_, r_375__35_, r_375__34_, r_375__33_, r_375__32_, r_375__31_, r_375__30_, r_375__29_, r_375__28_, r_375__27_, r_375__26_, r_375__25_, r_375__24_, r_375__23_, r_375__22_, r_375__21_, r_375__20_, r_375__19_, r_375__18_, r_375__17_, r_375__16_, r_375__15_, r_375__14_, r_375__13_, r_375__12_, r_375__11_, r_375__10_, r_375__9_, r_375__8_, r_375__7_, r_375__6_, r_375__5_, r_375__4_, r_375__3_, r_375__2_, r_375__1_, r_375__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N749)? data_i : 1'b0;
  assign N748 = sel_i[748];
  assign N749 = N2898;
  assign { r_n_375__63_, r_n_375__62_, r_n_375__61_, r_n_375__60_, r_n_375__59_, r_n_375__58_, r_n_375__57_, r_n_375__56_, r_n_375__55_, r_n_375__54_, r_n_375__53_, r_n_375__52_, r_n_375__51_, r_n_375__50_, r_n_375__49_, r_n_375__48_, r_n_375__47_, r_n_375__46_, r_n_375__45_, r_n_375__44_, r_n_375__43_, r_n_375__42_, r_n_375__41_, r_n_375__40_, r_n_375__39_, r_n_375__38_, r_n_375__37_, r_n_375__36_, r_n_375__35_, r_n_375__34_, r_n_375__33_, r_n_375__32_, r_n_375__31_, r_n_375__30_, r_n_375__29_, r_n_375__28_, r_n_375__27_, r_n_375__26_, r_n_375__25_, r_n_375__24_, r_n_375__23_, r_n_375__22_, r_n_375__21_, r_n_375__20_, r_n_375__19_, r_n_375__18_, r_n_375__17_, r_n_375__16_, r_n_375__15_, r_n_375__14_, r_n_375__13_, r_n_375__12_, r_n_375__11_, r_n_375__10_, r_n_375__9_, r_n_375__8_, r_n_375__7_, r_n_375__6_, r_n_375__5_, r_n_375__4_, r_n_375__3_, r_n_375__2_, r_n_375__1_, r_n_375__0_ } = (N750)? { r_376__63_, r_376__62_, r_376__61_, r_376__60_, r_376__59_, r_376__58_, r_376__57_, r_376__56_, r_376__55_, r_376__54_, r_376__53_, r_376__52_, r_376__51_, r_376__50_, r_376__49_, r_376__48_, r_376__47_, r_376__46_, r_376__45_, r_376__44_, r_376__43_, r_376__42_, r_376__41_, r_376__40_, r_376__39_, r_376__38_, r_376__37_, r_376__36_, r_376__35_, r_376__34_, r_376__33_, r_376__32_, r_376__31_, r_376__30_, r_376__29_, r_376__28_, r_376__27_, r_376__26_, r_376__25_, r_376__24_, r_376__23_, r_376__22_, r_376__21_, r_376__20_, r_376__19_, r_376__18_, r_376__17_, r_376__16_, r_376__15_, r_376__14_, r_376__13_, r_376__12_, r_376__11_, r_376__10_, r_376__9_, r_376__8_, r_376__7_, r_376__6_, r_376__5_, r_376__4_, r_376__3_, r_376__2_, r_376__1_, r_376__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N751)? data_i : 1'b0;
  assign N750 = sel_i[750];
  assign N751 = N2903;
  assign { r_n_376__63_, r_n_376__62_, r_n_376__61_, r_n_376__60_, r_n_376__59_, r_n_376__58_, r_n_376__57_, r_n_376__56_, r_n_376__55_, r_n_376__54_, r_n_376__53_, r_n_376__52_, r_n_376__51_, r_n_376__50_, r_n_376__49_, r_n_376__48_, r_n_376__47_, r_n_376__46_, r_n_376__45_, r_n_376__44_, r_n_376__43_, r_n_376__42_, r_n_376__41_, r_n_376__40_, r_n_376__39_, r_n_376__38_, r_n_376__37_, r_n_376__36_, r_n_376__35_, r_n_376__34_, r_n_376__33_, r_n_376__32_, r_n_376__31_, r_n_376__30_, r_n_376__29_, r_n_376__28_, r_n_376__27_, r_n_376__26_, r_n_376__25_, r_n_376__24_, r_n_376__23_, r_n_376__22_, r_n_376__21_, r_n_376__20_, r_n_376__19_, r_n_376__18_, r_n_376__17_, r_n_376__16_, r_n_376__15_, r_n_376__14_, r_n_376__13_, r_n_376__12_, r_n_376__11_, r_n_376__10_, r_n_376__9_, r_n_376__8_, r_n_376__7_, r_n_376__6_, r_n_376__5_, r_n_376__4_, r_n_376__3_, r_n_376__2_, r_n_376__1_, r_n_376__0_ } = (N752)? { r_377__63_, r_377__62_, r_377__61_, r_377__60_, r_377__59_, r_377__58_, r_377__57_, r_377__56_, r_377__55_, r_377__54_, r_377__53_, r_377__52_, r_377__51_, r_377__50_, r_377__49_, r_377__48_, r_377__47_, r_377__46_, r_377__45_, r_377__44_, r_377__43_, r_377__42_, r_377__41_, r_377__40_, r_377__39_, r_377__38_, r_377__37_, r_377__36_, r_377__35_, r_377__34_, r_377__33_, r_377__32_, r_377__31_, r_377__30_, r_377__29_, r_377__28_, r_377__27_, r_377__26_, r_377__25_, r_377__24_, r_377__23_, r_377__22_, r_377__21_, r_377__20_, r_377__19_, r_377__18_, r_377__17_, r_377__16_, r_377__15_, r_377__14_, r_377__13_, r_377__12_, r_377__11_, r_377__10_, r_377__9_, r_377__8_, r_377__7_, r_377__6_, r_377__5_, r_377__4_, r_377__3_, r_377__2_, r_377__1_, r_377__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N753)? data_i : 1'b0;
  assign N752 = sel_i[752];
  assign N753 = N2908;
  assign { r_n_377__63_, r_n_377__62_, r_n_377__61_, r_n_377__60_, r_n_377__59_, r_n_377__58_, r_n_377__57_, r_n_377__56_, r_n_377__55_, r_n_377__54_, r_n_377__53_, r_n_377__52_, r_n_377__51_, r_n_377__50_, r_n_377__49_, r_n_377__48_, r_n_377__47_, r_n_377__46_, r_n_377__45_, r_n_377__44_, r_n_377__43_, r_n_377__42_, r_n_377__41_, r_n_377__40_, r_n_377__39_, r_n_377__38_, r_n_377__37_, r_n_377__36_, r_n_377__35_, r_n_377__34_, r_n_377__33_, r_n_377__32_, r_n_377__31_, r_n_377__30_, r_n_377__29_, r_n_377__28_, r_n_377__27_, r_n_377__26_, r_n_377__25_, r_n_377__24_, r_n_377__23_, r_n_377__22_, r_n_377__21_, r_n_377__20_, r_n_377__19_, r_n_377__18_, r_n_377__17_, r_n_377__16_, r_n_377__15_, r_n_377__14_, r_n_377__13_, r_n_377__12_, r_n_377__11_, r_n_377__10_, r_n_377__9_, r_n_377__8_, r_n_377__7_, r_n_377__6_, r_n_377__5_, r_n_377__4_, r_n_377__3_, r_n_377__2_, r_n_377__1_, r_n_377__0_ } = (N754)? { r_378__63_, r_378__62_, r_378__61_, r_378__60_, r_378__59_, r_378__58_, r_378__57_, r_378__56_, r_378__55_, r_378__54_, r_378__53_, r_378__52_, r_378__51_, r_378__50_, r_378__49_, r_378__48_, r_378__47_, r_378__46_, r_378__45_, r_378__44_, r_378__43_, r_378__42_, r_378__41_, r_378__40_, r_378__39_, r_378__38_, r_378__37_, r_378__36_, r_378__35_, r_378__34_, r_378__33_, r_378__32_, r_378__31_, r_378__30_, r_378__29_, r_378__28_, r_378__27_, r_378__26_, r_378__25_, r_378__24_, r_378__23_, r_378__22_, r_378__21_, r_378__20_, r_378__19_, r_378__18_, r_378__17_, r_378__16_, r_378__15_, r_378__14_, r_378__13_, r_378__12_, r_378__11_, r_378__10_, r_378__9_, r_378__8_, r_378__7_, r_378__6_, r_378__5_, r_378__4_, r_378__3_, r_378__2_, r_378__1_, r_378__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N755)? data_i : 1'b0;
  assign N754 = sel_i[754];
  assign N755 = N2913;
  assign { r_n_378__63_, r_n_378__62_, r_n_378__61_, r_n_378__60_, r_n_378__59_, r_n_378__58_, r_n_378__57_, r_n_378__56_, r_n_378__55_, r_n_378__54_, r_n_378__53_, r_n_378__52_, r_n_378__51_, r_n_378__50_, r_n_378__49_, r_n_378__48_, r_n_378__47_, r_n_378__46_, r_n_378__45_, r_n_378__44_, r_n_378__43_, r_n_378__42_, r_n_378__41_, r_n_378__40_, r_n_378__39_, r_n_378__38_, r_n_378__37_, r_n_378__36_, r_n_378__35_, r_n_378__34_, r_n_378__33_, r_n_378__32_, r_n_378__31_, r_n_378__30_, r_n_378__29_, r_n_378__28_, r_n_378__27_, r_n_378__26_, r_n_378__25_, r_n_378__24_, r_n_378__23_, r_n_378__22_, r_n_378__21_, r_n_378__20_, r_n_378__19_, r_n_378__18_, r_n_378__17_, r_n_378__16_, r_n_378__15_, r_n_378__14_, r_n_378__13_, r_n_378__12_, r_n_378__11_, r_n_378__10_, r_n_378__9_, r_n_378__8_, r_n_378__7_, r_n_378__6_, r_n_378__5_, r_n_378__4_, r_n_378__3_, r_n_378__2_, r_n_378__1_, r_n_378__0_ } = (N756)? { r_379__63_, r_379__62_, r_379__61_, r_379__60_, r_379__59_, r_379__58_, r_379__57_, r_379__56_, r_379__55_, r_379__54_, r_379__53_, r_379__52_, r_379__51_, r_379__50_, r_379__49_, r_379__48_, r_379__47_, r_379__46_, r_379__45_, r_379__44_, r_379__43_, r_379__42_, r_379__41_, r_379__40_, r_379__39_, r_379__38_, r_379__37_, r_379__36_, r_379__35_, r_379__34_, r_379__33_, r_379__32_, r_379__31_, r_379__30_, r_379__29_, r_379__28_, r_379__27_, r_379__26_, r_379__25_, r_379__24_, r_379__23_, r_379__22_, r_379__21_, r_379__20_, r_379__19_, r_379__18_, r_379__17_, r_379__16_, r_379__15_, r_379__14_, r_379__13_, r_379__12_, r_379__11_, r_379__10_, r_379__9_, r_379__8_, r_379__7_, r_379__6_, r_379__5_, r_379__4_, r_379__3_, r_379__2_, r_379__1_, r_379__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N757)? data_i : 1'b0;
  assign N756 = sel_i[756];
  assign N757 = N2918;
  assign { r_n_379__63_, r_n_379__62_, r_n_379__61_, r_n_379__60_, r_n_379__59_, r_n_379__58_, r_n_379__57_, r_n_379__56_, r_n_379__55_, r_n_379__54_, r_n_379__53_, r_n_379__52_, r_n_379__51_, r_n_379__50_, r_n_379__49_, r_n_379__48_, r_n_379__47_, r_n_379__46_, r_n_379__45_, r_n_379__44_, r_n_379__43_, r_n_379__42_, r_n_379__41_, r_n_379__40_, r_n_379__39_, r_n_379__38_, r_n_379__37_, r_n_379__36_, r_n_379__35_, r_n_379__34_, r_n_379__33_, r_n_379__32_, r_n_379__31_, r_n_379__30_, r_n_379__29_, r_n_379__28_, r_n_379__27_, r_n_379__26_, r_n_379__25_, r_n_379__24_, r_n_379__23_, r_n_379__22_, r_n_379__21_, r_n_379__20_, r_n_379__19_, r_n_379__18_, r_n_379__17_, r_n_379__16_, r_n_379__15_, r_n_379__14_, r_n_379__13_, r_n_379__12_, r_n_379__11_, r_n_379__10_, r_n_379__9_, r_n_379__8_, r_n_379__7_, r_n_379__6_, r_n_379__5_, r_n_379__4_, r_n_379__3_, r_n_379__2_, r_n_379__1_, r_n_379__0_ } = (N758)? { r_380__63_, r_380__62_, r_380__61_, r_380__60_, r_380__59_, r_380__58_, r_380__57_, r_380__56_, r_380__55_, r_380__54_, r_380__53_, r_380__52_, r_380__51_, r_380__50_, r_380__49_, r_380__48_, r_380__47_, r_380__46_, r_380__45_, r_380__44_, r_380__43_, r_380__42_, r_380__41_, r_380__40_, r_380__39_, r_380__38_, r_380__37_, r_380__36_, r_380__35_, r_380__34_, r_380__33_, r_380__32_, r_380__31_, r_380__30_, r_380__29_, r_380__28_, r_380__27_, r_380__26_, r_380__25_, r_380__24_, r_380__23_, r_380__22_, r_380__21_, r_380__20_, r_380__19_, r_380__18_, r_380__17_, r_380__16_, r_380__15_, r_380__14_, r_380__13_, r_380__12_, r_380__11_, r_380__10_, r_380__9_, r_380__8_, r_380__7_, r_380__6_, r_380__5_, r_380__4_, r_380__3_, r_380__2_, r_380__1_, r_380__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N759)? data_i : 1'b0;
  assign N758 = sel_i[758];
  assign N759 = N2923;
  assign { r_n_380__63_, r_n_380__62_, r_n_380__61_, r_n_380__60_, r_n_380__59_, r_n_380__58_, r_n_380__57_, r_n_380__56_, r_n_380__55_, r_n_380__54_, r_n_380__53_, r_n_380__52_, r_n_380__51_, r_n_380__50_, r_n_380__49_, r_n_380__48_, r_n_380__47_, r_n_380__46_, r_n_380__45_, r_n_380__44_, r_n_380__43_, r_n_380__42_, r_n_380__41_, r_n_380__40_, r_n_380__39_, r_n_380__38_, r_n_380__37_, r_n_380__36_, r_n_380__35_, r_n_380__34_, r_n_380__33_, r_n_380__32_, r_n_380__31_, r_n_380__30_, r_n_380__29_, r_n_380__28_, r_n_380__27_, r_n_380__26_, r_n_380__25_, r_n_380__24_, r_n_380__23_, r_n_380__22_, r_n_380__21_, r_n_380__20_, r_n_380__19_, r_n_380__18_, r_n_380__17_, r_n_380__16_, r_n_380__15_, r_n_380__14_, r_n_380__13_, r_n_380__12_, r_n_380__11_, r_n_380__10_, r_n_380__9_, r_n_380__8_, r_n_380__7_, r_n_380__6_, r_n_380__5_, r_n_380__4_, r_n_380__3_, r_n_380__2_, r_n_380__1_, r_n_380__0_ } = (N760)? { r_381__63_, r_381__62_, r_381__61_, r_381__60_, r_381__59_, r_381__58_, r_381__57_, r_381__56_, r_381__55_, r_381__54_, r_381__53_, r_381__52_, r_381__51_, r_381__50_, r_381__49_, r_381__48_, r_381__47_, r_381__46_, r_381__45_, r_381__44_, r_381__43_, r_381__42_, r_381__41_, r_381__40_, r_381__39_, r_381__38_, r_381__37_, r_381__36_, r_381__35_, r_381__34_, r_381__33_, r_381__32_, r_381__31_, r_381__30_, r_381__29_, r_381__28_, r_381__27_, r_381__26_, r_381__25_, r_381__24_, r_381__23_, r_381__22_, r_381__21_, r_381__20_, r_381__19_, r_381__18_, r_381__17_, r_381__16_, r_381__15_, r_381__14_, r_381__13_, r_381__12_, r_381__11_, r_381__10_, r_381__9_, r_381__8_, r_381__7_, r_381__6_, r_381__5_, r_381__4_, r_381__3_, r_381__2_, r_381__1_, r_381__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N761)? data_i : 1'b0;
  assign N760 = sel_i[760];
  assign N761 = N2928;
  assign { r_n_381__63_, r_n_381__62_, r_n_381__61_, r_n_381__60_, r_n_381__59_, r_n_381__58_, r_n_381__57_, r_n_381__56_, r_n_381__55_, r_n_381__54_, r_n_381__53_, r_n_381__52_, r_n_381__51_, r_n_381__50_, r_n_381__49_, r_n_381__48_, r_n_381__47_, r_n_381__46_, r_n_381__45_, r_n_381__44_, r_n_381__43_, r_n_381__42_, r_n_381__41_, r_n_381__40_, r_n_381__39_, r_n_381__38_, r_n_381__37_, r_n_381__36_, r_n_381__35_, r_n_381__34_, r_n_381__33_, r_n_381__32_, r_n_381__31_, r_n_381__30_, r_n_381__29_, r_n_381__28_, r_n_381__27_, r_n_381__26_, r_n_381__25_, r_n_381__24_, r_n_381__23_, r_n_381__22_, r_n_381__21_, r_n_381__20_, r_n_381__19_, r_n_381__18_, r_n_381__17_, r_n_381__16_, r_n_381__15_, r_n_381__14_, r_n_381__13_, r_n_381__12_, r_n_381__11_, r_n_381__10_, r_n_381__9_, r_n_381__8_, r_n_381__7_, r_n_381__6_, r_n_381__5_, r_n_381__4_, r_n_381__3_, r_n_381__2_, r_n_381__1_, r_n_381__0_ } = (N762)? { r_382__63_, r_382__62_, r_382__61_, r_382__60_, r_382__59_, r_382__58_, r_382__57_, r_382__56_, r_382__55_, r_382__54_, r_382__53_, r_382__52_, r_382__51_, r_382__50_, r_382__49_, r_382__48_, r_382__47_, r_382__46_, r_382__45_, r_382__44_, r_382__43_, r_382__42_, r_382__41_, r_382__40_, r_382__39_, r_382__38_, r_382__37_, r_382__36_, r_382__35_, r_382__34_, r_382__33_, r_382__32_, r_382__31_, r_382__30_, r_382__29_, r_382__28_, r_382__27_, r_382__26_, r_382__25_, r_382__24_, r_382__23_, r_382__22_, r_382__21_, r_382__20_, r_382__19_, r_382__18_, r_382__17_, r_382__16_, r_382__15_, r_382__14_, r_382__13_, r_382__12_, r_382__11_, r_382__10_, r_382__9_, r_382__8_, r_382__7_, r_382__6_, r_382__5_, r_382__4_, r_382__3_, r_382__2_, r_382__1_, r_382__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N763)? data_i : 1'b0;
  assign N762 = sel_i[762];
  assign N763 = N2933;
  assign { r_n_382__63_, r_n_382__62_, r_n_382__61_, r_n_382__60_, r_n_382__59_, r_n_382__58_, r_n_382__57_, r_n_382__56_, r_n_382__55_, r_n_382__54_, r_n_382__53_, r_n_382__52_, r_n_382__51_, r_n_382__50_, r_n_382__49_, r_n_382__48_, r_n_382__47_, r_n_382__46_, r_n_382__45_, r_n_382__44_, r_n_382__43_, r_n_382__42_, r_n_382__41_, r_n_382__40_, r_n_382__39_, r_n_382__38_, r_n_382__37_, r_n_382__36_, r_n_382__35_, r_n_382__34_, r_n_382__33_, r_n_382__32_, r_n_382__31_, r_n_382__30_, r_n_382__29_, r_n_382__28_, r_n_382__27_, r_n_382__26_, r_n_382__25_, r_n_382__24_, r_n_382__23_, r_n_382__22_, r_n_382__21_, r_n_382__20_, r_n_382__19_, r_n_382__18_, r_n_382__17_, r_n_382__16_, r_n_382__15_, r_n_382__14_, r_n_382__13_, r_n_382__12_, r_n_382__11_, r_n_382__10_, r_n_382__9_, r_n_382__8_, r_n_382__7_, r_n_382__6_, r_n_382__5_, r_n_382__4_, r_n_382__3_, r_n_382__2_, r_n_382__1_, r_n_382__0_ } = (N764)? { r_383__63_, r_383__62_, r_383__61_, r_383__60_, r_383__59_, r_383__58_, r_383__57_, r_383__56_, r_383__55_, r_383__54_, r_383__53_, r_383__52_, r_383__51_, r_383__50_, r_383__49_, r_383__48_, r_383__47_, r_383__46_, r_383__45_, r_383__44_, r_383__43_, r_383__42_, r_383__41_, r_383__40_, r_383__39_, r_383__38_, r_383__37_, r_383__36_, r_383__35_, r_383__34_, r_383__33_, r_383__32_, r_383__31_, r_383__30_, r_383__29_, r_383__28_, r_383__27_, r_383__26_, r_383__25_, r_383__24_, r_383__23_, r_383__22_, r_383__21_, r_383__20_, r_383__19_, r_383__18_, r_383__17_, r_383__16_, r_383__15_, r_383__14_, r_383__13_, r_383__12_, r_383__11_, r_383__10_, r_383__9_, r_383__8_, r_383__7_, r_383__6_, r_383__5_, r_383__4_, r_383__3_, r_383__2_, r_383__1_, r_383__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N765)? data_i : 1'b0;
  assign N764 = sel_i[764];
  assign N765 = N2938;
  assign { r_n_383__63_, r_n_383__62_, r_n_383__61_, r_n_383__60_, r_n_383__59_, r_n_383__58_, r_n_383__57_, r_n_383__56_, r_n_383__55_, r_n_383__54_, r_n_383__53_, r_n_383__52_, r_n_383__51_, r_n_383__50_, r_n_383__49_, r_n_383__48_, r_n_383__47_, r_n_383__46_, r_n_383__45_, r_n_383__44_, r_n_383__43_, r_n_383__42_, r_n_383__41_, r_n_383__40_, r_n_383__39_, r_n_383__38_, r_n_383__37_, r_n_383__36_, r_n_383__35_, r_n_383__34_, r_n_383__33_, r_n_383__32_, r_n_383__31_, r_n_383__30_, r_n_383__29_, r_n_383__28_, r_n_383__27_, r_n_383__26_, r_n_383__25_, r_n_383__24_, r_n_383__23_, r_n_383__22_, r_n_383__21_, r_n_383__20_, r_n_383__19_, r_n_383__18_, r_n_383__17_, r_n_383__16_, r_n_383__15_, r_n_383__14_, r_n_383__13_, r_n_383__12_, r_n_383__11_, r_n_383__10_, r_n_383__9_, r_n_383__8_, r_n_383__7_, r_n_383__6_, r_n_383__5_, r_n_383__4_, r_n_383__3_, r_n_383__2_, r_n_383__1_, r_n_383__0_ } = (N766)? { r_384__63_, r_384__62_, r_384__61_, r_384__60_, r_384__59_, r_384__58_, r_384__57_, r_384__56_, r_384__55_, r_384__54_, r_384__53_, r_384__52_, r_384__51_, r_384__50_, r_384__49_, r_384__48_, r_384__47_, r_384__46_, r_384__45_, r_384__44_, r_384__43_, r_384__42_, r_384__41_, r_384__40_, r_384__39_, r_384__38_, r_384__37_, r_384__36_, r_384__35_, r_384__34_, r_384__33_, r_384__32_, r_384__31_, r_384__30_, r_384__29_, r_384__28_, r_384__27_, r_384__26_, r_384__25_, r_384__24_, r_384__23_, r_384__22_, r_384__21_, r_384__20_, r_384__19_, r_384__18_, r_384__17_, r_384__16_, r_384__15_, r_384__14_, r_384__13_, r_384__12_, r_384__11_, r_384__10_, r_384__9_, r_384__8_, r_384__7_, r_384__6_, r_384__5_, r_384__4_, r_384__3_, r_384__2_, r_384__1_, r_384__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N767)? data_i : 1'b0;
  assign N766 = sel_i[766];
  assign N767 = N2943;
  assign { r_n_384__63_, r_n_384__62_, r_n_384__61_, r_n_384__60_, r_n_384__59_, r_n_384__58_, r_n_384__57_, r_n_384__56_, r_n_384__55_, r_n_384__54_, r_n_384__53_, r_n_384__52_, r_n_384__51_, r_n_384__50_, r_n_384__49_, r_n_384__48_, r_n_384__47_, r_n_384__46_, r_n_384__45_, r_n_384__44_, r_n_384__43_, r_n_384__42_, r_n_384__41_, r_n_384__40_, r_n_384__39_, r_n_384__38_, r_n_384__37_, r_n_384__36_, r_n_384__35_, r_n_384__34_, r_n_384__33_, r_n_384__32_, r_n_384__31_, r_n_384__30_, r_n_384__29_, r_n_384__28_, r_n_384__27_, r_n_384__26_, r_n_384__25_, r_n_384__24_, r_n_384__23_, r_n_384__22_, r_n_384__21_, r_n_384__20_, r_n_384__19_, r_n_384__18_, r_n_384__17_, r_n_384__16_, r_n_384__15_, r_n_384__14_, r_n_384__13_, r_n_384__12_, r_n_384__11_, r_n_384__10_, r_n_384__9_, r_n_384__8_, r_n_384__7_, r_n_384__6_, r_n_384__5_, r_n_384__4_, r_n_384__3_, r_n_384__2_, r_n_384__1_, r_n_384__0_ } = (N768)? { r_385__63_, r_385__62_, r_385__61_, r_385__60_, r_385__59_, r_385__58_, r_385__57_, r_385__56_, r_385__55_, r_385__54_, r_385__53_, r_385__52_, r_385__51_, r_385__50_, r_385__49_, r_385__48_, r_385__47_, r_385__46_, r_385__45_, r_385__44_, r_385__43_, r_385__42_, r_385__41_, r_385__40_, r_385__39_, r_385__38_, r_385__37_, r_385__36_, r_385__35_, r_385__34_, r_385__33_, r_385__32_, r_385__31_, r_385__30_, r_385__29_, r_385__28_, r_385__27_, r_385__26_, r_385__25_, r_385__24_, r_385__23_, r_385__22_, r_385__21_, r_385__20_, r_385__19_, r_385__18_, r_385__17_, r_385__16_, r_385__15_, r_385__14_, r_385__13_, r_385__12_, r_385__11_, r_385__10_, r_385__9_, r_385__8_, r_385__7_, r_385__6_, r_385__5_, r_385__4_, r_385__3_, r_385__2_, r_385__1_, r_385__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N769)? data_i : 1'b0;
  assign N768 = sel_i[768];
  assign N769 = N2948;
  assign { r_n_385__63_, r_n_385__62_, r_n_385__61_, r_n_385__60_, r_n_385__59_, r_n_385__58_, r_n_385__57_, r_n_385__56_, r_n_385__55_, r_n_385__54_, r_n_385__53_, r_n_385__52_, r_n_385__51_, r_n_385__50_, r_n_385__49_, r_n_385__48_, r_n_385__47_, r_n_385__46_, r_n_385__45_, r_n_385__44_, r_n_385__43_, r_n_385__42_, r_n_385__41_, r_n_385__40_, r_n_385__39_, r_n_385__38_, r_n_385__37_, r_n_385__36_, r_n_385__35_, r_n_385__34_, r_n_385__33_, r_n_385__32_, r_n_385__31_, r_n_385__30_, r_n_385__29_, r_n_385__28_, r_n_385__27_, r_n_385__26_, r_n_385__25_, r_n_385__24_, r_n_385__23_, r_n_385__22_, r_n_385__21_, r_n_385__20_, r_n_385__19_, r_n_385__18_, r_n_385__17_, r_n_385__16_, r_n_385__15_, r_n_385__14_, r_n_385__13_, r_n_385__12_, r_n_385__11_, r_n_385__10_, r_n_385__9_, r_n_385__8_, r_n_385__7_, r_n_385__6_, r_n_385__5_, r_n_385__4_, r_n_385__3_, r_n_385__2_, r_n_385__1_, r_n_385__0_ } = (N770)? { r_386__63_, r_386__62_, r_386__61_, r_386__60_, r_386__59_, r_386__58_, r_386__57_, r_386__56_, r_386__55_, r_386__54_, r_386__53_, r_386__52_, r_386__51_, r_386__50_, r_386__49_, r_386__48_, r_386__47_, r_386__46_, r_386__45_, r_386__44_, r_386__43_, r_386__42_, r_386__41_, r_386__40_, r_386__39_, r_386__38_, r_386__37_, r_386__36_, r_386__35_, r_386__34_, r_386__33_, r_386__32_, r_386__31_, r_386__30_, r_386__29_, r_386__28_, r_386__27_, r_386__26_, r_386__25_, r_386__24_, r_386__23_, r_386__22_, r_386__21_, r_386__20_, r_386__19_, r_386__18_, r_386__17_, r_386__16_, r_386__15_, r_386__14_, r_386__13_, r_386__12_, r_386__11_, r_386__10_, r_386__9_, r_386__8_, r_386__7_, r_386__6_, r_386__5_, r_386__4_, r_386__3_, r_386__2_, r_386__1_, r_386__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N771)? data_i : 1'b0;
  assign N770 = sel_i[770];
  assign N771 = N2953;
  assign { r_n_386__63_, r_n_386__62_, r_n_386__61_, r_n_386__60_, r_n_386__59_, r_n_386__58_, r_n_386__57_, r_n_386__56_, r_n_386__55_, r_n_386__54_, r_n_386__53_, r_n_386__52_, r_n_386__51_, r_n_386__50_, r_n_386__49_, r_n_386__48_, r_n_386__47_, r_n_386__46_, r_n_386__45_, r_n_386__44_, r_n_386__43_, r_n_386__42_, r_n_386__41_, r_n_386__40_, r_n_386__39_, r_n_386__38_, r_n_386__37_, r_n_386__36_, r_n_386__35_, r_n_386__34_, r_n_386__33_, r_n_386__32_, r_n_386__31_, r_n_386__30_, r_n_386__29_, r_n_386__28_, r_n_386__27_, r_n_386__26_, r_n_386__25_, r_n_386__24_, r_n_386__23_, r_n_386__22_, r_n_386__21_, r_n_386__20_, r_n_386__19_, r_n_386__18_, r_n_386__17_, r_n_386__16_, r_n_386__15_, r_n_386__14_, r_n_386__13_, r_n_386__12_, r_n_386__11_, r_n_386__10_, r_n_386__9_, r_n_386__8_, r_n_386__7_, r_n_386__6_, r_n_386__5_, r_n_386__4_, r_n_386__3_, r_n_386__2_, r_n_386__1_, r_n_386__0_ } = (N772)? { r_387__63_, r_387__62_, r_387__61_, r_387__60_, r_387__59_, r_387__58_, r_387__57_, r_387__56_, r_387__55_, r_387__54_, r_387__53_, r_387__52_, r_387__51_, r_387__50_, r_387__49_, r_387__48_, r_387__47_, r_387__46_, r_387__45_, r_387__44_, r_387__43_, r_387__42_, r_387__41_, r_387__40_, r_387__39_, r_387__38_, r_387__37_, r_387__36_, r_387__35_, r_387__34_, r_387__33_, r_387__32_, r_387__31_, r_387__30_, r_387__29_, r_387__28_, r_387__27_, r_387__26_, r_387__25_, r_387__24_, r_387__23_, r_387__22_, r_387__21_, r_387__20_, r_387__19_, r_387__18_, r_387__17_, r_387__16_, r_387__15_, r_387__14_, r_387__13_, r_387__12_, r_387__11_, r_387__10_, r_387__9_, r_387__8_, r_387__7_, r_387__6_, r_387__5_, r_387__4_, r_387__3_, r_387__2_, r_387__1_, r_387__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N773)? data_i : 1'b0;
  assign N772 = sel_i[772];
  assign N773 = N2958;
  assign { r_n_387__63_, r_n_387__62_, r_n_387__61_, r_n_387__60_, r_n_387__59_, r_n_387__58_, r_n_387__57_, r_n_387__56_, r_n_387__55_, r_n_387__54_, r_n_387__53_, r_n_387__52_, r_n_387__51_, r_n_387__50_, r_n_387__49_, r_n_387__48_, r_n_387__47_, r_n_387__46_, r_n_387__45_, r_n_387__44_, r_n_387__43_, r_n_387__42_, r_n_387__41_, r_n_387__40_, r_n_387__39_, r_n_387__38_, r_n_387__37_, r_n_387__36_, r_n_387__35_, r_n_387__34_, r_n_387__33_, r_n_387__32_, r_n_387__31_, r_n_387__30_, r_n_387__29_, r_n_387__28_, r_n_387__27_, r_n_387__26_, r_n_387__25_, r_n_387__24_, r_n_387__23_, r_n_387__22_, r_n_387__21_, r_n_387__20_, r_n_387__19_, r_n_387__18_, r_n_387__17_, r_n_387__16_, r_n_387__15_, r_n_387__14_, r_n_387__13_, r_n_387__12_, r_n_387__11_, r_n_387__10_, r_n_387__9_, r_n_387__8_, r_n_387__7_, r_n_387__6_, r_n_387__5_, r_n_387__4_, r_n_387__3_, r_n_387__2_, r_n_387__1_, r_n_387__0_ } = (N774)? { r_388__63_, r_388__62_, r_388__61_, r_388__60_, r_388__59_, r_388__58_, r_388__57_, r_388__56_, r_388__55_, r_388__54_, r_388__53_, r_388__52_, r_388__51_, r_388__50_, r_388__49_, r_388__48_, r_388__47_, r_388__46_, r_388__45_, r_388__44_, r_388__43_, r_388__42_, r_388__41_, r_388__40_, r_388__39_, r_388__38_, r_388__37_, r_388__36_, r_388__35_, r_388__34_, r_388__33_, r_388__32_, r_388__31_, r_388__30_, r_388__29_, r_388__28_, r_388__27_, r_388__26_, r_388__25_, r_388__24_, r_388__23_, r_388__22_, r_388__21_, r_388__20_, r_388__19_, r_388__18_, r_388__17_, r_388__16_, r_388__15_, r_388__14_, r_388__13_, r_388__12_, r_388__11_, r_388__10_, r_388__9_, r_388__8_, r_388__7_, r_388__6_, r_388__5_, r_388__4_, r_388__3_, r_388__2_, r_388__1_, r_388__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N775)? data_i : 1'b0;
  assign N774 = sel_i[774];
  assign N775 = N2963;
  assign { r_n_388__63_, r_n_388__62_, r_n_388__61_, r_n_388__60_, r_n_388__59_, r_n_388__58_, r_n_388__57_, r_n_388__56_, r_n_388__55_, r_n_388__54_, r_n_388__53_, r_n_388__52_, r_n_388__51_, r_n_388__50_, r_n_388__49_, r_n_388__48_, r_n_388__47_, r_n_388__46_, r_n_388__45_, r_n_388__44_, r_n_388__43_, r_n_388__42_, r_n_388__41_, r_n_388__40_, r_n_388__39_, r_n_388__38_, r_n_388__37_, r_n_388__36_, r_n_388__35_, r_n_388__34_, r_n_388__33_, r_n_388__32_, r_n_388__31_, r_n_388__30_, r_n_388__29_, r_n_388__28_, r_n_388__27_, r_n_388__26_, r_n_388__25_, r_n_388__24_, r_n_388__23_, r_n_388__22_, r_n_388__21_, r_n_388__20_, r_n_388__19_, r_n_388__18_, r_n_388__17_, r_n_388__16_, r_n_388__15_, r_n_388__14_, r_n_388__13_, r_n_388__12_, r_n_388__11_, r_n_388__10_, r_n_388__9_, r_n_388__8_, r_n_388__7_, r_n_388__6_, r_n_388__5_, r_n_388__4_, r_n_388__3_, r_n_388__2_, r_n_388__1_, r_n_388__0_ } = (N776)? { r_389__63_, r_389__62_, r_389__61_, r_389__60_, r_389__59_, r_389__58_, r_389__57_, r_389__56_, r_389__55_, r_389__54_, r_389__53_, r_389__52_, r_389__51_, r_389__50_, r_389__49_, r_389__48_, r_389__47_, r_389__46_, r_389__45_, r_389__44_, r_389__43_, r_389__42_, r_389__41_, r_389__40_, r_389__39_, r_389__38_, r_389__37_, r_389__36_, r_389__35_, r_389__34_, r_389__33_, r_389__32_, r_389__31_, r_389__30_, r_389__29_, r_389__28_, r_389__27_, r_389__26_, r_389__25_, r_389__24_, r_389__23_, r_389__22_, r_389__21_, r_389__20_, r_389__19_, r_389__18_, r_389__17_, r_389__16_, r_389__15_, r_389__14_, r_389__13_, r_389__12_, r_389__11_, r_389__10_, r_389__9_, r_389__8_, r_389__7_, r_389__6_, r_389__5_, r_389__4_, r_389__3_, r_389__2_, r_389__1_, r_389__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N777)? data_i : 1'b0;
  assign N776 = sel_i[776];
  assign N777 = N2968;
  assign { r_n_389__63_, r_n_389__62_, r_n_389__61_, r_n_389__60_, r_n_389__59_, r_n_389__58_, r_n_389__57_, r_n_389__56_, r_n_389__55_, r_n_389__54_, r_n_389__53_, r_n_389__52_, r_n_389__51_, r_n_389__50_, r_n_389__49_, r_n_389__48_, r_n_389__47_, r_n_389__46_, r_n_389__45_, r_n_389__44_, r_n_389__43_, r_n_389__42_, r_n_389__41_, r_n_389__40_, r_n_389__39_, r_n_389__38_, r_n_389__37_, r_n_389__36_, r_n_389__35_, r_n_389__34_, r_n_389__33_, r_n_389__32_, r_n_389__31_, r_n_389__30_, r_n_389__29_, r_n_389__28_, r_n_389__27_, r_n_389__26_, r_n_389__25_, r_n_389__24_, r_n_389__23_, r_n_389__22_, r_n_389__21_, r_n_389__20_, r_n_389__19_, r_n_389__18_, r_n_389__17_, r_n_389__16_, r_n_389__15_, r_n_389__14_, r_n_389__13_, r_n_389__12_, r_n_389__11_, r_n_389__10_, r_n_389__9_, r_n_389__8_, r_n_389__7_, r_n_389__6_, r_n_389__5_, r_n_389__4_, r_n_389__3_, r_n_389__2_, r_n_389__1_, r_n_389__0_ } = (N778)? { r_390__63_, r_390__62_, r_390__61_, r_390__60_, r_390__59_, r_390__58_, r_390__57_, r_390__56_, r_390__55_, r_390__54_, r_390__53_, r_390__52_, r_390__51_, r_390__50_, r_390__49_, r_390__48_, r_390__47_, r_390__46_, r_390__45_, r_390__44_, r_390__43_, r_390__42_, r_390__41_, r_390__40_, r_390__39_, r_390__38_, r_390__37_, r_390__36_, r_390__35_, r_390__34_, r_390__33_, r_390__32_, r_390__31_, r_390__30_, r_390__29_, r_390__28_, r_390__27_, r_390__26_, r_390__25_, r_390__24_, r_390__23_, r_390__22_, r_390__21_, r_390__20_, r_390__19_, r_390__18_, r_390__17_, r_390__16_, r_390__15_, r_390__14_, r_390__13_, r_390__12_, r_390__11_, r_390__10_, r_390__9_, r_390__8_, r_390__7_, r_390__6_, r_390__5_, r_390__4_, r_390__3_, r_390__2_, r_390__1_, r_390__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N779)? data_i : 1'b0;
  assign N778 = sel_i[778];
  assign N779 = N2973;
  assign { r_n_390__63_, r_n_390__62_, r_n_390__61_, r_n_390__60_, r_n_390__59_, r_n_390__58_, r_n_390__57_, r_n_390__56_, r_n_390__55_, r_n_390__54_, r_n_390__53_, r_n_390__52_, r_n_390__51_, r_n_390__50_, r_n_390__49_, r_n_390__48_, r_n_390__47_, r_n_390__46_, r_n_390__45_, r_n_390__44_, r_n_390__43_, r_n_390__42_, r_n_390__41_, r_n_390__40_, r_n_390__39_, r_n_390__38_, r_n_390__37_, r_n_390__36_, r_n_390__35_, r_n_390__34_, r_n_390__33_, r_n_390__32_, r_n_390__31_, r_n_390__30_, r_n_390__29_, r_n_390__28_, r_n_390__27_, r_n_390__26_, r_n_390__25_, r_n_390__24_, r_n_390__23_, r_n_390__22_, r_n_390__21_, r_n_390__20_, r_n_390__19_, r_n_390__18_, r_n_390__17_, r_n_390__16_, r_n_390__15_, r_n_390__14_, r_n_390__13_, r_n_390__12_, r_n_390__11_, r_n_390__10_, r_n_390__9_, r_n_390__8_, r_n_390__7_, r_n_390__6_, r_n_390__5_, r_n_390__4_, r_n_390__3_, r_n_390__2_, r_n_390__1_, r_n_390__0_ } = (N780)? { r_391__63_, r_391__62_, r_391__61_, r_391__60_, r_391__59_, r_391__58_, r_391__57_, r_391__56_, r_391__55_, r_391__54_, r_391__53_, r_391__52_, r_391__51_, r_391__50_, r_391__49_, r_391__48_, r_391__47_, r_391__46_, r_391__45_, r_391__44_, r_391__43_, r_391__42_, r_391__41_, r_391__40_, r_391__39_, r_391__38_, r_391__37_, r_391__36_, r_391__35_, r_391__34_, r_391__33_, r_391__32_, r_391__31_, r_391__30_, r_391__29_, r_391__28_, r_391__27_, r_391__26_, r_391__25_, r_391__24_, r_391__23_, r_391__22_, r_391__21_, r_391__20_, r_391__19_, r_391__18_, r_391__17_, r_391__16_, r_391__15_, r_391__14_, r_391__13_, r_391__12_, r_391__11_, r_391__10_, r_391__9_, r_391__8_, r_391__7_, r_391__6_, r_391__5_, r_391__4_, r_391__3_, r_391__2_, r_391__1_, r_391__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N781)? data_i : 1'b0;
  assign N780 = sel_i[780];
  assign N781 = N2978;
  assign { r_n_391__63_, r_n_391__62_, r_n_391__61_, r_n_391__60_, r_n_391__59_, r_n_391__58_, r_n_391__57_, r_n_391__56_, r_n_391__55_, r_n_391__54_, r_n_391__53_, r_n_391__52_, r_n_391__51_, r_n_391__50_, r_n_391__49_, r_n_391__48_, r_n_391__47_, r_n_391__46_, r_n_391__45_, r_n_391__44_, r_n_391__43_, r_n_391__42_, r_n_391__41_, r_n_391__40_, r_n_391__39_, r_n_391__38_, r_n_391__37_, r_n_391__36_, r_n_391__35_, r_n_391__34_, r_n_391__33_, r_n_391__32_, r_n_391__31_, r_n_391__30_, r_n_391__29_, r_n_391__28_, r_n_391__27_, r_n_391__26_, r_n_391__25_, r_n_391__24_, r_n_391__23_, r_n_391__22_, r_n_391__21_, r_n_391__20_, r_n_391__19_, r_n_391__18_, r_n_391__17_, r_n_391__16_, r_n_391__15_, r_n_391__14_, r_n_391__13_, r_n_391__12_, r_n_391__11_, r_n_391__10_, r_n_391__9_, r_n_391__8_, r_n_391__7_, r_n_391__6_, r_n_391__5_, r_n_391__4_, r_n_391__3_, r_n_391__2_, r_n_391__1_, r_n_391__0_ } = (N782)? { r_392__63_, r_392__62_, r_392__61_, r_392__60_, r_392__59_, r_392__58_, r_392__57_, r_392__56_, r_392__55_, r_392__54_, r_392__53_, r_392__52_, r_392__51_, r_392__50_, r_392__49_, r_392__48_, r_392__47_, r_392__46_, r_392__45_, r_392__44_, r_392__43_, r_392__42_, r_392__41_, r_392__40_, r_392__39_, r_392__38_, r_392__37_, r_392__36_, r_392__35_, r_392__34_, r_392__33_, r_392__32_, r_392__31_, r_392__30_, r_392__29_, r_392__28_, r_392__27_, r_392__26_, r_392__25_, r_392__24_, r_392__23_, r_392__22_, r_392__21_, r_392__20_, r_392__19_, r_392__18_, r_392__17_, r_392__16_, r_392__15_, r_392__14_, r_392__13_, r_392__12_, r_392__11_, r_392__10_, r_392__9_, r_392__8_, r_392__7_, r_392__6_, r_392__5_, r_392__4_, r_392__3_, r_392__2_, r_392__1_, r_392__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N783)? data_i : 1'b0;
  assign N782 = sel_i[782];
  assign N783 = N2983;
  assign { r_n_392__63_, r_n_392__62_, r_n_392__61_, r_n_392__60_, r_n_392__59_, r_n_392__58_, r_n_392__57_, r_n_392__56_, r_n_392__55_, r_n_392__54_, r_n_392__53_, r_n_392__52_, r_n_392__51_, r_n_392__50_, r_n_392__49_, r_n_392__48_, r_n_392__47_, r_n_392__46_, r_n_392__45_, r_n_392__44_, r_n_392__43_, r_n_392__42_, r_n_392__41_, r_n_392__40_, r_n_392__39_, r_n_392__38_, r_n_392__37_, r_n_392__36_, r_n_392__35_, r_n_392__34_, r_n_392__33_, r_n_392__32_, r_n_392__31_, r_n_392__30_, r_n_392__29_, r_n_392__28_, r_n_392__27_, r_n_392__26_, r_n_392__25_, r_n_392__24_, r_n_392__23_, r_n_392__22_, r_n_392__21_, r_n_392__20_, r_n_392__19_, r_n_392__18_, r_n_392__17_, r_n_392__16_, r_n_392__15_, r_n_392__14_, r_n_392__13_, r_n_392__12_, r_n_392__11_, r_n_392__10_, r_n_392__9_, r_n_392__8_, r_n_392__7_, r_n_392__6_, r_n_392__5_, r_n_392__4_, r_n_392__3_, r_n_392__2_, r_n_392__1_, r_n_392__0_ } = (N784)? { r_393__63_, r_393__62_, r_393__61_, r_393__60_, r_393__59_, r_393__58_, r_393__57_, r_393__56_, r_393__55_, r_393__54_, r_393__53_, r_393__52_, r_393__51_, r_393__50_, r_393__49_, r_393__48_, r_393__47_, r_393__46_, r_393__45_, r_393__44_, r_393__43_, r_393__42_, r_393__41_, r_393__40_, r_393__39_, r_393__38_, r_393__37_, r_393__36_, r_393__35_, r_393__34_, r_393__33_, r_393__32_, r_393__31_, r_393__30_, r_393__29_, r_393__28_, r_393__27_, r_393__26_, r_393__25_, r_393__24_, r_393__23_, r_393__22_, r_393__21_, r_393__20_, r_393__19_, r_393__18_, r_393__17_, r_393__16_, r_393__15_, r_393__14_, r_393__13_, r_393__12_, r_393__11_, r_393__10_, r_393__9_, r_393__8_, r_393__7_, r_393__6_, r_393__5_, r_393__4_, r_393__3_, r_393__2_, r_393__1_, r_393__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N785)? data_i : 1'b0;
  assign N784 = sel_i[784];
  assign N785 = N2988;
  assign { r_n_393__63_, r_n_393__62_, r_n_393__61_, r_n_393__60_, r_n_393__59_, r_n_393__58_, r_n_393__57_, r_n_393__56_, r_n_393__55_, r_n_393__54_, r_n_393__53_, r_n_393__52_, r_n_393__51_, r_n_393__50_, r_n_393__49_, r_n_393__48_, r_n_393__47_, r_n_393__46_, r_n_393__45_, r_n_393__44_, r_n_393__43_, r_n_393__42_, r_n_393__41_, r_n_393__40_, r_n_393__39_, r_n_393__38_, r_n_393__37_, r_n_393__36_, r_n_393__35_, r_n_393__34_, r_n_393__33_, r_n_393__32_, r_n_393__31_, r_n_393__30_, r_n_393__29_, r_n_393__28_, r_n_393__27_, r_n_393__26_, r_n_393__25_, r_n_393__24_, r_n_393__23_, r_n_393__22_, r_n_393__21_, r_n_393__20_, r_n_393__19_, r_n_393__18_, r_n_393__17_, r_n_393__16_, r_n_393__15_, r_n_393__14_, r_n_393__13_, r_n_393__12_, r_n_393__11_, r_n_393__10_, r_n_393__9_, r_n_393__8_, r_n_393__7_, r_n_393__6_, r_n_393__5_, r_n_393__4_, r_n_393__3_, r_n_393__2_, r_n_393__1_, r_n_393__0_ } = (N786)? { r_394__63_, r_394__62_, r_394__61_, r_394__60_, r_394__59_, r_394__58_, r_394__57_, r_394__56_, r_394__55_, r_394__54_, r_394__53_, r_394__52_, r_394__51_, r_394__50_, r_394__49_, r_394__48_, r_394__47_, r_394__46_, r_394__45_, r_394__44_, r_394__43_, r_394__42_, r_394__41_, r_394__40_, r_394__39_, r_394__38_, r_394__37_, r_394__36_, r_394__35_, r_394__34_, r_394__33_, r_394__32_, r_394__31_, r_394__30_, r_394__29_, r_394__28_, r_394__27_, r_394__26_, r_394__25_, r_394__24_, r_394__23_, r_394__22_, r_394__21_, r_394__20_, r_394__19_, r_394__18_, r_394__17_, r_394__16_, r_394__15_, r_394__14_, r_394__13_, r_394__12_, r_394__11_, r_394__10_, r_394__9_, r_394__8_, r_394__7_, r_394__6_, r_394__5_, r_394__4_, r_394__3_, r_394__2_, r_394__1_, r_394__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N787)? data_i : 1'b0;
  assign N786 = sel_i[786];
  assign N787 = N2993;
  assign { r_n_394__63_, r_n_394__62_, r_n_394__61_, r_n_394__60_, r_n_394__59_, r_n_394__58_, r_n_394__57_, r_n_394__56_, r_n_394__55_, r_n_394__54_, r_n_394__53_, r_n_394__52_, r_n_394__51_, r_n_394__50_, r_n_394__49_, r_n_394__48_, r_n_394__47_, r_n_394__46_, r_n_394__45_, r_n_394__44_, r_n_394__43_, r_n_394__42_, r_n_394__41_, r_n_394__40_, r_n_394__39_, r_n_394__38_, r_n_394__37_, r_n_394__36_, r_n_394__35_, r_n_394__34_, r_n_394__33_, r_n_394__32_, r_n_394__31_, r_n_394__30_, r_n_394__29_, r_n_394__28_, r_n_394__27_, r_n_394__26_, r_n_394__25_, r_n_394__24_, r_n_394__23_, r_n_394__22_, r_n_394__21_, r_n_394__20_, r_n_394__19_, r_n_394__18_, r_n_394__17_, r_n_394__16_, r_n_394__15_, r_n_394__14_, r_n_394__13_, r_n_394__12_, r_n_394__11_, r_n_394__10_, r_n_394__9_, r_n_394__8_, r_n_394__7_, r_n_394__6_, r_n_394__5_, r_n_394__4_, r_n_394__3_, r_n_394__2_, r_n_394__1_, r_n_394__0_ } = (N788)? { r_395__63_, r_395__62_, r_395__61_, r_395__60_, r_395__59_, r_395__58_, r_395__57_, r_395__56_, r_395__55_, r_395__54_, r_395__53_, r_395__52_, r_395__51_, r_395__50_, r_395__49_, r_395__48_, r_395__47_, r_395__46_, r_395__45_, r_395__44_, r_395__43_, r_395__42_, r_395__41_, r_395__40_, r_395__39_, r_395__38_, r_395__37_, r_395__36_, r_395__35_, r_395__34_, r_395__33_, r_395__32_, r_395__31_, r_395__30_, r_395__29_, r_395__28_, r_395__27_, r_395__26_, r_395__25_, r_395__24_, r_395__23_, r_395__22_, r_395__21_, r_395__20_, r_395__19_, r_395__18_, r_395__17_, r_395__16_, r_395__15_, r_395__14_, r_395__13_, r_395__12_, r_395__11_, r_395__10_, r_395__9_, r_395__8_, r_395__7_, r_395__6_, r_395__5_, r_395__4_, r_395__3_, r_395__2_, r_395__1_, r_395__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N789)? data_i : 1'b0;
  assign N788 = sel_i[788];
  assign N789 = N2998;
  assign { r_n_395__63_, r_n_395__62_, r_n_395__61_, r_n_395__60_, r_n_395__59_, r_n_395__58_, r_n_395__57_, r_n_395__56_, r_n_395__55_, r_n_395__54_, r_n_395__53_, r_n_395__52_, r_n_395__51_, r_n_395__50_, r_n_395__49_, r_n_395__48_, r_n_395__47_, r_n_395__46_, r_n_395__45_, r_n_395__44_, r_n_395__43_, r_n_395__42_, r_n_395__41_, r_n_395__40_, r_n_395__39_, r_n_395__38_, r_n_395__37_, r_n_395__36_, r_n_395__35_, r_n_395__34_, r_n_395__33_, r_n_395__32_, r_n_395__31_, r_n_395__30_, r_n_395__29_, r_n_395__28_, r_n_395__27_, r_n_395__26_, r_n_395__25_, r_n_395__24_, r_n_395__23_, r_n_395__22_, r_n_395__21_, r_n_395__20_, r_n_395__19_, r_n_395__18_, r_n_395__17_, r_n_395__16_, r_n_395__15_, r_n_395__14_, r_n_395__13_, r_n_395__12_, r_n_395__11_, r_n_395__10_, r_n_395__9_, r_n_395__8_, r_n_395__7_, r_n_395__6_, r_n_395__5_, r_n_395__4_, r_n_395__3_, r_n_395__2_, r_n_395__1_, r_n_395__0_ } = (N790)? { r_396__63_, r_396__62_, r_396__61_, r_396__60_, r_396__59_, r_396__58_, r_396__57_, r_396__56_, r_396__55_, r_396__54_, r_396__53_, r_396__52_, r_396__51_, r_396__50_, r_396__49_, r_396__48_, r_396__47_, r_396__46_, r_396__45_, r_396__44_, r_396__43_, r_396__42_, r_396__41_, r_396__40_, r_396__39_, r_396__38_, r_396__37_, r_396__36_, r_396__35_, r_396__34_, r_396__33_, r_396__32_, r_396__31_, r_396__30_, r_396__29_, r_396__28_, r_396__27_, r_396__26_, r_396__25_, r_396__24_, r_396__23_, r_396__22_, r_396__21_, r_396__20_, r_396__19_, r_396__18_, r_396__17_, r_396__16_, r_396__15_, r_396__14_, r_396__13_, r_396__12_, r_396__11_, r_396__10_, r_396__9_, r_396__8_, r_396__7_, r_396__6_, r_396__5_, r_396__4_, r_396__3_, r_396__2_, r_396__1_, r_396__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N791)? data_i : 1'b0;
  assign N790 = sel_i[790];
  assign N791 = N3003;
  assign { r_n_396__63_, r_n_396__62_, r_n_396__61_, r_n_396__60_, r_n_396__59_, r_n_396__58_, r_n_396__57_, r_n_396__56_, r_n_396__55_, r_n_396__54_, r_n_396__53_, r_n_396__52_, r_n_396__51_, r_n_396__50_, r_n_396__49_, r_n_396__48_, r_n_396__47_, r_n_396__46_, r_n_396__45_, r_n_396__44_, r_n_396__43_, r_n_396__42_, r_n_396__41_, r_n_396__40_, r_n_396__39_, r_n_396__38_, r_n_396__37_, r_n_396__36_, r_n_396__35_, r_n_396__34_, r_n_396__33_, r_n_396__32_, r_n_396__31_, r_n_396__30_, r_n_396__29_, r_n_396__28_, r_n_396__27_, r_n_396__26_, r_n_396__25_, r_n_396__24_, r_n_396__23_, r_n_396__22_, r_n_396__21_, r_n_396__20_, r_n_396__19_, r_n_396__18_, r_n_396__17_, r_n_396__16_, r_n_396__15_, r_n_396__14_, r_n_396__13_, r_n_396__12_, r_n_396__11_, r_n_396__10_, r_n_396__9_, r_n_396__8_, r_n_396__7_, r_n_396__6_, r_n_396__5_, r_n_396__4_, r_n_396__3_, r_n_396__2_, r_n_396__1_, r_n_396__0_ } = (N792)? { r_397__63_, r_397__62_, r_397__61_, r_397__60_, r_397__59_, r_397__58_, r_397__57_, r_397__56_, r_397__55_, r_397__54_, r_397__53_, r_397__52_, r_397__51_, r_397__50_, r_397__49_, r_397__48_, r_397__47_, r_397__46_, r_397__45_, r_397__44_, r_397__43_, r_397__42_, r_397__41_, r_397__40_, r_397__39_, r_397__38_, r_397__37_, r_397__36_, r_397__35_, r_397__34_, r_397__33_, r_397__32_, r_397__31_, r_397__30_, r_397__29_, r_397__28_, r_397__27_, r_397__26_, r_397__25_, r_397__24_, r_397__23_, r_397__22_, r_397__21_, r_397__20_, r_397__19_, r_397__18_, r_397__17_, r_397__16_, r_397__15_, r_397__14_, r_397__13_, r_397__12_, r_397__11_, r_397__10_, r_397__9_, r_397__8_, r_397__7_, r_397__6_, r_397__5_, r_397__4_, r_397__3_, r_397__2_, r_397__1_, r_397__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N793)? data_i : 1'b0;
  assign N792 = sel_i[792];
  assign N793 = N3008;
  assign { r_n_397__63_, r_n_397__62_, r_n_397__61_, r_n_397__60_, r_n_397__59_, r_n_397__58_, r_n_397__57_, r_n_397__56_, r_n_397__55_, r_n_397__54_, r_n_397__53_, r_n_397__52_, r_n_397__51_, r_n_397__50_, r_n_397__49_, r_n_397__48_, r_n_397__47_, r_n_397__46_, r_n_397__45_, r_n_397__44_, r_n_397__43_, r_n_397__42_, r_n_397__41_, r_n_397__40_, r_n_397__39_, r_n_397__38_, r_n_397__37_, r_n_397__36_, r_n_397__35_, r_n_397__34_, r_n_397__33_, r_n_397__32_, r_n_397__31_, r_n_397__30_, r_n_397__29_, r_n_397__28_, r_n_397__27_, r_n_397__26_, r_n_397__25_, r_n_397__24_, r_n_397__23_, r_n_397__22_, r_n_397__21_, r_n_397__20_, r_n_397__19_, r_n_397__18_, r_n_397__17_, r_n_397__16_, r_n_397__15_, r_n_397__14_, r_n_397__13_, r_n_397__12_, r_n_397__11_, r_n_397__10_, r_n_397__9_, r_n_397__8_, r_n_397__7_, r_n_397__6_, r_n_397__5_, r_n_397__4_, r_n_397__3_, r_n_397__2_, r_n_397__1_, r_n_397__0_ } = (N794)? { r_398__63_, r_398__62_, r_398__61_, r_398__60_, r_398__59_, r_398__58_, r_398__57_, r_398__56_, r_398__55_, r_398__54_, r_398__53_, r_398__52_, r_398__51_, r_398__50_, r_398__49_, r_398__48_, r_398__47_, r_398__46_, r_398__45_, r_398__44_, r_398__43_, r_398__42_, r_398__41_, r_398__40_, r_398__39_, r_398__38_, r_398__37_, r_398__36_, r_398__35_, r_398__34_, r_398__33_, r_398__32_, r_398__31_, r_398__30_, r_398__29_, r_398__28_, r_398__27_, r_398__26_, r_398__25_, r_398__24_, r_398__23_, r_398__22_, r_398__21_, r_398__20_, r_398__19_, r_398__18_, r_398__17_, r_398__16_, r_398__15_, r_398__14_, r_398__13_, r_398__12_, r_398__11_, r_398__10_, r_398__9_, r_398__8_, r_398__7_, r_398__6_, r_398__5_, r_398__4_, r_398__3_, r_398__2_, r_398__1_, r_398__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N795)? data_i : 1'b0;
  assign N794 = sel_i[794];
  assign N795 = N3013;
  assign { r_n_398__63_, r_n_398__62_, r_n_398__61_, r_n_398__60_, r_n_398__59_, r_n_398__58_, r_n_398__57_, r_n_398__56_, r_n_398__55_, r_n_398__54_, r_n_398__53_, r_n_398__52_, r_n_398__51_, r_n_398__50_, r_n_398__49_, r_n_398__48_, r_n_398__47_, r_n_398__46_, r_n_398__45_, r_n_398__44_, r_n_398__43_, r_n_398__42_, r_n_398__41_, r_n_398__40_, r_n_398__39_, r_n_398__38_, r_n_398__37_, r_n_398__36_, r_n_398__35_, r_n_398__34_, r_n_398__33_, r_n_398__32_, r_n_398__31_, r_n_398__30_, r_n_398__29_, r_n_398__28_, r_n_398__27_, r_n_398__26_, r_n_398__25_, r_n_398__24_, r_n_398__23_, r_n_398__22_, r_n_398__21_, r_n_398__20_, r_n_398__19_, r_n_398__18_, r_n_398__17_, r_n_398__16_, r_n_398__15_, r_n_398__14_, r_n_398__13_, r_n_398__12_, r_n_398__11_, r_n_398__10_, r_n_398__9_, r_n_398__8_, r_n_398__7_, r_n_398__6_, r_n_398__5_, r_n_398__4_, r_n_398__3_, r_n_398__2_, r_n_398__1_, r_n_398__0_ } = (N796)? { r_399__63_, r_399__62_, r_399__61_, r_399__60_, r_399__59_, r_399__58_, r_399__57_, r_399__56_, r_399__55_, r_399__54_, r_399__53_, r_399__52_, r_399__51_, r_399__50_, r_399__49_, r_399__48_, r_399__47_, r_399__46_, r_399__45_, r_399__44_, r_399__43_, r_399__42_, r_399__41_, r_399__40_, r_399__39_, r_399__38_, r_399__37_, r_399__36_, r_399__35_, r_399__34_, r_399__33_, r_399__32_, r_399__31_, r_399__30_, r_399__29_, r_399__28_, r_399__27_, r_399__26_, r_399__25_, r_399__24_, r_399__23_, r_399__22_, r_399__21_, r_399__20_, r_399__19_, r_399__18_, r_399__17_, r_399__16_, r_399__15_, r_399__14_, r_399__13_, r_399__12_, r_399__11_, r_399__10_, r_399__9_, r_399__8_, r_399__7_, r_399__6_, r_399__5_, r_399__4_, r_399__3_, r_399__2_, r_399__1_, r_399__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N797)? data_i : 1'b0;
  assign N796 = sel_i[796];
  assign N797 = N3018;
  assign { r_n_399__63_, r_n_399__62_, r_n_399__61_, r_n_399__60_, r_n_399__59_, r_n_399__58_, r_n_399__57_, r_n_399__56_, r_n_399__55_, r_n_399__54_, r_n_399__53_, r_n_399__52_, r_n_399__51_, r_n_399__50_, r_n_399__49_, r_n_399__48_, r_n_399__47_, r_n_399__46_, r_n_399__45_, r_n_399__44_, r_n_399__43_, r_n_399__42_, r_n_399__41_, r_n_399__40_, r_n_399__39_, r_n_399__38_, r_n_399__37_, r_n_399__36_, r_n_399__35_, r_n_399__34_, r_n_399__33_, r_n_399__32_, r_n_399__31_, r_n_399__30_, r_n_399__29_, r_n_399__28_, r_n_399__27_, r_n_399__26_, r_n_399__25_, r_n_399__24_, r_n_399__23_, r_n_399__22_, r_n_399__21_, r_n_399__20_, r_n_399__19_, r_n_399__18_, r_n_399__17_, r_n_399__16_, r_n_399__15_, r_n_399__14_, r_n_399__13_, r_n_399__12_, r_n_399__11_, r_n_399__10_, r_n_399__9_, r_n_399__8_, r_n_399__7_, r_n_399__6_, r_n_399__5_, r_n_399__4_, r_n_399__3_, r_n_399__2_, r_n_399__1_, r_n_399__0_ } = (N798)? { r_400__63_, r_400__62_, r_400__61_, r_400__60_, r_400__59_, r_400__58_, r_400__57_, r_400__56_, r_400__55_, r_400__54_, r_400__53_, r_400__52_, r_400__51_, r_400__50_, r_400__49_, r_400__48_, r_400__47_, r_400__46_, r_400__45_, r_400__44_, r_400__43_, r_400__42_, r_400__41_, r_400__40_, r_400__39_, r_400__38_, r_400__37_, r_400__36_, r_400__35_, r_400__34_, r_400__33_, r_400__32_, r_400__31_, r_400__30_, r_400__29_, r_400__28_, r_400__27_, r_400__26_, r_400__25_, r_400__24_, r_400__23_, r_400__22_, r_400__21_, r_400__20_, r_400__19_, r_400__18_, r_400__17_, r_400__16_, r_400__15_, r_400__14_, r_400__13_, r_400__12_, r_400__11_, r_400__10_, r_400__9_, r_400__8_, r_400__7_, r_400__6_, r_400__5_, r_400__4_, r_400__3_, r_400__2_, r_400__1_, r_400__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N799)? data_i : 1'b0;
  assign N798 = sel_i[798];
  assign N799 = N3023;
  assign { r_n_400__63_, r_n_400__62_, r_n_400__61_, r_n_400__60_, r_n_400__59_, r_n_400__58_, r_n_400__57_, r_n_400__56_, r_n_400__55_, r_n_400__54_, r_n_400__53_, r_n_400__52_, r_n_400__51_, r_n_400__50_, r_n_400__49_, r_n_400__48_, r_n_400__47_, r_n_400__46_, r_n_400__45_, r_n_400__44_, r_n_400__43_, r_n_400__42_, r_n_400__41_, r_n_400__40_, r_n_400__39_, r_n_400__38_, r_n_400__37_, r_n_400__36_, r_n_400__35_, r_n_400__34_, r_n_400__33_, r_n_400__32_, r_n_400__31_, r_n_400__30_, r_n_400__29_, r_n_400__28_, r_n_400__27_, r_n_400__26_, r_n_400__25_, r_n_400__24_, r_n_400__23_, r_n_400__22_, r_n_400__21_, r_n_400__20_, r_n_400__19_, r_n_400__18_, r_n_400__17_, r_n_400__16_, r_n_400__15_, r_n_400__14_, r_n_400__13_, r_n_400__12_, r_n_400__11_, r_n_400__10_, r_n_400__9_, r_n_400__8_, r_n_400__7_, r_n_400__6_, r_n_400__5_, r_n_400__4_, r_n_400__3_, r_n_400__2_, r_n_400__1_, r_n_400__0_ } = (N800)? { r_401__63_, r_401__62_, r_401__61_, r_401__60_, r_401__59_, r_401__58_, r_401__57_, r_401__56_, r_401__55_, r_401__54_, r_401__53_, r_401__52_, r_401__51_, r_401__50_, r_401__49_, r_401__48_, r_401__47_, r_401__46_, r_401__45_, r_401__44_, r_401__43_, r_401__42_, r_401__41_, r_401__40_, r_401__39_, r_401__38_, r_401__37_, r_401__36_, r_401__35_, r_401__34_, r_401__33_, r_401__32_, r_401__31_, r_401__30_, r_401__29_, r_401__28_, r_401__27_, r_401__26_, r_401__25_, r_401__24_, r_401__23_, r_401__22_, r_401__21_, r_401__20_, r_401__19_, r_401__18_, r_401__17_, r_401__16_, r_401__15_, r_401__14_, r_401__13_, r_401__12_, r_401__11_, r_401__10_, r_401__9_, r_401__8_, r_401__7_, r_401__6_, r_401__5_, r_401__4_, r_401__3_, r_401__2_, r_401__1_, r_401__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N801)? data_i : 1'b0;
  assign N800 = sel_i[800];
  assign N801 = N3028;
  assign { r_n_401__63_, r_n_401__62_, r_n_401__61_, r_n_401__60_, r_n_401__59_, r_n_401__58_, r_n_401__57_, r_n_401__56_, r_n_401__55_, r_n_401__54_, r_n_401__53_, r_n_401__52_, r_n_401__51_, r_n_401__50_, r_n_401__49_, r_n_401__48_, r_n_401__47_, r_n_401__46_, r_n_401__45_, r_n_401__44_, r_n_401__43_, r_n_401__42_, r_n_401__41_, r_n_401__40_, r_n_401__39_, r_n_401__38_, r_n_401__37_, r_n_401__36_, r_n_401__35_, r_n_401__34_, r_n_401__33_, r_n_401__32_, r_n_401__31_, r_n_401__30_, r_n_401__29_, r_n_401__28_, r_n_401__27_, r_n_401__26_, r_n_401__25_, r_n_401__24_, r_n_401__23_, r_n_401__22_, r_n_401__21_, r_n_401__20_, r_n_401__19_, r_n_401__18_, r_n_401__17_, r_n_401__16_, r_n_401__15_, r_n_401__14_, r_n_401__13_, r_n_401__12_, r_n_401__11_, r_n_401__10_, r_n_401__9_, r_n_401__8_, r_n_401__7_, r_n_401__6_, r_n_401__5_, r_n_401__4_, r_n_401__3_, r_n_401__2_, r_n_401__1_, r_n_401__0_ } = (N802)? { r_402__63_, r_402__62_, r_402__61_, r_402__60_, r_402__59_, r_402__58_, r_402__57_, r_402__56_, r_402__55_, r_402__54_, r_402__53_, r_402__52_, r_402__51_, r_402__50_, r_402__49_, r_402__48_, r_402__47_, r_402__46_, r_402__45_, r_402__44_, r_402__43_, r_402__42_, r_402__41_, r_402__40_, r_402__39_, r_402__38_, r_402__37_, r_402__36_, r_402__35_, r_402__34_, r_402__33_, r_402__32_, r_402__31_, r_402__30_, r_402__29_, r_402__28_, r_402__27_, r_402__26_, r_402__25_, r_402__24_, r_402__23_, r_402__22_, r_402__21_, r_402__20_, r_402__19_, r_402__18_, r_402__17_, r_402__16_, r_402__15_, r_402__14_, r_402__13_, r_402__12_, r_402__11_, r_402__10_, r_402__9_, r_402__8_, r_402__7_, r_402__6_, r_402__5_, r_402__4_, r_402__3_, r_402__2_, r_402__1_, r_402__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N803)? data_i : 1'b0;
  assign N802 = sel_i[802];
  assign N803 = N3033;
  assign { r_n_402__63_, r_n_402__62_, r_n_402__61_, r_n_402__60_, r_n_402__59_, r_n_402__58_, r_n_402__57_, r_n_402__56_, r_n_402__55_, r_n_402__54_, r_n_402__53_, r_n_402__52_, r_n_402__51_, r_n_402__50_, r_n_402__49_, r_n_402__48_, r_n_402__47_, r_n_402__46_, r_n_402__45_, r_n_402__44_, r_n_402__43_, r_n_402__42_, r_n_402__41_, r_n_402__40_, r_n_402__39_, r_n_402__38_, r_n_402__37_, r_n_402__36_, r_n_402__35_, r_n_402__34_, r_n_402__33_, r_n_402__32_, r_n_402__31_, r_n_402__30_, r_n_402__29_, r_n_402__28_, r_n_402__27_, r_n_402__26_, r_n_402__25_, r_n_402__24_, r_n_402__23_, r_n_402__22_, r_n_402__21_, r_n_402__20_, r_n_402__19_, r_n_402__18_, r_n_402__17_, r_n_402__16_, r_n_402__15_, r_n_402__14_, r_n_402__13_, r_n_402__12_, r_n_402__11_, r_n_402__10_, r_n_402__9_, r_n_402__8_, r_n_402__7_, r_n_402__6_, r_n_402__5_, r_n_402__4_, r_n_402__3_, r_n_402__2_, r_n_402__1_, r_n_402__0_ } = (N804)? { r_403__63_, r_403__62_, r_403__61_, r_403__60_, r_403__59_, r_403__58_, r_403__57_, r_403__56_, r_403__55_, r_403__54_, r_403__53_, r_403__52_, r_403__51_, r_403__50_, r_403__49_, r_403__48_, r_403__47_, r_403__46_, r_403__45_, r_403__44_, r_403__43_, r_403__42_, r_403__41_, r_403__40_, r_403__39_, r_403__38_, r_403__37_, r_403__36_, r_403__35_, r_403__34_, r_403__33_, r_403__32_, r_403__31_, r_403__30_, r_403__29_, r_403__28_, r_403__27_, r_403__26_, r_403__25_, r_403__24_, r_403__23_, r_403__22_, r_403__21_, r_403__20_, r_403__19_, r_403__18_, r_403__17_, r_403__16_, r_403__15_, r_403__14_, r_403__13_, r_403__12_, r_403__11_, r_403__10_, r_403__9_, r_403__8_, r_403__7_, r_403__6_, r_403__5_, r_403__4_, r_403__3_, r_403__2_, r_403__1_, r_403__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N805)? data_i : 1'b0;
  assign N804 = sel_i[804];
  assign N805 = N3038;
  assign { r_n_403__63_, r_n_403__62_, r_n_403__61_, r_n_403__60_, r_n_403__59_, r_n_403__58_, r_n_403__57_, r_n_403__56_, r_n_403__55_, r_n_403__54_, r_n_403__53_, r_n_403__52_, r_n_403__51_, r_n_403__50_, r_n_403__49_, r_n_403__48_, r_n_403__47_, r_n_403__46_, r_n_403__45_, r_n_403__44_, r_n_403__43_, r_n_403__42_, r_n_403__41_, r_n_403__40_, r_n_403__39_, r_n_403__38_, r_n_403__37_, r_n_403__36_, r_n_403__35_, r_n_403__34_, r_n_403__33_, r_n_403__32_, r_n_403__31_, r_n_403__30_, r_n_403__29_, r_n_403__28_, r_n_403__27_, r_n_403__26_, r_n_403__25_, r_n_403__24_, r_n_403__23_, r_n_403__22_, r_n_403__21_, r_n_403__20_, r_n_403__19_, r_n_403__18_, r_n_403__17_, r_n_403__16_, r_n_403__15_, r_n_403__14_, r_n_403__13_, r_n_403__12_, r_n_403__11_, r_n_403__10_, r_n_403__9_, r_n_403__8_, r_n_403__7_, r_n_403__6_, r_n_403__5_, r_n_403__4_, r_n_403__3_, r_n_403__2_, r_n_403__1_, r_n_403__0_ } = (N806)? { r_404__63_, r_404__62_, r_404__61_, r_404__60_, r_404__59_, r_404__58_, r_404__57_, r_404__56_, r_404__55_, r_404__54_, r_404__53_, r_404__52_, r_404__51_, r_404__50_, r_404__49_, r_404__48_, r_404__47_, r_404__46_, r_404__45_, r_404__44_, r_404__43_, r_404__42_, r_404__41_, r_404__40_, r_404__39_, r_404__38_, r_404__37_, r_404__36_, r_404__35_, r_404__34_, r_404__33_, r_404__32_, r_404__31_, r_404__30_, r_404__29_, r_404__28_, r_404__27_, r_404__26_, r_404__25_, r_404__24_, r_404__23_, r_404__22_, r_404__21_, r_404__20_, r_404__19_, r_404__18_, r_404__17_, r_404__16_, r_404__15_, r_404__14_, r_404__13_, r_404__12_, r_404__11_, r_404__10_, r_404__9_, r_404__8_, r_404__7_, r_404__6_, r_404__5_, r_404__4_, r_404__3_, r_404__2_, r_404__1_, r_404__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N807)? data_i : 1'b0;
  assign N806 = sel_i[806];
  assign N807 = N3043;
  assign { r_n_404__63_, r_n_404__62_, r_n_404__61_, r_n_404__60_, r_n_404__59_, r_n_404__58_, r_n_404__57_, r_n_404__56_, r_n_404__55_, r_n_404__54_, r_n_404__53_, r_n_404__52_, r_n_404__51_, r_n_404__50_, r_n_404__49_, r_n_404__48_, r_n_404__47_, r_n_404__46_, r_n_404__45_, r_n_404__44_, r_n_404__43_, r_n_404__42_, r_n_404__41_, r_n_404__40_, r_n_404__39_, r_n_404__38_, r_n_404__37_, r_n_404__36_, r_n_404__35_, r_n_404__34_, r_n_404__33_, r_n_404__32_, r_n_404__31_, r_n_404__30_, r_n_404__29_, r_n_404__28_, r_n_404__27_, r_n_404__26_, r_n_404__25_, r_n_404__24_, r_n_404__23_, r_n_404__22_, r_n_404__21_, r_n_404__20_, r_n_404__19_, r_n_404__18_, r_n_404__17_, r_n_404__16_, r_n_404__15_, r_n_404__14_, r_n_404__13_, r_n_404__12_, r_n_404__11_, r_n_404__10_, r_n_404__9_, r_n_404__8_, r_n_404__7_, r_n_404__6_, r_n_404__5_, r_n_404__4_, r_n_404__3_, r_n_404__2_, r_n_404__1_, r_n_404__0_ } = (N808)? { r_405__63_, r_405__62_, r_405__61_, r_405__60_, r_405__59_, r_405__58_, r_405__57_, r_405__56_, r_405__55_, r_405__54_, r_405__53_, r_405__52_, r_405__51_, r_405__50_, r_405__49_, r_405__48_, r_405__47_, r_405__46_, r_405__45_, r_405__44_, r_405__43_, r_405__42_, r_405__41_, r_405__40_, r_405__39_, r_405__38_, r_405__37_, r_405__36_, r_405__35_, r_405__34_, r_405__33_, r_405__32_, r_405__31_, r_405__30_, r_405__29_, r_405__28_, r_405__27_, r_405__26_, r_405__25_, r_405__24_, r_405__23_, r_405__22_, r_405__21_, r_405__20_, r_405__19_, r_405__18_, r_405__17_, r_405__16_, r_405__15_, r_405__14_, r_405__13_, r_405__12_, r_405__11_, r_405__10_, r_405__9_, r_405__8_, r_405__7_, r_405__6_, r_405__5_, r_405__4_, r_405__3_, r_405__2_, r_405__1_, r_405__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N809)? data_i : 1'b0;
  assign N808 = sel_i[808];
  assign N809 = N3048;
  assign { r_n_405__63_, r_n_405__62_, r_n_405__61_, r_n_405__60_, r_n_405__59_, r_n_405__58_, r_n_405__57_, r_n_405__56_, r_n_405__55_, r_n_405__54_, r_n_405__53_, r_n_405__52_, r_n_405__51_, r_n_405__50_, r_n_405__49_, r_n_405__48_, r_n_405__47_, r_n_405__46_, r_n_405__45_, r_n_405__44_, r_n_405__43_, r_n_405__42_, r_n_405__41_, r_n_405__40_, r_n_405__39_, r_n_405__38_, r_n_405__37_, r_n_405__36_, r_n_405__35_, r_n_405__34_, r_n_405__33_, r_n_405__32_, r_n_405__31_, r_n_405__30_, r_n_405__29_, r_n_405__28_, r_n_405__27_, r_n_405__26_, r_n_405__25_, r_n_405__24_, r_n_405__23_, r_n_405__22_, r_n_405__21_, r_n_405__20_, r_n_405__19_, r_n_405__18_, r_n_405__17_, r_n_405__16_, r_n_405__15_, r_n_405__14_, r_n_405__13_, r_n_405__12_, r_n_405__11_, r_n_405__10_, r_n_405__9_, r_n_405__8_, r_n_405__7_, r_n_405__6_, r_n_405__5_, r_n_405__4_, r_n_405__3_, r_n_405__2_, r_n_405__1_, r_n_405__0_ } = (N810)? { r_406__63_, r_406__62_, r_406__61_, r_406__60_, r_406__59_, r_406__58_, r_406__57_, r_406__56_, r_406__55_, r_406__54_, r_406__53_, r_406__52_, r_406__51_, r_406__50_, r_406__49_, r_406__48_, r_406__47_, r_406__46_, r_406__45_, r_406__44_, r_406__43_, r_406__42_, r_406__41_, r_406__40_, r_406__39_, r_406__38_, r_406__37_, r_406__36_, r_406__35_, r_406__34_, r_406__33_, r_406__32_, r_406__31_, r_406__30_, r_406__29_, r_406__28_, r_406__27_, r_406__26_, r_406__25_, r_406__24_, r_406__23_, r_406__22_, r_406__21_, r_406__20_, r_406__19_, r_406__18_, r_406__17_, r_406__16_, r_406__15_, r_406__14_, r_406__13_, r_406__12_, r_406__11_, r_406__10_, r_406__9_, r_406__8_, r_406__7_, r_406__6_, r_406__5_, r_406__4_, r_406__3_, r_406__2_, r_406__1_, r_406__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N811)? data_i : 1'b0;
  assign N810 = sel_i[810];
  assign N811 = N3053;
  assign { r_n_406__63_, r_n_406__62_, r_n_406__61_, r_n_406__60_, r_n_406__59_, r_n_406__58_, r_n_406__57_, r_n_406__56_, r_n_406__55_, r_n_406__54_, r_n_406__53_, r_n_406__52_, r_n_406__51_, r_n_406__50_, r_n_406__49_, r_n_406__48_, r_n_406__47_, r_n_406__46_, r_n_406__45_, r_n_406__44_, r_n_406__43_, r_n_406__42_, r_n_406__41_, r_n_406__40_, r_n_406__39_, r_n_406__38_, r_n_406__37_, r_n_406__36_, r_n_406__35_, r_n_406__34_, r_n_406__33_, r_n_406__32_, r_n_406__31_, r_n_406__30_, r_n_406__29_, r_n_406__28_, r_n_406__27_, r_n_406__26_, r_n_406__25_, r_n_406__24_, r_n_406__23_, r_n_406__22_, r_n_406__21_, r_n_406__20_, r_n_406__19_, r_n_406__18_, r_n_406__17_, r_n_406__16_, r_n_406__15_, r_n_406__14_, r_n_406__13_, r_n_406__12_, r_n_406__11_, r_n_406__10_, r_n_406__9_, r_n_406__8_, r_n_406__7_, r_n_406__6_, r_n_406__5_, r_n_406__4_, r_n_406__3_, r_n_406__2_, r_n_406__1_, r_n_406__0_ } = (N812)? { r_407__63_, r_407__62_, r_407__61_, r_407__60_, r_407__59_, r_407__58_, r_407__57_, r_407__56_, r_407__55_, r_407__54_, r_407__53_, r_407__52_, r_407__51_, r_407__50_, r_407__49_, r_407__48_, r_407__47_, r_407__46_, r_407__45_, r_407__44_, r_407__43_, r_407__42_, r_407__41_, r_407__40_, r_407__39_, r_407__38_, r_407__37_, r_407__36_, r_407__35_, r_407__34_, r_407__33_, r_407__32_, r_407__31_, r_407__30_, r_407__29_, r_407__28_, r_407__27_, r_407__26_, r_407__25_, r_407__24_, r_407__23_, r_407__22_, r_407__21_, r_407__20_, r_407__19_, r_407__18_, r_407__17_, r_407__16_, r_407__15_, r_407__14_, r_407__13_, r_407__12_, r_407__11_, r_407__10_, r_407__9_, r_407__8_, r_407__7_, r_407__6_, r_407__5_, r_407__4_, r_407__3_, r_407__2_, r_407__1_, r_407__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N813)? data_i : 1'b0;
  assign N812 = sel_i[812];
  assign N813 = N3058;
  assign { r_n_407__63_, r_n_407__62_, r_n_407__61_, r_n_407__60_, r_n_407__59_, r_n_407__58_, r_n_407__57_, r_n_407__56_, r_n_407__55_, r_n_407__54_, r_n_407__53_, r_n_407__52_, r_n_407__51_, r_n_407__50_, r_n_407__49_, r_n_407__48_, r_n_407__47_, r_n_407__46_, r_n_407__45_, r_n_407__44_, r_n_407__43_, r_n_407__42_, r_n_407__41_, r_n_407__40_, r_n_407__39_, r_n_407__38_, r_n_407__37_, r_n_407__36_, r_n_407__35_, r_n_407__34_, r_n_407__33_, r_n_407__32_, r_n_407__31_, r_n_407__30_, r_n_407__29_, r_n_407__28_, r_n_407__27_, r_n_407__26_, r_n_407__25_, r_n_407__24_, r_n_407__23_, r_n_407__22_, r_n_407__21_, r_n_407__20_, r_n_407__19_, r_n_407__18_, r_n_407__17_, r_n_407__16_, r_n_407__15_, r_n_407__14_, r_n_407__13_, r_n_407__12_, r_n_407__11_, r_n_407__10_, r_n_407__9_, r_n_407__8_, r_n_407__7_, r_n_407__6_, r_n_407__5_, r_n_407__4_, r_n_407__3_, r_n_407__2_, r_n_407__1_, r_n_407__0_ } = (N814)? { r_408__63_, r_408__62_, r_408__61_, r_408__60_, r_408__59_, r_408__58_, r_408__57_, r_408__56_, r_408__55_, r_408__54_, r_408__53_, r_408__52_, r_408__51_, r_408__50_, r_408__49_, r_408__48_, r_408__47_, r_408__46_, r_408__45_, r_408__44_, r_408__43_, r_408__42_, r_408__41_, r_408__40_, r_408__39_, r_408__38_, r_408__37_, r_408__36_, r_408__35_, r_408__34_, r_408__33_, r_408__32_, r_408__31_, r_408__30_, r_408__29_, r_408__28_, r_408__27_, r_408__26_, r_408__25_, r_408__24_, r_408__23_, r_408__22_, r_408__21_, r_408__20_, r_408__19_, r_408__18_, r_408__17_, r_408__16_, r_408__15_, r_408__14_, r_408__13_, r_408__12_, r_408__11_, r_408__10_, r_408__9_, r_408__8_, r_408__7_, r_408__6_, r_408__5_, r_408__4_, r_408__3_, r_408__2_, r_408__1_, r_408__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N815)? data_i : 1'b0;
  assign N814 = sel_i[814];
  assign N815 = N3063;
  assign { r_n_408__63_, r_n_408__62_, r_n_408__61_, r_n_408__60_, r_n_408__59_, r_n_408__58_, r_n_408__57_, r_n_408__56_, r_n_408__55_, r_n_408__54_, r_n_408__53_, r_n_408__52_, r_n_408__51_, r_n_408__50_, r_n_408__49_, r_n_408__48_, r_n_408__47_, r_n_408__46_, r_n_408__45_, r_n_408__44_, r_n_408__43_, r_n_408__42_, r_n_408__41_, r_n_408__40_, r_n_408__39_, r_n_408__38_, r_n_408__37_, r_n_408__36_, r_n_408__35_, r_n_408__34_, r_n_408__33_, r_n_408__32_, r_n_408__31_, r_n_408__30_, r_n_408__29_, r_n_408__28_, r_n_408__27_, r_n_408__26_, r_n_408__25_, r_n_408__24_, r_n_408__23_, r_n_408__22_, r_n_408__21_, r_n_408__20_, r_n_408__19_, r_n_408__18_, r_n_408__17_, r_n_408__16_, r_n_408__15_, r_n_408__14_, r_n_408__13_, r_n_408__12_, r_n_408__11_, r_n_408__10_, r_n_408__9_, r_n_408__8_, r_n_408__7_, r_n_408__6_, r_n_408__5_, r_n_408__4_, r_n_408__3_, r_n_408__2_, r_n_408__1_, r_n_408__0_ } = (N816)? { r_409__63_, r_409__62_, r_409__61_, r_409__60_, r_409__59_, r_409__58_, r_409__57_, r_409__56_, r_409__55_, r_409__54_, r_409__53_, r_409__52_, r_409__51_, r_409__50_, r_409__49_, r_409__48_, r_409__47_, r_409__46_, r_409__45_, r_409__44_, r_409__43_, r_409__42_, r_409__41_, r_409__40_, r_409__39_, r_409__38_, r_409__37_, r_409__36_, r_409__35_, r_409__34_, r_409__33_, r_409__32_, r_409__31_, r_409__30_, r_409__29_, r_409__28_, r_409__27_, r_409__26_, r_409__25_, r_409__24_, r_409__23_, r_409__22_, r_409__21_, r_409__20_, r_409__19_, r_409__18_, r_409__17_, r_409__16_, r_409__15_, r_409__14_, r_409__13_, r_409__12_, r_409__11_, r_409__10_, r_409__9_, r_409__8_, r_409__7_, r_409__6_, r_409__5_, r_409__4_, r_409__3_, r_409__2_, r_409__1_, r_409__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N817)? data_i : 1'b0;
  assign N816 = sel_i[816];
  assign N817 = N3068;
  assign { r_n_409__63_, r_n_409__62_, r_n_409__61_, r_n_409__60_, r_n_409__59_, r_n_409__58_, r_n_409__57_, r_n_409__56_, r_n_409__55_, r_n_409__54_, r_n_409__53_, r_n_409__52_, r_n_409__51_, r_n_409__50_, r_n_409__49_, r_n_409__48_, r_n_409__47_, r_n_409__46_, r_n_409__45_, r_n_409__44_, r_n_409__43_, r_n_409__42_, r_n_409__41_, r_n_409__40_, r_n_409__39_, r_n_409__38_, r_n_409__37_, r_n_409__36_, r_n_409__35_, r_n_409__34_, r_n_409__33_, r_n_409__32_, r_n_409__31_, r_n_409__30_, r_n_409__29_, r_n_409__28_, r_n_409__27_, r_n_409__26_, r_n_409__25_, r_n_409__24_, r_n_409__23_, r_n_409__22_, r_n_409__21_, r_n_409__20_, r_n_409__19_, r_n_409__18_, r_n_409__17_, r_n_409__16_, r_n_409__15_, r_n_409__14_, r_n_409__13_, r_n_409__12_, r_n_409__11_, r_n_409__10_, r_n_409__9_, r_n_409__8_, r_n_409__7_, r_n_409__6_, r_n_409__5_, r_n_409__4_, r_n_409__3_, r_n_409__2_, r_n_409__1_, r_n_409__0_ } = (N818)? { r_410__63_, r_410__62_, r_410__61_, r_410__60_, r_410__59_, r_410__58_, r_410__57_, r_410__56_, r_410__55_, r_410__54_, r_410__53_, r_410__52_, r_410__51_, r_410__50_, r_410__49_, r_410__48_, r_410__47_, r_410__46_, r_410__45_, r_410__44_, r_410__43_, r_410__42_, r_410__41_, r_410__40_, r_410__39_, r_410__38_, r_410__37_, r_410__36_, r_410__35_, r_410__34_, r_410__33_, r_410__32_, r_410__31_, r_410__30_, r_410__29_, r_410__28_, r_410__27_, r_410__26_, r_410__25_, r_410__24_, r_410__23_, r_410__22_, r_410__21_, r_410__20_, r_410__19_, r_410__18_, r_410__17_, r_410__16_, r_410__15_, r_410__14_, r_410__13_, r_410__12_, r_410__11_, r_410__10_, r_410__9_, r_410__8_, r_410__7_, r_410__6_, r_410__5_, r_410__4_, r_410__3_, r_410__2_, r_410__1_, r_410__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N819)? data_i : 1'b0;
  assign N818 = sel_i[818];
  assign N819 = N3073;
  assign { r_n_410__63_, r_n_410__62_, r_n_410__61_, r_n_410__60_, r_n_410__59_, r_n_410__58_, r_n_410__57_, r_n_410__56_, r_n_410__55_, r_n_410__54_, r_n_410__53_, r_n_410__52_, r_n_410__51_, r_n_410__50_, r_n_410__49_, r_n_410__48_, r_n_410__47_, r_n_410__46_, r_n_410__45_, r_n_410__44_, r_n_410__43_, r_n_410__42_, r_n_410__41_, r_n_410__40_, r_n_410__39_, r_n_410__38_, r_n_410__37_, r_n_410__36_, r_n_410__35_, r_n_410__34_, r_n_410__33_, r_n_410__32_, r_n_410__31_, r_n_410__30_, r_n_410__29_, r_n_410__28_, r_n_410__27_, r_n_410__26_, r_n_410__25_, r_n_410__24_, r_n_410__23_, r_n_410__22_, r_n_410__21_, r_n_410__20_, r_n_410__19_, r_n_410__18_, r_n_410__17_, r_n_410__16_, r_n_410__15_, r_n_410__14_, r_n_410__13_, r_n_410__12_, r_n_410__11_, r_n_410__10_, r_n_410__9_, r_n_410__8_, r_n_410__7_, r_n_410__6_, r_n_410__5_, r_n_410__4_, r_n_410__3_, r_n_410__2_, r_n_410__1_, r_n_410__0_ } = (N820)? { r_411__63_, r_411__62_, r_411__61_, r_411__60_, r_411__59_, r_411__58_, r_411__57_, r_411__56_, r_411__55_, r_411__54_, r_411__53_, r_411__52_, r_411__51_, r_411__50_, r_411__49_, r_411__48_, r_411__47_, r_411__46_, r_411__45_, r_411__44_, r_411__43_, r_411__42_, r_411__41_, r_411__40_, r_411__39_, r_411__38_, r_411__37_, r_411__36_, r_411__35_, r_411__34_, r_411__33_, r_411__32_, r_411__31_, r_411__30_, r_411__29_, r_411__28_, r_411__27_, r_411__26_, r_411__25_, r_411__24_, r_411__23_, r_411__22_, r_411__21_, r_411__20_, r_411__19_, r_411__18_, r_411__17_, r_411__16_, r_411__15_, r_411__14_, r_411__13_, r_411__12_, r_411__11_, r_411__10_, r_411__9_, r_411__8_, r_411__7_, r_411__6_, r_411__5_, r_411__4_, r_411__3_, r_411__2_, r_411__1_, r_411__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N821)? data_i : 1'b0;
  assign N820 = sel_i[820];
  assign N821 = N3078;
  assign { r_n_411__63_, r_n_411__62_, r_n_411__61_, r_n_411__60_, r_n_411__59_, r_n_411__58_, r_n_411__57_, r_n_411__56_, r_n_411__55_, r_n_411__54_, r_n_411__53_, r_n_411__52_, r_n_411__51_, r_n_411__50_, r_n_411__49_, r_n_411__48_, r_n_411__47_, r_n_411__46_, r_n_411__45_, r_n_411__44_, r_n_411__43_, r_n_411__42_, r_n_411__41_, r_n_411__40_, r_n_411__39_, r_n_411__38_, r_n_411__37_, r_n_411__36_, r_n_411__35_, r_n_411__34_, r_n_411__33_, r_n_411__32_, r_n_411__31_, r_n_411__30_, r_n_411__29_, r_n_411__28_, r_n_411__27_, r_n_411__26_, r_n_411__25_, r_n_411__24_, r_n_411__23_, r_n_411__22_, r_n_411__21_, r_n_411__20_, r_n_411__19_, r_n_411__18_, r_n_411__17_, r_n_411__16_, r_n_411__15_, r_n_411__14_, r_n_411__13_, r_n_411__12_, r_n_411__11_, r_n_411__10_, r_n_411__9_, r_n_411__8_, r_n_411__7_, r_n_411__6_, r_n_411__5_, r_n_411__4_, r_n_411__3_, r_n_411__2_, r_n_411__1_, r_n_411__0_ } = (N822)? { r_412__63_, r_412__62_, r_412__61_, r_412__60_, r_412__59_, r_412__58_, r_412__57_, r_412__56_, r_412__55_, r_412__54_, r_412__53_, r_412__52_, r_412__51_, r_412__50_, r_412__49_, r_412__48_, r_412__47_, r_412__46_, r_412__45_, r_412__44_, r_412__43_, r_412__42_, r_412__41_, r_412__40_, r_412__39_, r_412__38_, r_412__37_, r_412__36_, r_412__35_, r_412__34_, r_412__33_, r_412__32_, r_412__31_, r_412__30_, r_412__29_, r_412__28_, r_412__27_, r_412__26_, r_412__25_, r_412__24_, r_412__23_, r_412__22_, r_412__21_, r_412__20_, r_412__19_, r_412__18_, r_412__17_, r_412__16_, r_412__15_, r_412__14_, r_412__13_, r_412__12_, r_412__11_, r_412__10_, r_412__9_, r_412__8_, r_412__7_, r_412__6_, r_412__5_, r_412__4_, r_412__3_, r_412__2_, r_412__1_, r_412__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N823)? data_i : 1'b0;
  assign N822 = sel_i[822];
  assign N823 = N3083;
  assign { r_n_412__63_, r_n_412__62_, r_n_412__61_, r_n_412__60_, r_n_412__59_, r_n_412__58_, r_n_412__57_, r_n_412__56_, r_n_412__55_, r_n_412__54_, r_n_412__53_, r_n_412__52_, r_n_412__51_, r_n_412__50_, r_n_412__49_, r_n_412__48_, r_n_412__47_, r_n_412__46_, r_n_412__45_, r_n_412__44_, r_n_412__43_, r_n_412__42_, r_n_412__41_, r_n_412__40_, r_n_412__39_, r_n_412__38_, r_n_412__37_, r_n_412__36_, r_n_412__35_, r_n_412__34_, r_n_412__33_, r_n_412__32_, r_n_412__31_, r_n_412__30_, r_n_412__29_, r_n_412__28_, r_n_412__27_, r_n_412__26_, r_n_412__25_, r_n_412__24_, r_n_412__23_, r_n_412__22_, r_n_412__21_, r_n_412__20_, r_n_412__19_, r_n_412__18_, r_n_412__17_, r_n_412__16_, r_n_412__15_, r_n_412__14_, r_n_412__13_, r_n_412__12_, r_n_412__11_, r_n_412__10_, r_n_412__9_, r_n_412__8_, r_n_412__7_, r_n_412__6_, r_n_412__5_, r_n_412__4_, r_n_412__3_, r_n_412__2_, r_n_412__1_, r_n_412__0_ } = (N824)? { r_413__63_, r_413__62_, r_413__61_, r_413__60_, r_413__59_, r_413__58_, r_413__57_, r_413__56_, r_413__55_, r_413__54_, r_413__53_, r_413__52_, r_413__51_, r_413__50_, r_413__49_, r_413__48_, r_413__47_, r_413__46_, r_413__45_, r_413__44_, r_413__43_, r_413__42_, r_413__41_, r_413__40_, r_413__39_, r_413__38_, r_413__37_, r_413__36_, r_413__35_, r_413__34_, r_413__33_, r_413__32_, r_413__31_, r_413__30_, r_413__29_, r_413__28_, r_413__27_, r_413__26_, r_413__25_, r_413__24_, r_413__23_, r_413__22_, r_413__21_, r_413__20_, r_413__19_, r_413__18_, r_413__17_, r_413__16_, r_413__15_, r_413__14_, r_413__13_, r_413__12_, r_413__11_, r_413__10_, r_413__9_, r_413__8_, r_413__7_, r_413__6_, r_413__5_, r_413__4_, r_413__3_, r_413__2_, r_413__1_, r_413__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N825)? data_i : 1'b0;
  assign N824 = sel_i[824];
  assign N825 = N3088;
  assign { r_n_413__63_, r_n_413__62_, r_n_413__61_, r_n_413__60_, r_n_413__59_, r_n_413__58_, r_n_413__57_, r_n_413__56_, r_n_413__55_, r_n_413__54_, r_n_413__53_, r_n_413__52_, r_n_413__51_, r_n_413__50_, r_n_413__49_, r_n_413__48_, r_n_413__47_, r_n_413__46_, r_n_413__45_, r_n_413__44_, r_n_413__43_, r_n_413__42_, r_n_413__41_, r_n_413__40_, r_n_413__39_, r_n_413__38_, r_n_413__37_, r_n_413__36_, r_n_413__35_, r_n_413__34_, r_n_413__33_, r_n_413__32_, r_n_413__31_, r_n_413__30_, r_n_413__29_, r_n_413__28_, r_n_413__27_, r_n_413__26_, r_n_413__25_, r_n_413__24_, r_n_413__23_, r_n_413__22_, r_n_413__21_, r_n_413__20_, r_n_413__19_, r_n_413__18_, r_n_413__17_, r_n_413__16_, r_n_413__15_, r_n_413__14_, r_n_413__13_, r_n_413__12_, r_n_413__11_, r_n_413__10_, r_n_413__9_, r_n_413__8_, r_n_413__7_, r_n_413__6_, r_n_413__5_, r_n_413__4_, r_n_413__3_, r_n_413__2_, r_n_413__1_, r_n_413__0_ } = (N826)? { r_414__63_, r_414__62_, r_414__61_, r_414__60_, r_414__59_, r_414__58_, r_414__57_, r_414__56_, r_414__55_, r_414__54_, r_414__53_, r_414__52_, r_414__51_, r_414__50_, r_414__49_, r_414__48_, r_414__47_, r_414__46_, r_414__45_, r_414__44_, r_414__43_, r_414__42_, r_414__41_, r_414__40_, r_414__39_, r_414__38_, r_414__37_, r_414__36_, r_414__35_, r_414__34_, r_414__33_, r_414__32_, r_414__31_, r_414__30_, r_414__29_, r_414__28_, r_414__27_, r_414__26_, r_414__25_, r_414__24_, r_414__23_, r_414__22_, r_414__21_, r_414__20_, r_414__19_, r_414__18_, r_414__17_, r_414__16_, r_414__15_, r_414__14_, r_414__13_, r_414__12_, r_414__11_, r_414__10_, r_414__9_, r_414__8_, r_414__7_, r_414__6_, r_414__5_, r_414__4_, r_414__3_, r_414__2_, r_414__1_, r_414__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N827)? data_i : 1'b0;
  assign N826 = sel_i[826];
  assign N827 = N3093;
  assign { r_n_414__63_, r_n_414__62_, r_n_414__61_, r_n_414__60_, r_n_414__59_, r_n_414__58_, r_n_414__57_, r_n_414__56_, r_n_414__55_, r_n_414__54_, r_n_414__53_, r_n_414__52_, r_n_414__51_, r_n_414__50_, r_n_414__49_, r_n_414__48_, r_n_414__47_, r_n_414__46_, r_n_414__45_, r_n_414__44_, r_n_414__43_, r_n_414__42_, r_n_414__41_, r_n_414__40_, r_n_414__39_, r_n_414__38_, r_n_414__37_, r_n_414__36_, r_n_414__35_, r_n_414__34_, r_n_414__33_, r_n_414__32_, r_n_414__31_, r_n_414__30_, r_n_414__29_, r_n_414__28_, r_n_414__27_, r_n_414__26_, r_n_414__25_, r_n_414__24_, r_n_414__23_, r_n_414__22_, r_n_414__21_, r_n_414__20_, r_n_414__19_, r_n_414__18_, r_n_414__17_, r_n_414__16_, r_n_414__15_, r_n_414__14_, r_n_414__13_, r_n_414__12_, r_n_414__11_, r_n_414__10_, r_n_414__9_, r_n_414__8_, r_n_414__7_, r_n_414__6_, r_n_414__5_, r_n_414__4_, r_n_414__3_, r_n_414__2_, r_n_414__1_, r_n_414__0_ } = (N828)? { r_415__63_, r_415__62_, r_415__61_, r_415__60_, r_415__59_, r_415__58_, r_415__57_, r_415__56_, r_415__55_, r_415__54_, r_415__53_, r_415__52_, r_415__51_, r_415__50_, r_415__49_, r_415__48_, r_415__47_, r_415__46_, r_415__45_, r_415__44_, r_415__43_, r_415__42_, r_415__41_, r_415__40_, r_415__39_, r_415__38_, r_415__37_, r_415__36_, r_415__35_, r_415__34_, r_415__33_, r_415__32_, r_415__31_, r_415__30_, r_415__29_, r_415__28_, r_415__27_, r_415__26_, r_415__25_, r_415__24_, r_415__23_, r_415__22_, r_415__21_, r_415__20_, r_415__19_, r_415__18_, r_415__17_, r_415__16_, r_415__15_, r_415__14_, r_415__13_, r_415__12_, r_415__11_, r_415__10_, r_415__9_, r_415__8_, r_415__7_, r_415__6_, r_415__5_, r_415__4_, r_415__3_, r_415__2_, r_415__1_, r_415__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N829)? data_i : 1'b0;
  assign N828 = sel_i[828];
  assign N829 = N3098;
  assign { r_n_415__63_, r_n_415__62_, r_n_415__61_, r_n_415__60_, r_n_415__59_, r_n_415__58_, r_n_415__57_, r_n_415__56_, r_n_415__55_, r_n_415__54_, r_n_415__53_, r_n_415__52_, r_n_415__51_, r_n_415__50_, r_n_415__49_, r_n_415__48_, r_n_415__47_, r_n_415__46_, r_n_415__45_, r_n_415__44_, r_n_415__43_, r_n_415__42_, r_n_415__41_, r_n_415__40_, r_n_415__39_, r_n_415__38_, r_n_415__37_, r_n_415__36_, r_n_415__35_, r_n_415__34_, r_n_415__33_, r_n_415__32_, r_n_415__31_, r_n_415__30_, r_n_415__29_, r_n_415__28_, r_n_415__27_, r_n_415__26_, r_n_415__25_, r_n_415__24_, r_n_415__23_, r_n_415__22_, r_n_415__21_, r_n_415__20_, r_n_415__19_, r_n_415__18_, r_n_415__17_, r_n_415__16_, r_n_415__15_, r_n_415__14_, r_n_415__13_, r_n_415__12_, r_n_415__11_, r_n_415__10_, r_n_415__9_, r_n_415__8_, r_n_415__7_, r_n_415__6_, r_n_415__5_, r_n_415__4_, r_n_415__3_, r_n_415__2_, r_n_415__1_, r_n_415__0_ } = (N830)? { r_416__63_, r_416__62_, r_416__61_, r_416__60_, r_416__59_, r_416__58_, r_416__57_, r_416__56_, r_416__55_, r_416__54_, r_416__53_, r_416__52_, r_416__51_, r_416__50_, r_416__49_, r_416__48_, r_416__47_, r_416__46_, r_416__45_, r_416__44_, r_416__43_, r_416__42_, r_416__41_, r_416__40_, r_416__39_, r_416__38_, r_416__37_, r_416__36_, r_416__35_, r_416__34_, r_416__33_, r_416__32_, r_416__31_, r_416__30_, r_416__29_, r_416__28_, r_416__27_, r_416__26_, r_416__25_, r_416__24_, r_416__23_, r_416__22_, r_416__21_, r_416__20_, r_416__19_, r_416__18_, r_416__17_, r_416__16_, r_416__15_, r_416__14_, r_416__13_, r_416__12_, r_416__11_, r_416__10_, r_416__9_, r_416__8_, r_416__7_, r_416__6_, r_416__5_, r_416__4_, r_416__3_, r_416__2_, r_416__1_, r_416__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N831)? data_i : 1'b0;
  assign N830 = sel_i[830];
  assign N831 = N3103;
  assign { r_n_416__63_, r_n_416__62_, r_n_416__61_, r_n_416__60_, r_n_416__59_, r_n_416__58_, r_n_416__57_, r_n_416__56_, r_n_416__55_, r_n_416__54_, r_n_416__53_, r_n_416__52_, r_n_416__51_, r_n_416__50_, r_n_416__49_, r_n_416__48_, r_n_416__47_, r_n_416__46_, r_n_416__45_, r_n_416__44_, r_n_416__43_, r_n_416__42_, r_n_416__41_, r_n_416__40_, r_n_416__39_, r_n_416__38_, r_n_416__37_, r_n_416__36_, r_n_416__35_, r_n_416__34_, r_n_416__33_, r_n_416__32_, r_n_416__31_, r_n_416__30_, r_n_416__29_, r_n_416__28_, r_n_416__27_, r_n_416__26_, r_n_416__25_, r_n_416__24_, r_n_416__23_, r_n_416__22_, r_n_416__21_, r_n_416__20_, r_n_416__19_, r_n_416__18_, r_n_416__17_, r_n_416__16_, r_n_416__15_, r_n_416__14_, r_n_416__13_, r_n_416__12_, r_n_416__11_, r_n_416__10_, r_n_416__9_, r_n_416__8_, r_n_416__7_, r_n_416__6_, r_n_416__5_, r_n_416__4_, r_n_416__3_, r_n_416__2_, r_n_416__1_, r_n_416__0_ } = (N832)? { r_417__63_, r_417__62_, r_417__61_, r_417__60_, r_417__59_, r_417__58_, r_417__57_, r_417__56_, r_417__55_, r_417__54_, r_417__53_, r_417__52_, r_417__51_, r_417__50_, r_417__49_, r_417__48_, r_417__47_, r_417__46_, r_417__45_, r_417__44_, r_417__43_, r_417__42_, r_417__41_, r_417__40_, r_417__39_, r_417__38_, r_417__37_, r_417__36_, r_417__35_, r_417__34_, r_417__33_, r_417__32_, r_417__31_, r_417__30_, r_417__29_, r_417__28_, r_417__27_, r_417__26_, r_417__25_, r_417__24_, r_417__23_, r_417__22_, r_417__21_, r_417__20_, r_417__19_, r_417__18_, r_417__17_, r_417__16_, r_417__15_, r_417__14_, r_417__13_, r_417__12_, r_417__11_, r_417__10_, r_417__9_, r_417__8_, r_417__7_, r_417__6_, r_417__5_, r_417__4_, r_417__3_, r_417__2_, r_417__1_, r_417__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N833)? data_i : 1'b0;
  assign N832 = sel_i[832];
  assign N833 = N3108;
  assign { r_n_417__63_, r_n_417__62_, r_n_417__61_, r_n_417__60_, r_n_417__59_, r_n_417__58_, r_n_417__57_, r_n_417__56_, r_n_417__55_, r_n_417__54_, r_n_417__53_, r_n_417__52_, r_n_417__51_, r_n_417__50_, r_n_417__49_, r_n_417__48_, r_n_417__47_, r_n_417__46_, r_n_417__45_, r_n_417__44_, r_n_417__43_, r_n_417__42_, r_n_417__41_, r_n_417__40_, r_n_417__39_, r_n_417__38_, r_n_417__37_, r_n_417__36_, r_n_417__35_, r_n_417__34_, r_n_417__33_, r_n_417__32_, r_n_417__31_, r_n_417__30_, r_n_417__29_, r_n_417__28_, r_n_417__27_, r_n_417__26_, r_n_417__25_, r_n_417__24_, r_n_417__23_, r_n_417__22_, r_n_417__21_, r_n_417__20_, r_n_417__19_, r_n_417__18_, r_n_417__17_, r_n_417__16_, r_n_417__15_, r_n_417__14_, r_n_417__13_, r_n_417__12_, r_n_417__11_, r_n_417__10_, r_n_417__9_, r_n_417__8_, r_n_417__7_, r_n_417__6_, r_n_417__5_, r_n_417__4_, r_n_417__3_, r_n_417__2_, r_n_417__1_, r_n_417__0_ } = (N834)? { r_418__63_, r_418__62_, r_418__61_, r_418__60_, r_418__59_, r_418__58_, r_418__57_, r_418__56_, r_418__55_, r_418__54_, r_418__53_, r_418__52_, r_418__51_, r_418__50_, r_418__49_, r_418__48_, r_418__47_, r_418__46_, r_418__45_, r_418__44_, r_418__43_, r_418__42_, r_418__41_, r_418__40_, r_418__39_, r_418__38_, r_418__37_, r_418__36_, r_418__35_, r_418__34_, r_418__33_, r_418__32_, r_418__31_, r_418__30_, r_418__29_, r_418__28_, r_418__27_, r_418__26_, r_418__25_, r_418__24_, r_418__23_, r_418__22_, r_418__21_, r_418__20_, r_418__19_, r_418__18_, r_418__17_, r_418__16_, r_418__15_, r_418__14_, r_418__13_, r_418__12_, r_418__11_, r_418__10_, r_418__9_, r_418__8_, r_418__7_, r_418__6_, r_418__5_, r_418__4_, r_418__3_, r_418__2_, r_418__1_, r_418__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N835)? data_i : 1'b0;
  assign N834 = sel_i[834];
  assign N835 = N3113;
  assign { r_n_418__63_, r_n_418__62_, r_n_418__61_, r_n_418__60_, r_n_418__59_, r_n_418__58_, r_n_418__57_, r_n_418__56_, r_n_418__55_, r_n_418__54_, r_n_418__53_, r_n_418__52_, r_n_418__51_, r_n_418__50_, r_n_418__49_, r_n_418__48_, r_n_418__47_, r_n_418__46_, r_n_418__45_, r_n_418__44_, r_n_418__43_, r_n_418__42_, r_n_418__41_, r_n_418__40_, r_n_418__39_, r_n_418__38_, r_n_418__37_, r_n_418__36_, r_n_418__35_, r_n_418__34_, r_n_418__33_, r_n_418__32_, r_n_418__31_, r_n_418__30_, r_n_418__29_, r_n_418__28_, r_n_418__27_, r_n_418__26_, r_n_418__25_, r_n_418__24_, r_n_418__23_, r_n_418__22_, r_n_418__21_, r_n_418__20_, r_n_418__19_, r_n_418__18_, r_n_418__17_, r_n_418__16_, r_n_418__15_, r_n_418__14_, r_n_418__13_, r_n_418__12_, r_n_418__11_, r_n_418__10_, r_n_418__9_, r_n_418__8_, r_n_418__7_, r_n_418__6_, r_n_418__5_, r_n_418__4_, r_n_418__3_, r_n_418__2_, r_n_418__1_, r_n_418__0_ } = (N836)? { r_419__63_, r_419__62_, r_419__61_, r_419__60_, r_419__59_, r_419__58_, r_419__57_, r_419__56_, r_419__55_, r_419__54_, r_419__53_, r_419__52_, r_419__51_, r_419__50_, r_419__49_, r_419__48_, r_419__47_, r_419__46_, r_419__45_, r_419__44_, r_419__43_, r_419__42_, r_419__41_, r_419__40_, r_419__39_, r_419__38_, r_419__37_, r_419__36_, r_419__35_, r_419__34_, r_419__33_, r_419__32_, r_419__31_, r_419__30_, r_419__29_, r_419__28_, r_419__27_, r_419__26_, r_419__25_, r_419__24_, r_419__23_, r_419__22_, r_419__21_, r_419__20_, r_419__19_, r_419__18_, r_419__17_, r_419__16_, r_419__15_, r_419__14_, r_419__13_, r_419__12_, r_419__11_, r_419__10_, r_419__9_, r_419__8_, r_419__7_, r_419__6_, r_419__5_, r_419__4_, r_419__3_, r_419__2_, r_419__1_, r_419__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N837)? data_i : 1'b0;
  assign N836 = sel_i[836];
  assign N837 = N3118;
  assign { r_n_419__63_, r_n_419__62_, r_n_419__61_, r_n_419__60_, r_n_419__59_, r_n_419__58_, r_n_419__57_, r_n_419__56_, r_n_419__55_, r_n_419__54_, r_n_419__53_, r_n_419__52_, r_n_419__51_, r_n_419__50_, r_n_419__49_, r_n_419__48_, r_n_419__47_, r_n_419__46_, r_n_419__45_, r_n_419__44_, r_n_419__43_, r_n_419__42_, r_n_419__41_, r_n_419__40_, r_n_419__39_, r_n_419__38_, r_n_419__37_, r_n_419__36_, r_n_419__35_, r_n_419__34_, r_n_419__33_, r_n_419__32_, r_n_419__31_, r_n_419__30_, r_n_419__29_, r_n_419__28_, r_n_419__27_, r_n_419__26_, r_n_419__25_, r_n_419__24_, r_n_419__23_, r_n_419__22_, r_n_419__21_, r_n_419__20_, r_n_419__19_, r_n_419__18_, r_n_419__17_, r_n_419__16_, r_n_419__15_, r_n_419__14_, r_n_419__13_, r_n_419__12_, r_n_419__11_, r_n_419__10_, r_n_419__9_, r_n_419__8_, r_n_419__7_, r_n_419__6_, r_n_419__5_, r_n_419__4_, r_n_419__3_, r_n_419__2_, r_n_419__1_, r_n_419__0_ } = (N838)? { r_420__63_, r_420__62_, r_420__61_, r_420__60_, r_420__59_, r_420__58_, r_420__57_, r_420__56_, r_420__55_, r_420__54_, r_420__53_, r_420__52_, r_420__51_, r_420__50_, r_420__49_, r_420__48_, r_420__47_, r_420__46_, r_420__45_, r_420__44_, r_420__43_, r_420__42_, r_420__41_, r_420__40_, r_420__39_, r_420__38_, r_420__37_, r_420__36_, r_420__35_, r_420__34_, r_420__33_, r_420__32_, r_420__31_, r_420__30_, r_420__29_, r_420__28_, r_420__27_, r_420__26_, r_420__25_, r_420__24_, r_420__23_, r_420__22_, r_420__21_, r_420__20_, r_420__19_, r_420__18_, r_420__17_, r_420__16_, r_420__15_, r_420__14_, r_420__13_, r_420__12_, r_420__11_, r_420__10_, r_420__9_, r_420__8_, r_420__7_, r_420__6_, r_420__5_, r_420__4_, r_420__3_, r_420__2_, r_420__1_, r_420__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N839)? data_i : 1'b0;
  assign N838 = sel_i[838];
  assign N839 = N3123;
  assign { r_n_420__63_, r_n_420__62_, r_n_420__61_, r_n_420__60_, r_n_420__59_, r_n_420__58_, r_n_420__57_, r_n_420__56_, r_n_420__55_, r_n_420__54_, r_n_420__53_, r_n_420__52_, r_n_420__51_, r_n_420__50_, r_n_420__49_, r_n_420__48_, r_n_420__47_, r_n_420__46_, r_n_420__45_, r_n_420__44_, r_n_420__43_, r_n_420__42_, r_n_420__41_, r_n_420__40_, r_n_420__39_, r_n_420__38_, r_n_420__37_, r_n_420__36_, r_n_420__35_, r_n_420__34_, r_n_420__33_, r_n_420__32_, r_n_420__31_, r_n_420__30_, r_n_420__29_, r_n_420__28_, r_n_420__27_, r_n_420__26_, r_n_420__25_, r_n_420__24_, r_n_420__23_, r_n_420__22_, r_n_420__21_, r_n_420__20_, r_n_420__19_, r_n_420__18_, r_n_420__17_, r_n_420__16_, r_n_420__15_, r_n_420__14_, r_n_420__13_, r_n_420__12_, r_n_420__11_, r_n_420__10_, r_n_420__9_, r_n_420__8_, r_n_420__7_, r_n_420__6_, r_n_420__5_, r_n_420__4_, r_n_420__3_, r_n_420__2_, r_n_420__1_, r_n_420__0_ } = (N840)? { r_421__63_, r_421__62_, r_421__61_, r_421__60_, r_421__59_, r_421__58_, r_421__57_, r_421__56_, r_421__55_, r_421__54_, r_421__53_, r_421__52_, r_421__51_, r_421__50_, r_421__49_, r_421__48_, r_421__47_, r_421__46_, r_421__45_, r_421__44_, r_421__43_, r_421__42_, r_421__41_, r_421__40_, r_421__39_, r_421__38_, r_421__37_, r_421__36_, r_421__35_, r_421__34_, r_421__33_, r_421__32_, r_421__31_, r_421__30_, r_421__29_, r_421__28_, r_421__27_, r_421__26_, r_421__25_, r_421__24_, r_421__23_, r_421__22_, r_421__21_, r_421__20_, r_421__19_, r_421__18_, r_421__17_, r_421__16_, r_421__15_, r_421__14_, r_421__13_, r_421__12_, r_421__11_, r_421__10_, r_421__9_, r_421__8_, r_421__7_, r_421__6_, r_421__5_, r_421__4_, r_421__3_, r_421__2_, r_421__1_, r_421__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N841)? data_i : 1'b0;
  assign N840 = sel_i[840];
  assign N841 = N3128;
  assign { r_n_421__63_, r_n_421__62_, r_n_421__61_, r_n_421__60_, r_n_421__59_, r_n_421__58_, r_n_421__57_, r_n_421__56_, r_n_421__55_, r_n_421__54_, r_n_421__53_, r_n_421__52_, r_n_421__51_, r_n_421__50_, r_n_421__49_, r_n_421__48_, r_n_421__47_, r_n_421__46_, r_n_421__45_, r_n_421__44_, r_n_421__43_, r_n_421__42_, r_n_421__41_, r_n_421__40_, r_n_421__39_, r_n_421__38_, r_n_421__37_, r_n_421__36_, r_n_421__35_, r_n_421__34_, r_n_421__33_, r_n_421__32_, r_n_421__31_, r_n_421__30_, r_n_421__29_, r_n_421__28_, r_n_421__27_, r_n_421__26_, r_n_421__25_, r_n_421__24_, r_n_421__23_, r_n_421__22_, r_n_421__21_, r_n_421__20_, r_n_421__19_, r_n_421__18_, r_n_421__17_, r_n_421__16_, r_n_421__15_, r_n_421__14_, r_n_421__13_, r_n_421__12_, r_n_421__11_, r_n_421__10_, r_n_421__9_, r_n_421__8_, r_n_421__7_, r_n_421__6_, r_n_421__5_, r_n_421__4_, r_n_421__3_, r_n_421__2_, r_n_421__1_, r_n_421__0_ } = (N842)? { r_422__63_, r_422__62_, r_422__61_, r_422__60_, r_422__59_, r_422__58_, r_422__57_, r_422__56_, r_422__55_, r_422__54_, r_422__53_, r_422__52_, r_422__51_, r_422__50_, r_422__49_, r_422__48_, r_422__47_, r_422__46_, r_422__45_, r_422__44_, r_422__43_, r_422__42_, r_422__41_, r_422__40_, r_422__39_, r_422__38_, r_422__37_, r_422__36_, r_422__35_, r_422__34_, r_422__33_, r_422__32_, r_422__31_, r_422__30_, r_422__29_, r_422__28_, r_422__27_, r_422__26_, r_422__25_, r_422__24_, r_422__23_, r_422__22_, r_422__21_, r_422__20_, r_422__19_, r_422__18_, r_422__17_, r_422__16_, r_422__15_, r_422__14_, r_422__13_, r_422__12_, r_422__11_, r_422__10_, r_422__9_, r_422__8_, r_422__7_, r_422__6_, r_422__5_, r_422__4_, r_422__3_, r_422__2_, r_422__1_, r_422__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N843)? data_i : 1'b0;
  assign N842 = sel_i[842];
  assign N843 = N3133;
  assign { r_n_422__63_, r_n_422__62_, r_n_422__61_, r_n_422__60_, r_n_422__59_, r_n_422__58_, r_n_422__57_, r_n_422__56_, r_n_422__55_, r_n_422__54_, r_n_422__53_, r_n_422__52_, r_n_422__51_, r_n_422__50_, r_n_422__49_, r_n_422__48_, r_n_422__47_, r_n_422__46_, r_n_422__45_, r_n_422__44_, r_n_422__43_, r_n_422__42_, r_n_422__41_, r_n_422__40_, r_n_422__39_, r_n_422__38_, r_n_422__37_, r_n_422__36_, r_n_422__35_, r_n_422__34_, r_n_422__33_, r_n_422__32_, r_n_422__31_, r_n_422__30_, r_n_422__29_, r_n_422__28_, r_n_422__27_, r_n_422__26_, r_n_422__25_, r_n_422__24_, r_n_422__23_, r_n_422__22_, r_n_422__21_, r_n_422__20_, r_n_422__19_, r_n_422__18_, r_n_422__17_, r_n_422__16_, r_n_422__15_, r_n_422__14_, r_n_422__13_, r_n_422__12_, r_n_422__11_, r_n_422__10_, r_n_422__9_, r_n_422__8_, r_n_422__7_, r_n_422__6_, r_n_422__5_, r_n_422__4_, r_n_422__3_, r_n_422__2_, r_n_422__1_, r_n_422__0_ } = (N844)? { r_423__63_, r_423__62_, r_423__61_, r_423__60_, r_423__59_, r_423__58_, r_423__57_, r_423__56_, r_423__55_, r_423__54_, r_423__53_, r_423__52_, r_423__51_, r_423__50_, r_423__49_, r_423__48_, r_423__47_, r_423__46_, r_423__45_, r_423__44_, r_423__43_, r_423__42_, r_423__41_, r_423__40_, r_423__39_, r_423__38_, r_423__37_, r_423__36_, r_423__35_, r_423__34_, r_423__33_, r_423__32_, r_423__31_, r_423__30_, r_423__29_, r_423__28_, r_423__27_, r_423__26_, r_423__25_, r_423__24_, r_423__23_, r_423__22_, r_423__21_, r_423__20_, r_423__19_, r_423__18_, r_423__17_, r_423__16_, r_423__15_, r_423__14_, r_423__13_, r_423__12_, r_423__11_, r_423__10_, r_423__9_, r_423__8_, r_423__7_, r_423__6_, r_423__5_, r_423__4_, r_423__3_, r_423__2_, r_423__1_, r_423__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N845)? data_i : 1'b0;
  assign N844 = sel_i[844];
  assign N845 = N3138;
  assign { r_n_423__63_, r_n_423__62_, r_n_423__61_, r_n_423__60_, r_n_423__59_, r_n_423__58_, r_n_423__57_, r_n_423__56_, r_n_423__55_, r_n_423__54_, r_n_423__53_, r_n_423__52_, r_n_423__51_, r_n_423__50_, r_n_423__49_, r_n_423__48_, r_n_423__47_, r_n_423__46_, r_n_423__45_, r_n_423__44_, r_n_423__43_, r_n_423__42_, r_n_423__41_, r_n_423__40_, r_n_423__39_, r_n_423__38_, r_n_423__37_, r_n_423__36_, r_n_423__35_, r_n_423__34_, r_n_423__33_, r_n_423__32_, r_n_423__31_, r_n_423__30_, r_n_423__29_, r_n_423__28_, r_n_423__27_, r_n_423__26_, r_n_423__25_, r_n_423__24_, r_n_423__23_, r_n_423__22_, r_n_423__21_, r_n_423__20_, r_n_423__19_, r_n_423__18_, r_n_423__17_, r_n_423__16_, r_n_423__15_, r_n_423__14_, r_n_423__13_, r_n_423__12_, r_n_423__11_, r_n_423__10_, r_n_423__9_, r_n_423__8_, r_n_423__7_, r_n_423__6_, r_n_423__5_, r_n_423__4_, r_n_423__3_, r_n_423__2_, r_n_423__1_, r_n_423__0_ } = (N846)? { r_424__63_, r_424__62_, r_424__61_, r_424__60_, r_424__59_, r_424__58_, r_424__57_, r_424__56_, r_424__55_, r_424__54_, r_424__53_, r_424__52_, r_424__51_, r_424__50_, r_424__49_, r_424__48_, r_424__47_, r_424__46_, r_424__45_, r_424__44_, r_424__43_, r_424__42_, r_424__41_, r_424__40_, r_424__39_, r_424__38_, r_424__37_, r_424__36_, r_424__35_, r_424__34_, r_424__33_, r_424__32_, r_424__31_, r_424__30_, r_424__29_, r_424__28_, r_424__27_, r_424__26_, r_424__25_, r_424__24_, r_424__23_, r_424__22_, r_424__21_, r_424__20_, r_424__19_, r_424__18_, r_424__17_, r_424__16_, r_424__15_, r_424__14_, r_424__13_, r_424__12_, r_424__11_, r_424__10_, r_424__9_, r_424__8_, r_424__7_, r_424__6_, r_424__5_, r_424__4_, r_424__3_, r_424__2_, r_424__1_, r_424__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N847)? data_i : 1'b0;
  assign N846 = sel_i[846];
  assign N847 = N3143;
  assign { r_n_424__63_, r_n_424__62_, r_n_424__61_, r_n_424__60_, r_n_424__59_, r_n_424__58_, r_n_424__57_, r_n_424__56_, r_n_424__55_, r_n_424__54_, r_n_424__53_, r_n_424__52_, r_n_424__51_, r_n_424__50_, r_n_424__49_, r_n_424__48_, r_n_424__47_, r_n_424__46_, r_n_424__45_, r_n_424__44_, r_n_424__43_, r_n_424__42_, r_n_424__41_, r_n_424__40_, r_n_424__39_, r_n_424__38_, r_n_424__37_, r_n_424__36_, r_n_424__35_, r_n_424__34_, r_n_424__33_, r_n_424__32_, r_n_424__31_, r_n_424__30_, r_n_424__29_, r_n_424__28_, r_n_424__27_, r_n_424__26_, r_n_424__25_, r_n_424__24_, r_n_424__23_, r_n_424__22_, r_n_424__21_, r_n_424__20_, r_n_424__19_, r_n_424__18_, r_n_424__17_, r_n_424__16_, r_n_424__15_, r_n_424__14_, r_n_424__13_, r_n_424__12_, r_n_424__11_, r_n_424__10_, r_n_424__9_, r_n_424__8_, r_n_424__7_, r_n_424__6_, r_n_424__5_, r_n_424__4_, r_n_424__3_, r_n_424__2_, r_n_424__1_, r_n_424__0_ } = (N848)? { r_425__63_, r_425__62_, r_425__61_, r_425__60_, r_425__59_, r_425__58_, r_425__57_, r_425__56_, r_425__55_, r_425__54_, r_425__53_, r_425__52_, r_425__51_, r_425__50_, r_425__49_, r_425__48_, r_425__47_, r_425__46_, r_425__45_, r_425__44_, r_425__43_, r_425__42_, r_425__41_, r_425__40_, r_425__39_, r_425__38_, r_425__37_, r_425__36_, r_425__35_, r_425__34_, r_425__33_, r_425__32_, r_425__31_, r_425__30_, r_425__29_, r_425__28_, r_425__27_, r_425__26_, r_425__25_, r_425__24_, r_425__23_, r_425__22_, r_425__21_, r_425__20_, r_425__19_, r_425__18_, r_425__17_, r_425__16_, r_425__15_, r_425__14_, r_425__13_, r_425__12_, r_425__11_, r_425__10_, r_425__9_, r_425__8_, r_425__7_, r_425__6_, r_425__5_, r_425__4_, r_425__3_, r_425__2_, r_425__1_, r_425__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N849)? data_i : 1'b0;
  assign N848 = sel_i[848];
  assign N849 = N3148;
  assign { r_n_425__63_, r_n_425__62_, r_n_425__61_, r_n_425__60_, r_n_425__59_, r_n_425__58_, r_n_425__57_, r_n_425__56_, r_n_425__55_, r_n_425__54_, r_n_425__53_, r_n_425__52_, r_n_425__51_, r_n_425__50_, r_n_425__49_, r_n_425__48_, r_n_425__47_, r_n_425__46_, r_n_425__45_, r_n_425__44_, r_n_425__43_, r_n_425__42_, r_n_425__41_, r_n_425__40_, r_n_425__39_, r_n_425__38_, r_n_425__37_, r_n_425__36_, r_n_425__35_, r_n_425__34_, r_n_425__33_, r_n_425__32_, r_n_425__31_, r_n_425__30_, r_n_425__29_, r_n_425__28_, r_n_425__27_, r_n_425__26_, r_n_425__25_, r_n_425__24_, r_n_425__23_, r_n_425__22_, r_n_425__21_, r_n_425__20_, r_n_425__19_, r_n_425__18_, r_n_425__17_, r_n_425__16_, r_n_425__15_, r_n_425__14_, r_n_425__13_, r_n_425__12_, r_n_425__11_, r_n_425__10_, r_n_425__9_, r_n_425__8_, r_n_425__7_, r_n_425__6_, r_n_425__5_, r_n_425__4_, r_n_425__3_, r_n_425__2_, r_n_425__1_, r_n_425__0_ } = (N850)? { r_426__63_, r_426__62_, r_426__61_, r_426__60_, r_426__59_, r_426__58_, r_426__57_, r_426__56_, r_426__55_, r_426__54_, r_426__53_, r_426__52_, r_426__51_, r_426__50_, r_426__49_, r_426__48_, r_426__47_, r_426__46_, r_426__45_, r_426__44_, r_426__43_, r_426__42_, r_426__41_, r_426__40_, r_426__39_, r_426__38_, r_426__37_, r_426__36_, r_426__35_, r_426__34_, r_426__33_, r_426__32_, r_426__31_, r_426__30_, r_426__29_, r_426__28_, r_426__27_, r_426__26_, r_426__25_, r_426__24_, r_426__23_, r_426__22_, r_426__21_, r_426__20_, r_426__19_, r_426__18_, r_426__17_, r_426__16_, r_426__15_, r_426__14_, r_426__13_, r_426__12_, r_426__11_, r_426__10_, r_426__9_, r_426__8_, r_426__7_, r_426__6_, r_426__5_, r_426__4_, r_426__3_, r_426__2_, r_426__1_, r_426__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N851)? data_i : 1'b0;
  assign N850 = sel_i[850];
  assign N851 = N3153;
  assign { r_n_426__63_, r_n_426__62_, r_n_426__61_, r_n_426__60_, r_n_426__59_, r_n_426__58_, r_n_426__57_, r_n_426__56_, r_n_426__55_, r_n_426__54_, r_n_426__53_, r_n_426__52_, r_n_426__51_, r_n_426__50_, r_n_426__49_, r_n_426__48_, r_n_426__47_, r_n_426__46_, r_n_426__45_, r_n_426__44_, r_n_426__43_, r_n_426__42_, r_n_426__41_, r_n_426__40_, r_n_426__39_, r_n_426__38_, r_n_426__37_, r_n_426__36_, r_n_426__35_, r_n_426__34_, r_n_426__33_, r_n_426__32_, r_n_426__31_, r_n_426__30_, r_n_426__29_, r_n_426__28_, r_n_426__27_, r_n_426__26_, r_n_426__25_, r_n_426__24_, r_n_426__23_, r_n_426__22_, r_n_426__21_, r_n_426__20_, r_n_426__19_, r_n_426__18_, r_n_426__17_, r_n_426__16_, r_n_426__15_, r_n_426__14_, r_n_426__13_, r_n_426__12_, r_n_426__11_, r_n_426__10_, r_n_426__9_, r_n_426__8_, r_n_426__7_, r_n_426__6_, r_n_426__5_, r_n_426__4_, r_n_426__3_, r_n_426__2_, r_n_426__1_, r_n_426__0_ } = (N852)? { r_427__63_, r_427__62_, r_427__61_, r_427__60_, r_427__59_, r_427__58_, r_427__57_, r_427__56_, r_427__55_, r_427__54_, r_427__53_, r_427__52_, r_427__51_, r_427__50_, r_427__49_, r_427__48_, r_427__47_, r_427__46_, r_427__45_, r_427__44_, r_427__43_, r_427__42_, r_427__41_, r_427__40_, r_427__39_, r_427__38_, r_427__37_, r_427__36_, r_427__35_, r_427__34_, r_427__33_, r_427__32_, r_427__31_, r_427__30_, r_427__29_, r_427__28_, r_427__27_, r_427__26_, r_427__25_, r_427__24_, r_427__23_, r_427__22_, r_427__21_, r_427__20_, r_427__19_, r_427__18_, r_427__17_, r_427__16_, r_427__15_, r_427__14_, r_427__13_, r_427__12_, r_427__11_, r_427__10_, r_427__9_, r_427__8_, r_427__7_, r_427__6_, r_427__5_, r_427__4_, r_427__3_, r_427__2_, r_427__1_, r_427__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N853)? data_i : 1'b0;
  assign N852 = sel_i[852];
  assign N853 = N3158;
  assign { r_n_427__63_, r_n_427__62_, r_n_427__61_, r_n_427__60_, r_n_427__59_, r_n_427__58_, r_n_427__57_, r_n_427__56_, r_n_427__55_, r_n_427__54_, r_n_427__53_, r_n_427__52_, r_n_427__51_, r_n_427__50_, r_n_427__49_, r_n_427__48_, r_n_427__47_, r_n_427__46_, r_n_427__45_, r_n_427__44_, r_n_427__43_, r_n_427__42_, r_n_427__41_, r_n_427__40_, r_n_427__39_, r_n_427__38_, r_n_427__37_, r_n_427__36_, r_n_427__35_, r_n_427__34_, r_n_427__33_, r_n_427__32_, r_n_427__31_, r_n_427__30_, r_n_427__29_, r_n_427__28_, r_n_427__27_, r_n_427__26_, r_n_427__25_, r_n_427__24_, r_n_427__23_, r_n_427__22_, r_n_427__21_, r_n_427__20_, r_n_427__19_, r_n_427__18_, r_n_427__17_, r_n_427__16_, r_n_427__15_, r_n_427__14_, r_n_427__13_, r_n_427__12_, r_n_427__11_, r_n_427__10_, r_n_427__9_, r_n_427__8_, r_n_427__7_, r_n_427__6_, r_n_427__5_, r_n_427__4_, r_n_427__3_, r_n_427__2_, r_n_427__1_, r_n_427__0_ } = (N854)? { r_428__63_, r_428__62_, r_428__61_, r_428__60_, r_428__59_, r_428__58_, r_428__57_, r_428__56_, r_428__55_, r_428__54_, r_428__53_, r_428__52_, r_428__51_, r_428__50_, r_428__49_, r_428__48_, r_428__47_, r_428__46_, r_428__45_, r_428__44_, r_428__43_, r_428__42_, r_428__41_, r_428__40_, r_428__39_, r_428__38_, r_428__37_, r_428__36_, r_428__35_, r_428__34_, r_428__33_, r_428__32_, r_428__31_, r_428__30_, r_428__29_, r_428__28_, r_428__27_, r_428__26_, r_428__25_, r_428__24_, r_428__23_, r_428__22_, r_428__21_, r_428__20_, r_428__19_, r_428__18_, r_428__17_, r_428__16_, r_428__15_, r_428__14_, r_428__13_, r_428__12_, r_428__11_, r_428__10_, r_428__9_, r_428__8_, r_428__7_, r_428__6_, r_428__5_, r_428__4_, r_428__3_, r_428__2_, r_428__1_, r_428__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N855)? data_i : 1'b0;
  assign N854 = sel_i[854];
  assign N855 = N3163;
  assign { r_n_428__63_, r_n_428__62_, r_n_428__61_, r_n_428__60_, r_n_428__59_, r_n_428__58_, r_n_428__57_, r_n_428__56_, r_n_428__55_, r_n_428__54_, r_n_428__53_, r_n_428__52_, r_n_428__51_, r_n_428__50_, r_n_428__49_, r_n_428__48_, r_n_428__47_, r_n_428__46_, r_n_428__45_, r_n_428__44_, r_n_428__43_, r_n_428__42_, r_n_428__41_, r_n_428__40_, r_n_428__39_, r_n_428__38_, r_n_428__37_, r_n_428__36_, r_n_428__35_, r_n_428__34_, r_n_428__33_, r_n_428__32_, r_n_428__31_, r_n_428__30_, r_n_428__29_, r_n_428__28_, r_n_428__27_, r_n_428__26_, r_n_428__25_, r_n_428__24_, r_n_428__23_, r_n_428__22_, r_n_428__21_, r_n_428__20_, r_n_428__19_, r_n_428__18_, r_n_428__17_, r_n_428__16_, r_n_428__15_, r_n_428__14_, r_n_428__13_, r_n_428__12_, r_n_428__11_, r_n_428__10_, r_n_428__9_, r_n_428__8_, r_n_428__7_, r_n_428__6_, r_n_428__5_, r_n_428__4_, r_n_428__3_, r_n_428__2_, r_n_428__1_, r_n_428__0_ } = (N856)? { r_429__63_, r_429__62_, r_429__61_, r_429__60_, r_429__59_, r_429__58_, r_429__57_, r_429__56_, r_429__55_, r_429__54_, r_429__53_, r_429__52_, r_429__51_, r_429__50_, r_429__49_, r_429__48_, r_429__47_, r_429__46_, r_429__45_, r_429__44_, r_429__43_, r_429__42_, r_429__41_, r_429__40_, r_429__39_, r_429__38_, r_429__37_, r_429__36_, r_429__35_, r_429__34_, r_429__33_, r_429__32_, r_429__31_, r_429__30_, r_429__29_, r_429__28_, r_429__27_, r_429__26_, r_429__25_, r_429__24_, r_429__23_, r_429__22_, r_429__21_, r_429__20_, r_429__19_, r_429__18_, r_429__17_, r_429__16_, r_429__15_, r_429__14_, r_429__13_, r_429__12_, r_429__11_, r_429__10_, r_429__9_, r_429__8_, r_429__7_, r_429__6_, r_429__5_, r_429__4_, r_429__3_, r_429__2_, r_429__1_, r_429__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N857)? data_i : 1'b0;
  assign N856 = sel_i[856];
  assign N857 = N3168;
  assign { r_n_429__63_, r_n_429__62_, r_n_429__61_, r_n_429__60_, r_n_429__59_, r_n_429__58_, r_n_429__57_, r_n_429__56_, r_n_429__55_, r_n_429__54_, r_n_429__53_, r_n_429__52_, r_n_429__51_, r_n_429__50_, r_n_429__49_, r_n_429__48_, r_n_429__47_, r_n_429__46_, r_n_429__45_, r_n_429__44_, r_n_429__43_, r_n_429__42_, r_n_429__41_, r_n_429__40_, r_n_429__39_, r_n_429__38_, r_n_429__37_, r_n_429__36_, r_n_429__35_, r_n_429__34_, r_n_429__33_, r_n_429__32_, r_n_429__31_, r_n_429__30_, r_n_429__29_, r_n_429__28_, r_n_429__27_, r_n_429__26_, r_n_429__25_, r_n_429__24_, r_n_429__23_, r_n_429__22_, r_n_429__21_, r_n_429__20_, r_n_429__19_, r_n_429__18_, r_n_429__17_, r_n_429__16_, r_n_429__15_, r_n_429__14_, r_n_429__13_, r_n_429__12_, r_n_429__11_, r_n_429__10_, r_n_429__9_, r_n_429__8_, r_n_429__7_, r_n_429__6_, r_n_429__5_, r_n_429__4_, r_n_429__3_, r_n_429__2_, r_n_429__1_, r_n_429__0_ } = (N858)? { r_430__63_, r_430__62_, r_430__61_, r_430__60_, r_430__59_, r_430__58_, r_430__57_, r_430__56_, r_430__55_, r_430__54_, r_430__53_, r_430__52_, r_430__51_, r_430__50_, r_430__49_, r_430__48_, r_430__47_, r_430__46_, r_430__45_, r_430__44_, r_430__43_, r_430__42_, r_430__41_, r_430__40_, r_430__39_, r_430__38_, r_430__37_, r_430__36_, r_430__35_, r_430__34_, r_430__33_, r_430__32_, r_430__31_, r_430__30_, r_430__29_, r_430__28_, r_430__27_, r_430__26_, r_430__25_, r_430__24_, r_430__23_, r_430__22_, r_430__21_, r_430__20_, r_430__19_, r_430__18_, r_430__17_, r_430__16_, r_430__15_, r_430__14_, r_430__13_, r_430__12_, r_430__11_, r_430__10_, r_430__9_, r_430__8_, r_430__7_, r_430__6_, r_430__5_, r_430__4_, r_430__3_, r_430__2_, r_430__1_, r_430__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N859)? data_i : 1'b0;
  assign N858 = sel_i[858];
  assign N859 = N3173;
  assign { r_n_430__63_, r_n_430__62_, r_n_430__61_, r_n_430__60_, r_n_430__59_, r_n_430__58_, r_n_430__57_, r_n_430__56_, r_n_430__55_, r_n_430__54_, r_n_430__53_, r_n_430__52_, r_n_430__51_, r_n_430__50_, r_n_430__49_, r_n_430__48_, r_n_430__47_, r_n_430__46_, r_n_430__45_, r_n_430__44_, r_n_430__43_, r_n_430__42_, r_n_430__41_, r_n_430__40_, r_n_430__39_, r_n_430__38_, r_n_430__37_, r_n_430__36_, r_n_430__35_, r_n_430__34_, r_n_430__33_, r_n_430__32_, r_n_430__31_, r_n_430__30_, r_n_430__29_, r_n_430__28_, r_n_430__27_, r_n_430__26_, r_n_430__25_, r_n_430__24_, r_n_430__23_, r_n_430__22_, r_n_430__21_, r_n_430__20_, r_n_430__19_, r_n_430__18_, r_n_430__17_, r_n_430__16_, r_n_430__15_, r_n_430__14_, r_n_430__13_, r_n_430__12_, r_n_430__11_, r_n_430__10_, r_n_430__9_, r_n_430__8_, r_n_430__7_, r_n_430__6_, r_n_430__5_, r_n_430__4_, r_n_430__3_, r_n_430__2_, r_n_430__1_, r_n_430__0_ } = (N860)? { r_431__63_, r_431__62_, r_431__61_, r_431__60_, r_431__59_, r_431__58_, r_431__57_, r_431__56_, r_431__55_, r_431__54_, r_431__53_, r_431__52_, r_431__51_, r_431__50_, r_431__49_, r_431__48_, r_431__47_, r_431__46_, r_431__45_, r_431__44_, r_431__43_, r_431__42_, r_431__41_, r_431__40_, r_431__39_, r_431__38_, r_431__37_, r_431__36_, r_431__35_, r_431__34_, r_431__33_, r_431__32_, r_431__31_, r_431__30_, r_431__29_, r_431__28_, r_431__27_, r_431__26_, r_431__25_, r_431__24_, r_431__23_, r_431__22_, r_431__21_, r_431__20_, r_431__19_, r_431__18_, r_431__17_, r_431__16_, r_431__15_, r_431__14_, r_431__13_, r_431__12_, r_431__11_, r_431__10_, r_431__9_, r_431__8_, r_431__7_, r_431__6_, r_431__5_, r_431__4_, r_431__3_, r_431__2_, r_431__1_, r_431__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N861)? data_i : 1'b0;
  assign N860 = sel_i[860];
  assign N861 = N3178;
  assign { r_n_431__63_, r_n_431__62_, r_n_431__61_, r_n_431__60_, r_n_431__59_, r_n_431__58_, r_n_431__57_, r_n_431__56_, r_n_431__55_, r_n_431__54_, r_n_431__53_, r_n_431__52_, r_n_431__51_, r_n_431__50_, r_n_431__49_, r_n_431__48_, r_n_431__47_, r_n_431__46_, r_n_431__45_, r_n_431__44_, r_n_431__43_, r_n_431__42_, r_n_431__41_, r_n_431__40_, r_n_431__39_, r_n_431__38_, r_n_431__37_, r_n_431__36_, r_n_431__35_, r_n_431__34_, r_n_431__33_, r_n_431__32_, r_n_431__31_, r_n_431__30_, r_n_431__29_, r_n_431__28_, r_n_431__27_, r_n_431__26_, r_n_431__25_, r_n_431__24_, r_n_431__23_, r_n_431__22_, r_n_431__21_, r_n_431__20_, r_n_431__19_, r_n_431__18_, r_n_431__17_, r_n_431__16_, r_n_431__15_, r_n_431__14_, r_n_431__13_, r_n_431__12_, r_n_431__11_, r_n_431__10_, r_n_431__9_, r_n_431__8_, r_n_431__7_, r_n_431__6_, r_n_431__5_, r_n_431__4_, r_n_431__3_, r_n_431__2_, r_n_431__1_, r_n_431__0_ } = (N862)? { r_432__63_, r_432__62_, r_432__61_, r_432__60_, r_432__59_, r_432__58_, r_432__57_, r_432__56_, r_432__55_, r_432__54_, r_432__53_, r_432__52_, r_432__51_, r_432__50_, r_432__49_, r_432__48_, r_432__47_, r_432__46_, r_432__45_, r_432__44_, r_432__43_, r_432__42_, r_432__41_, r_432__40_, r_432__39_, r_432__38_, r_432__37_, r_432__36_, r_432__35_, r_432__34_, r_432__33_, r_432__32_, r_432__31_, r_432__30_, r_432__29_, r_432__28_, r_432__27_, r_432__26_, r_432__25_, r_432__24_, r_432__23_, r_432__22_, r_432__21_, r_432__20_, r_432__19_, r_432__18_, r_432__17_, r_432__16_, r_432__15_, r_432__14_, r_432__13_, r_432__12_, r_432__11_, r_432__10_, r_432__9_, r_432__8_, r_432__7_, r_432__6_, r_432__5_, r_432__4_, r_432__3_, r_432__2_, r_432__1_, r_432__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N863)? data_i : 1'b0;
  assign N862 = sel_i[862];
  assign N863 = N3183;
  assign { r_n_432__63_, r_n_432__62_, r_n_432__61_, r_n_432__60_, r_n_432__59_, r_n_432__58_, r_n_432__57_, r_n_432__56_, r_n_432__55_, r_n_432__54_, r_n_432__53_, r_n_432__52_, r_n_432__51_, r_n_432__50_, r_n_432__49_, r_n_432__48_, r_n_432__47_, r_n_432__46_, r_n_432__45_, r_n_432__44_, r_n_432__43_, r_n_432__42_, r_n_432__41_, r_n_432__40_, r_n_432__39_, r_n_432__38_, r_n_432__37_, r_n_432__36_, r_n_432__35_, r_n_432__34_, r_n_432__33_, r_n_432__32_, r_n_432__31_, r_n_432__30_, r_n_432__29_, r_n_432__28_, r_n_432__27_, r_n_432__26_, r_n_432__25_, r_n_432__24_, r_n_432__23_, r_n_432__22_, r_n_432__21_, r_n_432__20_, r_n_432__19_, r_n_432__18_, r_n_432__17_, r_n_432__16_, r_n_432__15_, r_n_432__14_, r_n_432__13_, r_n_432__12_, r_n_432__11_, r_n_432__10_, r_n_432__9_, r_n_432__8_, r_n_432__7_, r_n_432__6_, r_n_432__5_, r_n_432__4_, r_n_432__3_, r_n_432__2_, r_n_432__1_, r_n_432__0_ } = (N864)? { r_433__63_, r_433__62_, r_433__61_, r_433__60_, r_433__59_, r_433__58_, r_433__57_, r_433__56_, r_433__55_, r_433__54_, r_433__53_, r_433__52_, r_433__51_, r_433__50_, r_433__49_, r_433__48_, r_433__47_, r_433__46_, r_433__45_, r_433__44_, r_433__43_, r_433__42_, r_433__41_, r_433__40_, r_433__39_, r_433__38_, r_433__37_, r_433__36_, r_433__35_, r_433__34_, r_433__33_, r_433__32_, r_433__31_, r_433__30_, r_433__29_, r_433__28_, r_433__27_, r_433__26_, r_433__25_, r_433__24_, r_433__23_, r_433__22_, r_433__21_, r_433__20_, r_433__19_, r_433__18_, r_433__17_, r_433__16_, r_433__15_, r_433__14_, r_433__13_, r_433__12_, r_433__11_, r_433__10_, r_433__9_, r_433__8_, r_433__7_, r_433__6_, r_433__5_, r_433__4_, r_433__3_, r_433__2_, r_433__1_, r_433__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N865)? data_i : 1'b0;
  assign N864 = sel_i[864];
  assign N865 = N3188;
  assign { r_n_433__63_, r_n_433__62_, r_n_433__61_, r_n_433__60_, r_n_433__59_, r_n_433__58_, r_n_433__57_, r_n_433__56_, r_n_433__55_, r_n_433__54_, r_n_433__53_, r_n_433__52_, r_n_433__51_, r_n_433__50_, r_n_433__49_, r_n_433__48_, r_n_433__47_, r_n_433__46_, r_n_433__45_, r_n_433__44_, r_n_433__43_, r_n_433__42_, r_n_433__41_, r_n_433__40_, r_n_433__39_, r_n_433__38_, r_n_433__37_, r_n_433__36_, r_n_433__35_, r_n_433__34_, r_n_433__33_, r_n_433__32_, r_n_433__31_, r_n_433__30_, r_n_433__29_, r_n_433__28_, r_n_433__27_, r_n_433__26_, r_n_433__25_, r_n_433__24_, r_n_433__23_, r_n_433__22_, r_n_433__21_, r_n_433__20_, r_n_433__19_, r_n_433__18_, r_n_433__17_, r_n_433__16_, r_n_433__15_, r_n_433__14_, r_n_433__13_, r_n_433__12_, r_n_433__11_, r_n_433__10_, r_n_433__9_, r_n_433__8_, r_n_433__7_, r_n_433__6_, r_n_433__5_, r_n_433__4_, r_n_433__3_, r_n_433__2_, r_n_433__1_, r_n_433__0_ } = (N866)? { r_434__63_, r_434__62_, r_434__61_, r_434__60_, r_434__59_, r_434__58_, r_434__57_, r_434__56_, r_434__55_, r_434__54_, r_434__53_, r_434__52_, r_434__51_, r_434__50_, r_434__49_, r_434__48_, r_434__47_, r_434__46_, r_434__45_, r_434__44_, r_434__43_, r_434__42_, r_434__41_, r_434__40_, r_434__39_, r_434__38_, r_434__37_, r_434__36_, r_434__35_, r_434__34_, r_434__33_, r_434__32_, r_434__31_, r_434__30_, r_434__29_, r_434__28_, r_434__27_, r_434__26_, r_434__25_, r_434__24_, r_434__23_, r_434__22_, r_434__21_, r_434__20_, r_434__19_, r_434__18_, r_434__17_, r_434__16_, r_434__15_, r_434__14_, r_434__13_, r_434__12_, r_434__11_, r_434__10_, r_434__9_, r_434__8_, r_434__7_, r_434__6_, r_434__5_, r_434__4_, r_434__3_, r_434__2_, r_434__1_, r_434__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N867)? data_i : 1'b0;
  assign N866 = sel_i[866];
  assign N867 = N3193;
  assign { r_n_434__63_, r_n_434__62_, r_n_434__61_, r_n_434__60_, r_n_434__59_, r_n_434__58_, r_n_434__57_, r_n_434__56_, r_n_434__55_, r_n_434__54_, r_n_434__53_, r_n_434__52_, r_n_434__51_, r_n_434__50_, r_n_434__49_, r_n_434__48_, r_n_434__47_, r_n_434__46_, r_n_434__45_, r_n_434__44_, r_n_434__43_, r_n_434__42_, r_n_434__41_, r_n_434__40_, r_n_434__39_, r_n_434__38_, r_n_434__37_, r_n_434__36_, r_n_434__35_, r_n_434__34_, r_n_434__33_, r_n_434__32_, r_n_434__31_, r_n_434__30_, r_n_434__29_, r_n_434__28_, r_n_434__27_, r_n_434__26_, r_n_434__25_, r_n_434__24_, r_n_434__23_, r_n_434__22_, r_n_434__21_, r_n_434__20_, r_n_434__19_, r_n_434__18_, r_n_434__17_, r_n_434__16_, r_n_434__15_, r_n_434__14_, r_n_434__13_, r_n_434__12_, r_n_434__11_, r_n_434__10_, r_n_434__9_, r_n_434__8_, r_n_434__7_, r_n_434__6_, r_n_434__5_, r_n_434__4_, r_n_434__3_, r_n_434__2_, r_n_434__1_, r_n_434__0_ } = (N868)? { r_435__63_, r_435__62_, r_435__61_, r_435__60_, r_435__59_, r_435__58_, r_435__57_, r_435__56_, r_435__55_, r_435__54_, r_435__53_, r_435__52_, r_435__51_, r_435__50_, r_435__49_, r_435__48_, r_435__47_, r_435__46_, r_435__45_, r_435__44_, r_435__43_, r_435__42_, r_435__41_, r_435__40_, r_435__39_, r_435__38_, r_435__37_, r_435__36_, r_435__35_, r_435__34_, r_435__33_, r_435__32_, r_435__31_, r_435__30_, r_435__29_, r_435__28_, r_435__27_, r_435__26_, r_435__25_, r_435__24_, r_435__23_, r_435__22_, r_435__21_, r_435__20_, r_435__19_, r_435__18_, r_435__17_, r_435__16_, r_435__15_, r_435__14_, r_435__13_, r_435__12_, r_435__11_, r_435__10_, r_435__9_, r_435__8_, r_435__7_, r_435__6_, r_435__5_, r_435__4_, r_435__3_, r_435__2_, r_435__1_, r_435__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N869)? data_i : 1'b0;
  assign N868 = sel_i[868];
  assign N869 = N3198;
  assign { r_n_435__63_, r_n_435__62_, r_n_435__61_, r_n_435__60_, r_n_435__59_, r_n_435__58_, r_n_435__57_, r_n_435__56_, r_n_435__55_, r_n_435__54_, r_n_435__53_, r_n_435__52_, r_n_435__51_, r_n_435__50_, r_n_435__49_, r_n_435__48_, r_n_435__47_, r_n_435__46_, r_n_435__45_, r_n_435__44_, r_n_435__43_, r_n_435__42_, r_n_435__41_, r_n_435__40_, r_n_435__39_, r_n_435__38_, r_n_435__37_, r_n_435__36_, r_n_435__35_, r_n_435__34_, r_n_435__33_, r_n_435__32_, r_n_435__31_, r_n_435__30_, r_n_435__29_, r_n_435__28_, r_n_435__27_, r_n_435__26_, r_n_435__25_, r_n_435__24_, r_n_435__23_, r_n_435__22_, r_n_435__21_, r_n_435__20_, r_n_435__19_, r_n_435__18_, r_n_435__17_, r_n_435__16_, r_n_435__15_, r_n_435__14_, r_n_435__13_, r_n_435__12_, r_n_435__11_, r_n_435__10_, r_n_435__9_, r_n_435__8_, r_n_435__7_, r_n_435__6_, r_n_435__5_, r_n_435__4_, r_n_435__3_, r_n_435__2_, r_n_435__1_, r_n_435__0_ } = (N870)? { r_436__63_, r_436__62_, r_436__61_, r_436__60_, r_436__59_, r_436__58_, r_436__57_, r_436__56_, r_436__55_, r_436__54_, r_436__53_, r_436__52_, r_436__51_, r_436__50_, r_436__49_, r_436__48_, r_436__47_, r_436__46_, r_436__45_, r_436__44_, r_436__43_, r_436__42_, r_436__41_, r_436__40_, r_436__39_, r_436__38_, r_436__37_, r_436__36_, r_436__35_, r_436__34_, r_436__33_, r_436__32_, r_436__31_, r_436__30_, r_436__29_, r_436__28_, r_436__27_, r_436__26_, r_436__25_, r_436__24_, r_436__23_, r_436__22_, r_436__21_, r_436__20_, r_436__19_, r_436__18_, r_436__17_, r_436__16_, r_436__15_, r_436__14_, r_436__13_, r_436__12_, r_436__11_, r_436__10_, r_436__9_, r_436__8_, r_436__7_, r_436__6_, r_436__5_, r_436__4_, r_436__3_, r_436__2_, r_436__1_, r_436__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N871)? data_i : 1'b0;
  assign N870 = sel_i[870];
  assign N871 = N3203;
  assign { r_n_436__63_, r_n_436__62_, r_n_436__61_, r_n_436__60_, r_n_436__59_, r_n_436__58_, r_n_436__57_, r_n_436__56_, r_n_436__55_, r_n_436__54_, r_n_436__53_, r_n_436__52_, r_n_436__51_, r_n_436__50_, r_n_436__49_, r_n_436__48_, r_n_436__47_, r_n_436__46_, r_n_436__45_, r_n_436__44_, r_n_436__43_, r_n_436__42_, r_n_436__41_, r_n_436__40_, r_n_436__39_, r_n_436__38_, r_n_436__37_, r_n_436__36_, r_n_436__35_, r_n_436__34_, r_n_436__33_, r_n_436__32_, r_n_436__31_, r_n_436__30_, r_n_436__29_, r_n_436__28_, r_n_436__27_, r_n_436__26_, r_n_436__25_, r_n_436__24_, r_n_436__23_, r_n_436__22_, r_n_436__21_, r_n_436__20_, r_n_436__19_, r_n_436__18_, r_n_436__17_, r_n_436__16_, r_n_436__15_, r_n_436__14_, r_n_436__13_, r_n_436__12_, r_n_436__11_, r_n_436__10_, r_n_436__9_, r_n_436__8_, r_n_436__7_, r_n_436__6_, r_n_436__5_, r_n_436__4_, r_n_436__3_, r_n_436__2_, r_n_436__1_, r_n_436__0_ } = (N872)? { r_437__63_, r_437__62_, r_437__61_, r_437__60_, r_437__59_, r_437__58_, r_437__57_, r_437__56_, r_437__55_, r_437__54_, r_437__53_, r_437__52_, r_437__51_, r_437__50_, r_437__49_, r_437__48_, r_437__47_, r_437__46_, r_437__45_, r_437__44_, r_437__43_, r_437__42_, r_437__41_, r_437__40_, r_437__39_, r_437__38_, r_437__37_, r_437__36_, r_437__35_, r_437__34_, r_437__33_, r_437__32_, r_437__31_, r_437__30_, r_437__29_, r_437__28_, r_437__27_, r_437__26_, r_437__25_, r_437__24_, r_437__23_, r_437__22_, r_437__21_, r_437__20_, r_437__19_, r_437__18_, r_437__17_, r_437__16_, r_437__15_, r_437__14_, r_437__13_, r_437__12_, r_437__11_, r_437__10_, r_437__9_, r_437__8_, r_437__7_, r_437__6_, r_437__5_, r_437__4_, r_437__3_, r_437__2_, r_437__1_, r_437__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N873)? data_i : 1'b0;
  assign N872 = sel_i[872];
  assign N873 = N3208;
  assign { r_n_437__63_, r_n_437__62_, r_n_437__61_, r_n_437__60_, r_n_437__59_, r_n_437__58_, r_n_437__57_, r_n_437__56_, r_n_437__55_, r_n_437__54_, r_n_437__53_, r_n_437__52_, r_n_437__51_, r_n_437__50_, r_n_437__49_, r_n_437__48_, r_n_437__47_, r_n_437__46_, r_n_437__45_, r_n_437__44_, r_n_437__43_, r_n_437__42_, r_n_437__41_, r_n_437__40_, r_n_437__39_, r_n_437__38_, r_n_437__37_, r_n_437__36_, r_n_437__35_, r_n_437__34_, r_n_437__33_, r_n_437__32_, r_n_437__31_, r_n_437__30_, r_n_437__29_, r_n_437__28_, r_n_437__27_, r_n_437__26_, r_n_437__25_, r_n_437__24_, r_n_437__23_, r_n_437__22_, r_n_437__21_, r_n_437__20_, r_n_437__19_, r_n_437__18_, r_n_437__17_, r_n_437__16_, r_n_437__15_, r_n_437__14_, r_n_437__13_, r_n_437__12_, r_n_437__11_, r_n_437__10_, r_n_437__9_, r_n_437__8_, r_n_437__7_, r_n_437__6_, r_n_437__5_, r_n_437__4_, r_n_437__3_, r_n_437__2_, r_n_437__1_, r_n_437__0_ } = (N874)? { r_438__63_, r_438__62_, r_438__61_, r_438__60_, r_438__59_, r_438__58_, r_438__57_, r_438__56_, r_438__55_, r_438__54_, r_438__53_, r_438__52_, r_438__51_, r_438__50_, r_438__49_, r_438__48_, r_438__47_, r_438__46_, r_438__45_, r_438__44_, r_438__43_, r_438__42_, r_438__41_, r_438__40_, r_438__39_, r_438__38_, r_438__37_, r_438__36_, r_438__35_, r_438__34_, r_438__33_, r_438__32_, r_438__31_, r_438__30_, r_438__29_, r_438__28_, r_438__27_, r_438__26_, r_438__25_, r_438__24_, r_438__23_, r_438__22_, r_438__21_, r_438__20_, r_438__19_, r_438__18_, r_438__17_, r_438__16_, r_438__15_, r_438__14_, r_438__13_, r_438__12_, r_438__11_, r_438__10_, r_438__9_, r_438__8_, r_438__7_, r_438__6_, r_438__5_, r_438__4_, r_438__3_, r_438__2_, r_438__1_, r_438__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N875)? data_i : 1'b0;
  assign N874 = sel_i[874];
  assign N875 = N3213;
  assign { r_n_438__63_, r_n_438__62_, r_n_438__61_, r_n_438__60_, r_n_438__59_, r_n_438__58_, r_n_438__57_, r_n_438__56_, r_n_438__55_, r_n_438__54_, r_n_438__53_, r_n_438__52_, r_n_438__51_, r_n_438__50_, r_n_438__49_, r_n_438__48_, r_n_438__47_, r_n_438__46_, r_n_438__45_, r_n_438__44_, r_n_438__43_, r_n_438__42_, r_n_438__41_, r_n_438__40_, r_n_438__39_, r_n_438__38_, r_n_438__37_, r_n_438__36_, r_n_438__35_, r_n_438__34_, r_n_438__33_, r_n_438__32_, r_n_438__31_, r_n_438__30_, r_n_438__29_, r_n_438__28_, r_n_438__27_, r_n_438__26_, r_n_438__25_, r_n_438__24_, r_n_438__23_, r_n_438__22_, r_n_438__21_, r_n_438__20_, r_n_438__19_, r_n_438__18_, r_n_438__17_, r_n_438__16_, r_n_438__15_, r_n_438__14_, r_n_438__13_, r_n_438__12_, r_n_438__11_, r_n_438__10_, r_n_438__9_, r_n_438__8_, r_n_438__7_, r_n_438__6_, r_n_438__5_, r_n_438__4_, r_n_438__3_, r_n_438__2_, r_n_438__1_, r_n_438__0_ } = (N876)? { r_439__63_, r_439__62_, r_439__61_, r_439__60_, r_439__59_, r_439__58_, r_439__57_, r_439__56_, r_439__55_, r_439__54_, r_439__53_, r_439__52_, r_439__51_, r_439__50_, r_439__49_, r_439__48_, r_439__47_, r_439__46_, r_439__45_, r_439__44_, r_439__43_, r_439__42_, r_439__41_, r_439__40_, r_439__39_, r_439__38_, r_439__37_, r_439__36_, r_439__35_, r_439__34_, r_439__33_, r_439__32_, r_439__31_, r_439__30_, r_439__29_, r_439__28_, r_439__27_, r_439__26_, r_439__25_, r_439__24_, r_439__23_, r_439__22_, r_439__21_, r_439__20_, r_439__19_, r_439__18_, r_439__17_, r_439__16_, r_439__15_, r_439__14_, r_439__13_, r_439__12_, r_439__11_, r_439__10_, r_439__9_, r_439__8_, r_439__7_, r_439__6_, r_439__5_, r_439__4_, r_439__3_, r_439__2_, r_439__1_, r_439__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N877)? data_i : 1'b0;
  assign N876 = sel_i[876];
  assign N877 = N3218;
  assign { r_n_439__63_, r_n_439__62_, r_n_439__61_, r_n_439__60_, r_n_439__59_, r_n_439__58_, r_n_439__57_, r_n_439__56_, r_n_439__55_, r_n_439__54_, r_n_439__53_, r_n_439__52_, r_n_439__51_, r_n_439__50_, r_n_439__49_, r_n_439__48_, r_n_439__47_, r_n_439__46_, r_n_439__45_, r_n_439__44_, r_n_439__43_, r_n_439__42_, r_n_439__41_, r_n_439__40_, r_n_439__39_, r_n_439__38_, r_n_439__37_, r_n_439__36_, r_n_439__35_, r_n_439__34_, r_n_439__33_, r_n_439__32_, r_n_439__31_, r_n_439__30_, r_n_439__29_, r_n_439__28_, r_n_439__27_, r_n_439__26_, r_n_439__25_, r_n_439__24_, r_n_439__23_, r_n_439__22_, r_n_439__21_, r_n_439__20_, r_n_439__19_, r_n_439__18_, r_n_439__17_, r_n_439__16_, r_n_439__15_, r_n_439__14_, r_n_439__13_, r_n_439__12_, r_n_439__11_, r_n_439__10_, r_n_439__9_, r_n_439__8_, r_n_439__7_, r_n_439__6_, r_n_439__5_, r_n_439__4_, r_n_439__3_, r_n_439__2_, r_n_439__1_, r_n_439__0_ } = (N878)? { r_440__63_, r_440__62_, r_440__61_, r_440__60_, r_440__59_, r_440__58_, r_440__57_, r_440__56_, r_440__55_, r_440__54_, r_440__53_, r_440__52_, r_440__51_, r_440__50_, r_440__49_, r_440__48_, r_440__47_, r_440__46_, r_440__45_, r_440__44_, r_440__43_, r_440__42_, r_440__41_, r_440__40_, r_440__39_, r_440__38_, r_440__37_, r_440__36_, r_440__35_, r_440__34_, r_440__33_, r_440__32_, r_440__31_, r_440__30_, r_440__29_, r_440__28_, r_440__27_, r_440__26_, r_440__25_, r_440__24_, r_440__23_, r_440__22_, r_440__21_, r_440__20_, r_440__19_, r_440__18_, r_440__17_, r_440__16_, r_440__15_, r_440__14_, r_440__13_, r_440__12_, r_440__11_, r_440__10_, r_440__9_, r_440__8_, r_440__7_, r_440__6_, r_440__5_, r_440__4_, r_440__3_, r_440__2_, r_440__1_, r_440__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N879)? data_i : 1'b0;
  assign N878 = sel_i[878];
  assign N879 = N3223;
  assign { r_n_440__63_, r_n_440__62_, r_n_440__61_, r_n_440__60_, r_n_440__59_, r_n_440__58_, r_n_440__57_, r_n_440__56_, r_n_440__55_, r_n_440__54_, r_n_440__53_, r_n_440__52_, r_n_440__51_, r_n_440__50_, r_n_440__49_, r_n_440__48_, r_n_440__47_, r_n_440__46_, r_n_440__45_, r_n_440__44_, r_n_440__43_, r_n_440__42_, r_n_440__41_, r_n_440__40_, r_n_440__39_, r_n_440__38_, r_n_440__37_, r_n_440__36_, r_n_440__35_, r_n_440__34_, r_n_440__33_, r_n_440__32_, r_n_440__31_, r_n_440__30_, r_n_440__29_, r_n_440__28_, r_n_440__27_, r_n_440__26_, r_n_440__25_, r_n_440__24_, r_n_440__23_, r_n_440__22_, r_n_440__21_, r_n_440__20_, r_n_440__19_, r_n_440__18_, r_n_440__17_, r_n_440__16_, r_n_440__15_, r_n_440__14_, r_n_440__13_, r_n_440__12_, r_n_440__11_, r_n_440__10_, r_n_440__9_, r_n_440__8_, r_n_440__7_, r_n_440__6_, r_n_440__5_, r_n_440__4_, r_n_440__3_, r_n_440__2_, r_n_440__1_, r_n_440__0_ } = (N880)? { r_441__63_, r_441__62_, r_441__61_, r_441__60_, r_441__59_, r_441__58_, r_441__57_, r_441__56_, r_441__55_, r_441__54_, r_441__53_, r_441__52_, r_441__51_, r_441__50_, r_441__49_, r_441__48_, r_441__47_, r_441__46_, r_441__45_, r_441__44_, r_441__43_, r_441__42_, r_441__41_, r_441__40_, r_441__39_, r_441__38_, r_441__37_, r_441__36_, r_441__35_, r_441__34_, r_441__33_, r_441__32_, r_441__31_, r_441__30_, r_441__29_, r_441__28_, r_441__27_, r_441__26_, r_441__25_, r_441__24_, r_441__23_, r_441__22_, r_441__21_, r_441__20_, r_441__19_, r_441__18_, r_441__17_, r_441__16_, r_441__15_, r_441__14_, r_441__13_, r_441__12_, r_441__11_, r_441__10_, r_441__9_, r_441__8_, r_441__7_, r_441__6_, r_441__5_, r_441__4_, r_441__3_, r_441__2_, r_441__1_, r_441__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N881)? data_i : 1'b0;
  assign N880 = sel_i[880];
  assign N881 = N3228;
  assign { r_n_441__63_, r_n_441__62_, r_n_441__61_, r_n_441__60_, r_n_441__59_, r_n_441__58_, r_n_441__57_, r_n_441__56_, r_n_441__55_, r_n_441__54_, r_n_441__53_, r_n_441__52_, r_n_441__51_, r_n_441__50_, r_n_441__49_, r_n_441__48_, r_n_441__47_, r_n_441__46_, r_n_441__45_, r_n_441__44_, r_n_441__43_, r_n_441__42_, r_n_441__41_, r_n_441__40_, r_n_441__39_, r_n_441__38_, r_n_441__37_, r_n_441__36_, r_n_441__35_, r_n_441__34_, r_n_441__33_, r_n_441__32_, r_n_441__31_, r_n_441__30_, r_n_441__29_, r_n_441__28_, r_n_441__27_, r_n_441__26_, r_n_441__25_, r_n_441__24_, r_n_441__23_, r_n_441__22_, r_n_441__21_, r_n_441__20_, r_n_441__19_, r_n_441__18_, r_n_441__17_, r_n_441__16_, r_n_441__15_, r_n_441__14_, r_n_441__13_, r_n_441__12_, r_n_441__11_, r_n_441__10_, r_n_441__9_, r_n_441__8_, r_n_441__7_, r_n_441__6_, r_n_441__5_, r_n_441__4_, r_n_441__3_, r_n_441__2_, r_n_441__1_, r_n_441__0_ } = (N882)? { r_442__63_, r_442__62_, r_442__61_, r_442__60_, r_442__59_, r_442__58_, r_442__57_, r_442__56_, r_442__55_, r_442__54_, r_442__53_, r_442__52_, r_442__51_, r_442__50_, r_442__49_, r_442__48_, r_442__47_, r_442__46_, r_442__45_, r_442__44_, r_442__43_, r_442__42_, r_442__41_, r_442__40_, r_442__39_, r_442__38_, r_442__37_, r_442__36_, r_442__35_, r_442__34_, r_442__33_, r_442__32_, r_442__31_, r_442__30_, r_442__29_, r_442__28_, r_442__27_, r_442__26_, r_442__25_, r_442__24_, r_442__23_, r_442__22_, r_442__21_, r_442__20_, r_442__19_, r_442__18_, r_442__17_, r_442__16_, r_442__15_, r_442__14_, r_442__13_, r_442__12_, r_442__11_, r_442__10_, r_442__9_, r_442__8_, r_442__7_, r_442__6_, r_442__5_, r_442__4_, r_442__3_, r_442__2_, r_442__1_, r_442__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N883)? data_i : 1'b0;
  assign N882 = sel_i[882];
  assign N883 = N3233;
  assign { r_n_442__63_, r_n_442__62_, r_n_442__61_, r_n_442__60_, r_n_442__59_, r_n_442__58_, r_n_442__57_, r_n_442__56_, r_n_442__55_, r_n_442__54_, r_n_442__53_, r_n_442__52_, r_n_442__51_, r_n_442__50_, r_n_442__49_, r_n_442__48_, r_n_442__47_, r_n_442__46_, r_n_442__45_, r_n_442__44_, r_n_442__43_, r_n_442__42_, r_n_442__41_, r_n_442__40_, r_n_442__39_, r_n_442__38_, r_n_442__37_, r_n_442__36_, r_n_442__35_, r_n_442__34_, r_n_442__33_, r_n_442__32_, r_n_442__31_, r_n_442__30_, r_n_442__29_, r_n_442__28_, r_n_442__27_, r_n_442__26_, r_n_442__25_, r_n_442__24_, r_n_442__23_, r_n_442__22_, r_n_442__21_, r_n_442__20_, r_n_442__19_, r_n_442__18_, r_n_442__17_, r_n_442__16_, r_n_442__15_, r_n_442__14_, r_n_442__13_, r_n_442__12_, r_n_442__11_, r_n_442__10_, r_n_442__9_, r_n_442__8_, r_n_442__7_, r_n_442__6_, r_n_442__5_, r_n_442__4_, r_n_442__3_, r_n_442__2_, r_n_442__1_, r_n_442__0_ } = (N884)? { r_443__63_, r_443__62_, r_443__61_, r_443__60_, r_443__59_, r_443__58_, r_443__57_, r_443__56_, r_443__55_, r_443__54_, r_443__53_, r_443__52_, r_443__51_, r_443__50_, r_443__49_, r_443__48_, r_443__47_, r_443__46_, r_443__45_, r_443__44_, r_443__43_, r_443__42_, r_443__41_, r_443__40_, r_443__39_, r_443__38_, r_443__37_, r_443__36_, r_443__35_, r_443__34_, r_443__33_, r_443__32_, r_443__31_, r_443__30_, r_443__29_, r_443__28_, r_443__27_, r_443__26_, r_443__25_, r_443__24_, r_443__23_, r_443__22_, r_443__21_, r_443__20_, r_443__19_, r_443__18_, r_443__17_, r_443__16_, r_443__15_, r_443__14_, r_443__13_, r_443__12_, r_443__11_, r_443__10_, r_443__9_, r_443__8_, r_443__7_, r_443__6_, r_443__5_, r_443__4_, r_443__3_, r_443__2_, r_443__1_, r_443__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N885)? data_i : 1'b0;
  assign N884 = sel_i[884];
  assign N885 = N3238;
  assign { r_n_443__63_, r_n_443__62_, r_n_443__61_, r_n_443__60_, r_n_443__59_, r_n_443__58_, r_n_443__57_, r_n_443__56_, r_n_443__55_, r_n_443__54_, r_n_443__53_, r_n_443__52_, r_n_443__51_, r_n_443__50_, r_n_443__49_, r_n_443__48_, r_n_443__47_, r_n_443__46_, r_n_443__45_, r_n_443__44_, r_n_443__43_, r_n_443__42_, r_n_443__41_, r_n_443__40_, r_n_443__39_, r_n_443__38_, r_n_443__37_, r_n_443__36_, r_n_443__35_, r_n_443__34_, r_n_443__33_, r_n_443__32_, r_n_443__31_, r_n_443__30_, r_n_443__29_, r_n_443__28_, r_n_443__27_, r_n_443__26_, r_n_443__25_, r_n_443__24_, r_n_443__23_, r_n_443__22_, r_n_443__21_, r_n_443__20_, r_n_443__19_, r_n_443__18_, r_n_443__17_, r_n_443__16_, r_n_443__15_, r_n_443__14_, r_n_443__13_, r_n_443__12_, r_n_443__11_, r_n_443__10_, r_n_443__9_, r_n_443__8_, r_n_443__7_, r_n_443__6_, r_n_443__5_, r_n_443__4_, r_n_443__3_, r_n_443__2_, r_n_443__1_, r_n_443__0_ } = (N886)? { r_444__63_, r_444__62_, r_444__61_, r_444__60_, r_444__59_, r_444__58_, r_444__57_, r_444__56_, r_444__55_, r_444__54_, r_444__53_, r_444__52_, r_444__51_, r_444__50_, r_444__49_, r_444__48_, r_444__47_, r_444__46_, r_444__45_, r_444__44_, r_444__43_, r_444__42_, r_444__41_, r_444__40_, r_444__39_, r_444__38_, r_444__37_, r_444__36_, r_444__35_, r_444__34_, r_444__33_, r_444__32_, r_444__31_, r_444__30_, r_444__29_, r_444__28_, r_444__27_, r_444__26_, r_444__25_, r_444__24_, r_444__23_, r_444__22_, r_444__21_, r_444__20_, r_444__19_, r_444__18_, r_444__17_, r_444__16_, r_444__15_, r_444__14_, r_444__13_, r_444__12_, r_444__11_, r_444__10_, r_444__9_, r_444__8_, r_444__7_, r_444__6_, r_444__5_, r_444__4_, r_444__3_, r_444__2_, r_444__1_, r_444__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N887)? data_i : 1'b0;
  assign N886 = sel_i[886];
  assign N887 = N3243;
  assign { r_n_444__63_, r_n_444__62_, r_n_444__61_, r_n_444__60_, r_n_444__59_, r_n_444__58_, r_n_444__57_, r_n_444__56_, r_n_444__55_, r_n_444__54_, r_n_444__53_, r_n_444__52_, r_n_444__51_, r_n_444__50_, r_n_444__49_, r_n_444__48_, r_n_444__47_, r_n_444__46_, r_n_444__45_, r_n_444__44_, r_n_444__43_, r_n_444__42_, r_n_444__41_, r_n_444__40_, r_n_444__39_, r_n_444__38_, r_n_444__37_, r_n_444__36_, r_n_444__35_, r_n_444__34_, r_n_444__33_, r_n_444__32_, r_n_444__31_, r_n_444__30_, r_n_444__29_, r_n_444__28_, r_n_444__27_, r_n_444__26_, r_n_444__25_, r_n_444__24_, r_n_444__23_, r_n_444__22_, r_n_444__21_, r_n_444__20_, r_n_444__19_, r_n_444__18_, r_n_444__17_, r_n_444__16_, r_n_444__15_, r_n_444__14_, r_n_444__13_, r_n_444__12_, r_n_444__11_, r_n_444__10_, r_n_444__9_, r_n_444__8_, r_n_444__7_, r_n_444__6_, r_n_444__5_, r_n_444__4_, r_n_444__3_, r_n_444__2_, r_n_444__1_, r_n_444__0_ } = (N888)? { r_445__63_, r_445__62_, r_445__61_, r_445__60_, r_445__59_, r_445__58_, r_445__57_, r_445__56_, r_445__55_, r_445__54_, r_445__53_, r_445__52_, r_445__51_, r_445__50_, r_445__49_, r_445__48_, r_445__47_, r_445__46_, r_445__45_, r_445__44_, r_445__43_, r_445__42_, r_445__41_, r_445__40_, r_445__39_, r_445__38_, r_445__37_, r_445__36_, r_445__35_, r_445__34_, r_445__33_, r_445__32_, r_445__31_, r_445__30_, r_445__29_, r_445__28_, r_445__27_, r_445__26_, r_445__25_, r_445__24_, r_445__23_, r_445__22_, r_445__21_, r_445__20_, r_445__19_, r_445__18_, r_445__17_, r_445__16_, r_445__15_, r_445__14_, r_445__13_, r_445__12_, r_445__11_, r_445__10_, r_445__9_, r_445__8_, r_445__7_, r_445__6_, r_445__5_, r_445__4_, r_445__3_, r_445__2_, r_445__1_, r_445__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N889)? data_i : 1'b0;
  assign N888 = sel_i[888];
  assign N889 = N3248;
  assign { r_n_445__63_, r_n_445__62_, r_n_445__61_, r_n_445__60_, r_n_445__59_, r_n_445__58_, r_n_445__57_, r_n_445__56_, r_n_445__55_, r_n_445__54_, r_n_445__53_, r_n_445__52_, r_n_445__51_, r_n_445__50_, r_n_445__49_, r_n_445__48_, r_n_445__47_, r_n_445__46_, r_n_445__45_, r_n_445__44_, r_n_445__43_, r_n_445__42_, r_n_445__41_, r_n_445__40_, r_n_445__39_, r_n_445__38_, r_n_445__37_, r_n_445__36_, r_n_445__35_, r_n_445__34_, r_n_445__33_, r_n_445__32_, r_n_445__31_, r_n_445__30_, r_n_445__29_, r_n_445__28_, r_n_445__27_, r_n_445__26_, r_n_445__25_, r_n_445__24_, r_n_445__23_, r_n_445__22_, r_n_445__21_, r_n_445__20_, r_n_445__19_, r_n_445__18_, r_n_445__17_, r_n_445__16_, r_n_445__15_, r_n_445__14_, r_n_445__13_, r_n_445__12_, r_n_445__11_, r_n_445__10_, r_n_445__9_, r_n_445__8_, r_n_445__7_, r_n_445__6_, r_n_445__5_, r_n_445__4_, r_n_445__3_, r_n_445__2_, r_n_445__1_, r_n_445__0_ } = (N890)? { r_446__63_, r_446__62_, r_446__61_, r_446__60_, r_446__59_, r_446__58_, r_446__57_, r_446__56_, r_446__55_, r_446__54_, r_446__53_, r_446__52_, r_446__51_, r_446__50_, r_446__49_, r_446__48_, r_446__47_, r_446__46_, r_446__45_, r_446__44_, r_446__43_, r_446__42_, r_446__41_, r_446__40_, r_446__39_, r_446__38_, r_446__37_, r_446__36_, r_446__35_, r_446__34_, r_446__33_, r_446__32_, r_446__31_, r_446__30_, r_446__29_, r_446__28_, r_446__27_, r_446__26_, r_446__25_, r_446__24_, r_446__23_, r_446__22_, r_446__21_, r_446__20_, r_446__19_, r_446__18_, r_446__17_, r_446__16_, r_446__15_, r_446__14_, r_446__13_, r_446__12_, r_446__11_, r_446__10_, r_446__9_, r_446__8_, r_446__7_, r_446__6_, r_446__5_, r_446__4_, r_446__3_, r_446__2_, r_446__1_, r_446__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N891)? data_i : 1'b0;
  assign N890 = sel_i[890];
  assign N891 = N3253;
  assign { r_n_446__63_, r_n_446__62_, r_n_446__61_, r_n_446__60_, r_n_446__59_, r_n_446__58_, r_n_446__57_, r_n_446__56_, r_n_446__55_, r_n_446__54_, r_n_446__53_, r_n_446__52_, r_n_446__51_, r_n_446__50_, r_n_446__49_, r_n_446__48_, r_n_446__47_, r_n_446__46_, r_n_446__45_, r_n_446__44_, r_n_446__43_, r_n_446__42_, r_n_446__41_, r_n_446__40_, r_n_446__39_, r_n_446__38_, r_n_446__37_, r_n_446__36_, r_n_446__35_, r_n_446__34_, r_n_446__33_, r_n_446__32_, r_n_446__31_, r_n_446__30_, r_n_446__29_, r_n_446__28_, r_n_446__27_, r_n_446__26_, r_n_446__25_, r_n_446__24_, r_n_446__23_, r_n_446__22_, r_n_446__21_, r_n_446__20_, r_n_446__19_, r_n_446__18_, r_n_446__17_, r_n_446__16_, r_n_446__15_, r_n_446__14_, r_n_446__13_, r_n_446__12_, r_n_446__11_, r_n_446__10_, r_n_446__9_, r_n_446__8_, r_n_446__7_, r_n_446__6_, r_n_446__5_, r_n_446__4_, r_n_446__3_, r_n_446__2_, r_n_446__1_, r_n_446__0_ } = (N892)? { r_447__63_, r_447__62_, r_447__61_, r_447__60_, r_447__59_, r_447__58_, r_447__57_, r_447__56_, r_447__55_, r_447__54_, r_447__53_, r_447__52_, r_447__51_, r_447__50_, r_447__49_, r_447__48_, r_447__47_, r_447__46_, r_447__45_, r_447__44_, r_447__43_, r_447__42_, r_447__41_, r_447__40_, r_447__39_, r_447__38_, r_447__37_, r_447__36_, r_447__35_, r_447__34_, r_447__33_, r_447__32_, r_447__31_, r_447__30_, r_447__29_, r_447__28_, r_447__27_, r_447__26_, r_447__25_, r_447__24_, r_447__23_, r_447__22_, r_447__21_, r_447__20_, r_447__19_, r_447__18_, r_447__17_, r_447__16_, r_447__15_, r_447__14_, r_447__13_, r_447__12_, r_447__11_, r_447__10_, r_447__9_, r_447__8_, r_447__7_, r_447__6_, r_447__5_, r_447__4_, r_447__3_, r_447__2_, r_447__1_, r_447__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N893)? data_i : 1'b0;
  assign N892 = sel_i[892];
  assign N893 = N3258;
  assign { r_n_447__63_, r_n_447__62_, r_n_447__61_, r_n_447__60_, r_n_447__59_, r_n_447__58_, r_n_447__57_, r_n_447__56_, r_n_447__55_, r_n_447__54_, r_n_447__53_, r_n_447__52_, r_n_447__51_, r_n_447__50_, r_n_447__49_, r_n_447__48_, r_n_447__47_, r_n_447__46_, r_n_447__45_, r_n_447__44_, r_n_447__43_, r_n_447__42_, r_n_447__41_, r_n_447__40_, r_n_447__39_, r_n_447__38_, r_n_447__37_, r_n_447__36_, r_n_447__35_, r_n_447__34_, r_n_447__33_, r_n_447__32_, r_n_447__31_, r_n_447__30_, r_n_447__29_, r_n_447__28_, r_n_447__27_, r_n_447__26_, r_n_447__25_, r_n_447__24_, r_n_447__23_, r_n_447__22_, r_n_447__21_, r_n_447__20_, r_n_447__19_, r_n_447__18_, r_n_447__17_, r_n_447__16_, r_n_447__15_, r_n_447__14_, r_n_447__13_, r_n_447__12_, r_n_447__11_, r_n_447__10_, r_n_447__9_, r_n_447__8_, r_n_447__7_, r_n_447__6_, r_n_447__5_, r_n_447__4_, r_n_447__3_, r_n_447__2_, r_n_447__1_, r_n_447__0_ } = (N894)? { r_448__63_, r_448__62_, r_448__61_, r_448__60_, r_448__59_, r_448__58_, r_448__57_, r_448__56_, r_448__55_, r_448__54_, r_448__53_, r_448__52_, r_448__51_, r_448__50_, r_448__49_, r_448__48_, r_448__47_, r_448__46_, r_448__45_, r_448__44_, r_448__43_, r_448__42_, r_448__41_, r_448__40_, r_448__39_, r_448__38_, r_448__37_, r_448__36_, r_448__35_, r_448__34_, r_448__33_, r_448__32_, r_448__31_, r_448__30_, r_448__29_, r_448__28_, r_448__27_, r_448__26_, r_448__25_, r_448__24_, r_448__23_, r_448__22_, r_448__21_, r_448__20_, r_448__19_, r_448__18_, r_448__17_, r_448__16_, r_448__15_, r_448__14_, r_448__13_, r_448__12_, r_448__11_, r_448__10_, r_448__9_, r_448__8_, r_448__7_, r_448__6_, r_448__5_, r_448__4_, r_448__3_, r_448__2_, r_448__1_, r_448__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N895)? data_i : 1'b0;
  assign N894 = sel_i[894];
  assign N895 = N3263;
  assign { r_n_448__63_, r_n_448__62_, r_n_448__61_, r_n_448__60_, r_n_448__59_, r_n_448__58_, r_n_448__57_, r_n_448__56_, r_n_448__55_, r_n_448__54_, r_n_448__53_, r_n_448__52_, r_n_448__51_, r_n_448__50_, r_n_448__49_, r_n_448__48_, r_n_448__47_, r_n_448__46_, r_n_448__45_, r_n_448__44_, r_n_448__43_, r_n_448__42_, r_n_448__41_, r_n_448__40_, r_n_448__39_, r_n_448__38_, r_n_448__37_, r_n_448__36_, r_n_448__35_, r_n_448__34_, r_n_448__33_, r_n_448__32_, r_n_448__31_, r_n_448__30_, r_n_448__29_, r_n_448__28_, r_n_448__27_, r_n_448__26_, r_n_448__25_, r_n_448__24_, r_n_448__23_, r_n_448__22_, r_n_448__21_, r_n_448__20_, r_n_448__19_, r_n_448__18_, r_n_448__17_, r_n_448__16_, r_n_448__15_, r_n_448__14_, r_n_448__13_, r_n_448__12_, r_n_448__11_, r_n_448__10_, r_n_448__9_, r_n_448__8_, r_n_448__7_, r_n_448__6_, r_n_448__5_, r_n_448__4_, r_n_448__3_, r_n_448__2_, r_n_448__1_, r_n_448__0_ } = (N896)? { r_449__63_, r_449__62_, r_449__61_, r_449__60_, r_449__59_, r_449__58_, r_449__57_, r_449__56_, r_449__55_, r_449__54_, r_449__53_, r_449__52_, r_449__51_, r_449__50_, r_449__49_, r_449__48_, r_449__47_, r_449__46_, r_449__45_, r_449__44_, r_449__43_, r_449__42_, r_449__41_, r_449__40_, r_449__39_, r_449__38_, r_449__37_, r_449__36_, r_449__35_, r_449__34_, r_449__33_, r_449__32_, r_449__31_, r_449__30_, r_449__29_, r_449__28_, r_449__27_, r_449__26_, r_449__25_, r_449__24_, r_449__23_, r_449__22_, r_449__21_, r_449__20_, r_449__19_, r_449__18_, r_449__17_, r_449__16_, r_449__15_, r_449__14_, r_449__13_, r_449__12_, r_449__11_, r_449__10_, r_449__9_, r_449__8_, r_449__7_, r_449__6_, r_449__5_, r_449__4_, r_449__3_, r_449__2_, r_449__1_, r_449__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N897)? data_i : 1'b0;
  assign N896 = sel_i[896];
  assign N897 = N3268;
  assign { r_n_449__63_, r_n_449__62_, r_n_449__61_, r_n_449__60_, r_n_449__59_, r_n_449__58_, r_n_449__57_, r_n_449__56_, r_n_449__55_, r_n_449__54_, r_n_449__53_, r_n_449__52_, r_n_449__51_, r_n_449__50_, r_n_449__49_, r_n_449__48_, r_n_449__47_, r_n_449__46_, r_n_449__45_, r_n_449__44_, r_n_449__43_, r_n_449__42_, r_n_449__41_, r_n_449__40_, r_n_449__39_, r_n_449__38_, r_n_449__37_, r_n_449__36_, r_n_449__35_, r_n_449__34_, r_n_449__33_, r_n_449__32_, r_n_449__31_, r_n_449__30_, r_n_449__29_, r_n_449__28_, r_n_449__27_, r_n_449__26_, r_n_449__25_, r_n_449__24_, r_n_449__23_, r_n_449__22_, r_n_449__21_, r_n_449__20_, r_n_449__19_, r_n_449__18_, r_n_449__17_, r_n_449__16_, r_n_449__15_, r_n_449__14_, r_n_449__13_, r_n_449__12_, r_n_449__11_, r_n_449__10_, r_n_449__9_, r_n_449__8_, r_n_449__7_, r_n_449__6_, r_n_449__5_, r_n_449__4_, r_n_449__3_, r_n_449__2_, r_n_449__1_, r_n_449__0_ } = (N898)? { r_450__63_, r_450__62_, r_450__61_, r_450__60_, r_450__59_, r_450__58_, r_450__57_, r_450__56_, r_450__55_, r_450__54_, r_450__53_, r_450__52_, r_450__51_, r_450__50_, r_450__49_, r_450__48_, r_450__47_, r_450__46_, r_450__45_, r_450__44_, r_450__43_, r_450__42_, r_450__41_, r_450__40_, r_450__39_, r_450__38_, r_450__37_, r_450__36_, r_450__35_, r_450__34_, r_450__33_, r_450__32_, r_450__31_, r_450__30_, r_450__29_, r_450__28_, r_450__27_, r_450__26_, r_450__25_, r_450__24_, r_450__23_, r_450__22_, r_450__21_, r_450__20_, r_450__19_, r_450__18_, r_450__17_, r_450__16_, r_450__15_, r_450__14_, r_450__13_, r_450__12_, r_450__11_, r_450__10_, r_450__9_, r_450__8_, r_450__7_, r_450__6_, r_450__5_, r_450__4_, r_450__3_, r_450__2_, r_450__1_, r_450__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N899)? data_i : 1'b0;
  assign N898 = sel_i[898];
  assign N899 = N3273;
  assign { r_n_450__63_, r_n_450__62_, r_n_450__61_, r_n_450__60_, r_n_450__59_, r_n_450__58_, r_n_450__57_, r_n_450__56_, r_n_450__55_, r_n_450__54_, r_n_450__53_, r_n_450__52_, r_n_450__51_, r_n_450__50_, r_n_450__49_, r_n_450__48_, r_n_450__47_, r_n_450__46_, r_n_450__45_, r_n_450__44_, r_n_450__43_, r_n_450__42_, r_n_450__41_, r_n_450__40_, r_n_450__39_, r_n_450__38_, r_n_450__37_, r_n_450__36_, r_n_450__35_, r_n_450__34_, r_n_450__33_, r_n_450__32_, r_n_450__31_, r_n_450__30_, r_n_450__29_, r_n_450__28_, r_n_450__27_, r_n_450__26_, r_n_450__25_, r_n_450__24_, r_n_450__23_, r_n_450__22_, r_n_450__21_, r_n_450__20_, r_n_450__19_, r_n_450__18_, r_n_450__17_, r_n_450__16_, r_n_450__15_, r_n_450__14_, r_n_450__13_, r_n_450__12_, r_n_450__11_, r_n_450__10_, r_n_450__9_, r_n_450__8_, r_n_450__7_, r_n_450__6_, r_n_450__5_, r_n_450__4_, r_n_450__3_, r_n_450__2_, r_n_450__1_, r_n_450__0_ } = (N900)? { r_451__63_, r_451__62_, r_451__61_, r_451__60_, r_451__59_, r_451__58_, r_451__57_, r_451__56_, r_451__55_, r_451__54_, r_451__53_, r_451__52_, r_451__51_, r_451__50_, r_451__49_, r_451__48_, r_451__47_, r_451__46_, r_451__45_, r_451__44_, r_451__43_, r_451__42_, r_451__41_, r_451__40_, r_451__39_, r_451__38_, r_451__37_, r_451__36_, r_451__35_, r_451__34_, r_451__33_, r_451__32_, r_451__31_, r_451__30_, r_451__29_, r_451__28_, r_451__27_, r_451__26_, r_451__25_, r_451__24_, r_451__23_, r_451__22_, r_451__21_, r_451__20_, r_451__19_, r_451__18_, r_451__17_, r_451__16_, r_451__15_, r_451__14_, r_451__13_, r_451__12_, r_451__11_, r_451__10_, r_451__9_, r_451__8_, r_451__7_, r_451__6_, r_451__5_, r_451__4_, r_451__3_, r_451__2_, r_451__1_, r_451__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N901)? data_i : 1'b0;
  assign N900 = sel_i[900];
  assign N901 = N3278;
  assign { r_n_451__63_, r_n_451__62_, r_n_451__61_, r_n_451__60_, r_n_451__59_, r_n_451__58_, r_n_451__57_, r_n_451__56_, r_n_451__55_, r_n_451__54_, r_n_451__53_, r_n_451__52_, r_n_451__51_, r_n_451__50_, r_n_451__49_, r_n_451__48_, r_n_451__47_, r_n_451__46_, r_n_451__45_, r_n_451__44_, r_n_451__43_, r_n_451__42_, r_n_451__41_, r_n_451__40_, r_n_451__39_, r_n_451__38_, r_n_451__37_, r_n_451__36_, r_n_451__35_, r_n_451__34_, r_n_451__33_, r_n_451__32_, r_n_451__31_, r_n_451__30_, r_n_451__29_, r_n_451__28_, r_n_451__27_, r_n_451__26_, r_n_451__25_, r_n_451__24_, r_n_451__23_, r_n_451__22_, r_n_451__21_, r_n_451__20_, r_n_451__19_, r_n_451__18_, r_n_451__17_, r_n_451__16_, r_n_451__15_, r_n_451__14_, r_n_451__13_, r_n_451__12_, r_n_451__11_, r_n_451__10_, r_n_451__9_, r_n_451__8_, r_n_451__7_, r_n_451__6_, r_n_451__5_, r_n_451__4_, r_n_451__3_, r_n_451__2_, r_n_451__1_, r_n_451__0_ } = (N902)? { r_452__63_, r_452__62_, r_452__61_, r_452__60_, r_452__59_, r_452__58_, r_452__57_, r_452__56_, r_452__55_, r_452__54_, r_452__53_, r_452__52_, r_452__51_, r_452__50_, r_452__49_, r_452__48_, r_452__47_, r_452__46_, r_452__45_, r_452__44_, r_452__43_, r_452__42_, r_452__41_, r_452__40_, r_452__39_, r_452__38_, r_452__37_, r_452__36_, r_452__35_, r_452__34_, r_452__33_, r_452__32_, r_452__31_, r_452__30_, r_452__29_, r_452__28_, r_452__27_, r_452__26_, r_452__25_, r_452__24_, r_452__23_, r_452__22_, r_452__21_, r_452__20_, r_452__19_, r_452__18_, r_452__17_, r_452__16_, r_452__15_, r_452__14_, r_452__13_, r_452__12_, r_452__11_, r_452__10_, r_452__9_, r_452__8_, r_452__7_, r_452__6_, r_452__5_, r_452__4_, r_452__3_, r_452__2_, r_452__1_, r_452__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N903)? data_i : 1'b0;
  assign N902 = sel_i[902];
  assign N903 = N3283;
  assign { r_n_452__63_, r_n_452__62_, r_n_452__61_, r_n_452__60_, r_n_452__59_, r_n_452__58_, r_n_452__57_, r_n_452__56_, r_n_452__55_, r_n_452__54_, r_n_452__53_, r_n_452__52_, r_n_452__51_, r_n_452__50_, r_n_452__49_, r_n_452__48_, r_n_452__47_, r_n_452__46_, r_n_452__45_, r_n_452__44_, r_n_452__43_, r_n_452__42_, r_n_452__41_, r_n_452__40_, r_n_452__39_, r_n_452__38_, r_n_452__37_, r_n_452__36_, r_n_452__35_, r_n_452__34_, r_n_452__33_, r_n_452__32_, r_n_452__31_, r_n_452__30_, r_n_452__29_, r_n_452__28_, r_n_452__27_, r_n_452__26_, r_n_452__25_, r_n_452__24_, r_n_452__23_, r_n_452__22_, r_n_452__21_, r_n_452__20_, r_n_452__19_, r_n_452__18_, r_n_452__17_, r_n_452__16_, r_n_452__15_, r_n_452__14_, r_n_452__13_, r_n_452__12_, r_n_452__11_, r_n_452__10_, r_n_452__9_, r_n_452__8_, r_n_452__7_, r_n_452__6_, r_n_452__5_, r_n_452__4_, r_n_452__3_, r_n_452__2_, r_n_452__1_, r_n_452__0_ } = (N904)? { r_453__63_, r_453__62_, r_453__61_, r_453__60_, r_453__59_, r_453__58_, r_453__57_, r_453__56_, r_453__55_, r_453__54_, r_453__53_, r_453__52_, r_453__51_, r_453__50_, r_453__49_, r_453__48_, r_453__47_, r_453__46_, r_453__45_, r_453__44_, r_453__43_, r_453__42_, r_453__41_, r_453__40_, r_453__39_, r_453__38_, r_453__37_, r_453__36_, r_453__35_, r_453__34_, r_453__33_, r_453__32_, r_453__31_, r_453__30_, r_453__29_, r_453__28_, r_453__27_, r_453__26_, r_453__25_, r_453__24_, r_453__23_, r_453__22_, r_453__21_, r_453__20_, r_453__19_, r_453__18_, r_453__17_, r_453__16_, r_453__15_, r_453__14_, r_453__13_, r_453__12_, r_453__11_, r_453__10_, r_453__9_, r_453__8_, r_453__7_, r_453__6_, r_453__5_, r_453__4_, r_453__3_, r_453__2_, r_453__1_, r_453__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N905)? data_i : 1'b0;
  assign N904 = sel_i[904];
  assign N905 = N3288;
  assign { r_n_453__63_, r_n_453__62_, r_n_453__61_, r_n_453__60_, r_n_453__59_, r_n_453__58_, r_n_453__57_, r_n_453__56_, r_n_453__55_, r_n_453__54_, r_n_453__53_, r_n_453__52_, r_n_453__51_, r_n_453__50_, r_n_453__49_, r_n_453__48_, r_n_453__47_, r_n_453__46_, r_n_453__45_, r_n_453__44_, r_n_453__43_, r_n_453__42_, r_n_453__41_, r_n_453__40_, r_n_453__39_, r_n_453__38_, r_n_453__37_, r_n_453__36_, r_n_453__35_, r_n_453__34_, r_n_453__33_, r_n_453__32_, r_n_453__31_, r_n_453__30_, r_n_453__29_, r_n_453__28_, r_n_453__27_, r_n_453__26_, r_n_453__25_, r_n_453__24_, r_n_453__23_, r_n_453__22_, r_n_453__21_, r_n_453__20_, r_n_453__19_, r_n_453__18_, r_n_453__17_, r_n_453__16_, r_n_453__15_, r_n_453__14_, r_n_453__13_, r_n_453__12_, r_n_453__11_, r_n_453__10_, r_n_453__9_, r_n_453__8_, r_n_453__7_, r_n_453__6_, r_n_453__5_, r_n_453__4_, r_n_453__3_, r_n_453__2_, r_n_453__1_, r_n_453__0_ } = (N906)? { r_454__63_, r_454__62_, r_454__61_, r_454__60_, r_454__59_, r_454__58_, r_454__57_, r_454__56_, r_454__55_, r_454__54_, r_454__53_, r_454__52_, r_454__51_, r_454__50_, r_454__49_, r_454__48_, r_454__47_, r_454__46_, r_454__45_, r_454__44_, r_454__43_, r_454__42_, r_454__41_, r_454__40_, r_454__39_, r_454__38_, r_454__37_, r_454__36_, r_454__35_, r_454__34_, r_454__33_, r_454__32_, r_454__31_, r_454__30_, r_454__29_, r_454__28_, r_454__27_, r_454__26_, r_454__25_, r_454__24_, r_454__23_, r_454__22_, r_454__21_, r_454__20_, r_454__19_, r_454__18_, r_454__17_, r_454__16_, r_454__15_, r_454__14_, r_454__13_, r_454__12_, r_454__11_, r_454__10_, r_454__9_, r_454__8_, r_454__7_, r_454__6_, r_454__5_, r_454__4_, r_454__3_, r_454__2_, r_454__1_, r_454__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N907)? data_i : 1'b0;
  assign N906 = sel_i[906];
  assign N907 = N3293;
  assign { r_n_454__63_, r_n_454__62_, r_n_454__61_, r_n_454__60_, r_n_454__59_, r_n_454__58_, r_n_454__57_, r_n_454__56_, r_n_454__55_, r_n_454__54_, r_n_454__53_, r_n_454__52_, r_n_454__51_, r_n_454__50_, r_n_454__49_, r_n_454__48_, r_n_454__47_, r_n_454__46_, r_n_454__45_, r_n_454__44_, r_n_454__43_, r_n_454__42_, r_n_454__41_, r_n_454__40_, r_n_454__39_, r_n_454__38_, r_n_454__37_, r_n_454__36_, r_n_454__35_, r_n_454__34_, r_n_454__33_, r_n_454__32_, r_n_454__31_, r_n_454__30_, r_n_454__29_, r_n_454__28_, r_n_454__27_, r_n_454__26_, r_n_454__25_, r_n_454__24_, r_n_454__23_, r_n_454__22_, r_n_454__21_, r_n_454__20_, r_n_454__19_, r_n_454__18_, r_n_454__17_, r_n_454__16_, r_n_454__15_, r_n_454__14_, r_n_454__13_, r_n_454__12_, r_n_454__11_, r_n_454__10_, r_n_454__9_, r_n_454__8_, r_n_454__7_, r_n_454__6_, r_n_454__5_, r_n_454__4_, r_n_454__3_, r_n_454__2_, r_n_454__1_, r_n_454__0_ } = (N908)? { r_455__63_, r_455__62_, r_455__61_, r_455__60_, r_455__59_, r_455__58_, r_455__57_, r_455__56_, r_455__55_, r_455__54_, r_455__53_, r_455__52_, r_455__51_, r_455__50_, r_455__49_, r_455__48_, r_455__47_, r_455__46_, r_455__45_, r_455__44_, r_455__43_, r_455__42_, r_455__41_, r_455__40_, r_455__39_, r_455__38_, r_455__37_, r_455__36_, r_455__35_, r_455__34_, r_455__33_, r_455__32_, r_455__31_, r_455__30_, r_455__29_, r_455__28_, r_455__27_, r_455__26_, r_455__25_, r_455__24_, r_455__23_, r_455__22_, r_455__21_, r_455__20_, r_455__19_, r_455__18_, r_455__17_, r_455__16_, r_455__15_, r_455__14_, r_455__13_, r_455__12_, r_455__11_, r_455__10_, r_455__9_, r_455__8_, r_455__7_, r_455__6_, r_455__5_, r_455__4_, r_455__3_, r_455__2_, r_455__1_, r_455__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N909)? data_i : 1'b0;
  assign N908 = sel_i[908];
  assign N909 = N3298;
  assign { r_n_455__63_, r_n_455__62_, r_n_455__61_, r_n_455__60_, r_n_455__59_, r_n_455__58_, r_n_455__57_, r_n_455__56_, r_n_455__55_, r_n_455__54_, r_n_455__53_, r_n_455__52_, r_n_455__51_, r_n_455__50_, r_n_455__49_, r_n_455__48_, r_n_455__47_, r_n_455__46_, r_n_455__45_, r_n_455__44_, r_n_455__43_, r_n_455__42_, r_n_455__41_, r_n_455__40_, r_n_455__39_, r_n_455__38_, r_n_455__37_, r_n_455__36_, r_n_455__35_, r_n_455__34_, r_n_455__33_, r_n_455__32_, r_n_455__31_, r_n_455__30_, r_n_455__29_, r_n_455__28_, r_n_455__27_, r_n_455__26_, r_n_455__25_, r_n_455__24_, r_n_455__23_, r_n_455__22_, r_n_455__21_, r_n_455__20_, r_n_455__19_, r_n_455__18_, r_n_455__17_, r_n_455__16_, r_n_455__15_, r_n_455__14_, r_n_455__13_, r_n_455__12_, r_n_455__11_, r_n_455__10_, r_n_455__9_, r_n_455__8_, r_n_455__7_, r_n_455__6_, r_n_455__5_, r_n_455__4_, r_n_455__3_, r_n_455__2_, r_n_455__1_, r_n_455__0_ } = (N910)? { r_456__63_, r_456__62_, r_456__61_, r_456__60_, r_456__59_, r_456__58_, r_456__57_, r_456__56_, r_456__55_, r_456__54_, r_456__53_, r_456__52_, r_456__51_, r_456__50_, r_456__49_, r_456__48_, r_456__47_, r_456__46_, r_456__45_, r_456__44_, r_456__43_, r_456__42_, r_456__41_, r_456__40_, r_456__39_, r_456__38_, r_456__37_, r_456__36_, r_456__35_, r_456__34_, r_456__33_, r_456__32_, r_456__31_, r_456__30_, r_456__29_, r_456__28_, r_456__27_, r_456__26_, r_456__25_, r_456__24_, r_456__23_, r_456__22_, r_456__21_, r_456__20_, r_456__19_, r_456__18_, r_456__17_, r_456__16_, r_456__15_, r_456__14_, r_456__13_, r_456__12_, r_456__11_, r_456__10_, r_456__9_, r_456__8_, r_456__7_, r_456__6_, r_456__5_, r_456__4_, r_456__3_, r_456__2_, r_456__1_, r_456__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N911)? data_i : 1'b0;
  assign N910 = sel_i[910];
  assign N911 = N3303;
  assign { r_n_456__63_, r_n_456__62_, r_n_456__61_, r_n_456__60_, r_n_456__59_, r_n_456__58_, r_n_456__57_, r_n_456__56_, r_n_456__55_, r_n_456__54_, r_n_456__53_, r_n_456__52_, r_n_456__51_, r_n_456__50_, r_n_456__49_, r_n_456__48_, r_n_456__47_, r_n_456__46_, r_n_456__45_, r_n_456__44_, r_n_456__43_, r_n_456__42_, r_n_456__41_, r_n_456__40_, r_n_456__39_, r_n_456__38_, r_n_456__37_, r_n_456__36_, r_n_456__35_, r_n_456__34_, r_n_456__33_, r_n_456__32_, r_n_456__31_, r_n_456__30_, r_n_456__29_, r_n_456__28_, r_n_456__27_, r_n_456__26_, r_n_456__25_, r_n_456__24_, r_n_456__23_, r_n_456__22_, r_n_456__21_, r_n_456__20_, r_n_456__19_, r_n_456__18_, r_n_456__17_, r_n_456__16_, r_n_456__15_, r_n_456__14_, r_n_456__13_, r_n_456__12_, r_n_456__11_, r_n_456__10_, r_n_456__9_, r_n_456__8_, r_n_456__7_, r_n_456__6_, r_n_456__5_, r_n_456__4_, r_n_456__3_, r_n_456__2_, r_n_456__1_, r_n_456__0_ } = (N912)? { r_457__63_, r_457__62_, r_457__61_, r_457__60_, r_457__59_, r_457__58_, r_457__57_, r_457__56_, r_457__55_, r_457__54_, r_457__53_, r_457__52_, r_457__51_, r_457__50_, r_457__49_, r_457__48_, r_457__47_, r_457__46_, r_457__45_, r_457__44_, r_457__43_, r_457__42_, r_457__41_, r_457__40_, r_457__39_, r_457__38_, r_457__37_, r_457__36_, r_457__35_, r_457__34_, r_457__33_, r_457__32_, r_457__31_, r_457__30_, r_457__29_, r_457__28_, r_457__27_, r_457__26_, r_457__25_, r_457__24_, r_457__23_, r_457__22_, r_457__21_, r_457__20_, r_457__19_, r_457__18_, r_457__17_, r_457__16_, r_457__15_, r_457__14_, r_457__13_, r_457__12_, r_457__11_, r_457__10_, r_457__9_, r_457__8_, r_457__7_, r_457__6_, r_457__5_, r_457__4_, r_457__3_, r_457__2_, r_457__1_, r_457__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N913)? data_i : 1'b0;
  assign N912 = sel_i[912];
  assign N913 = N3308;
  assign { r_n_457__63_, r_n_457__62_, r_n_457__61_, r_n_457__60_, r_n_457__59_, r_n_457__58_, r_n_457__57_, r_n_457__56_, r_n_457__55_, r_n_457__54_, r_n_457__53_, r_n_457__52_, r_n_457__51_, r_n_457__50_, r_n_457__49_, r_n_457__48_, r_n_457__47_, r_n_457__46_, r_n_457__45_, r_n_457__44_, r_n_457__43_, r_n_457__42_, r_n_457__41_, r_n_457__40_, r_n_457__39_, r_n_457__38_, r_n_457__37_, r_n_457__36_, r_n_457__35_, r_n_457__34_, r_n_457__33_, r_n_457__32_, r_n_457__31_, r_n_457__30_, r_n_457__29_, r_n_457__28_, r_n_457__27_, r_n_457__26_, r_n_457__25_, r_n_457__24_, r_n_457__23_, r_n_457__22_, r_n_457__21_, r_n_457__20_, r_n_457__19_, r_n_457__18_, r_n_457__17_, r_n_457__16_, r_n_457__15_, r_n_457__14_, r_n_457__13_, r_n_457__12_, r_n_457__11_, r_n_457__10_, r_n_457__9_, r_n_457__8_, r_n_457__7_, r_n_457__6_, r_n_457__5_, r_n_457__4_, r_n_457__3_, r_n_457__2_, r_n_457__1_, r_n_457__0_ } = (N914)? { r_458__63_, r_458__62_, r_458__61_, r_458__60_, r_458__59_, r_458__58_, r_458__57_, r_458__56_, r_458__55_, r_458__54_, r_458__53_, r_458__52_, r_458__51_, r_458__50_, r_458__49_, r_458__48_, r_458__47_, r_458__46_, r_458__45_, r_458__44_, r_458__43_, r_458__42_, r_458__41_, r_458__40_, r_458__39_, r_458__38_, r_458__37_, r_458__36_, r_458__35_, r_458__34_, r_458__33_, r_458__32_, r_458__31_, r_458__30_, r_458__29_, r_458__28_, r_458__27_, r_458__26_, r_458__25_, r_458__24_, r_458__23_, r_458__22_, r_458__21_, r_458__20_, r_458__19_, r_458__18_, r_458__17_, r_458__16_, r_458__15_, r_458__14_, r_458__13_, r_458__12_, r_458__11_, r_458__10_, r_458__9_, r_458__8_, r_458__7_, r_458__6_, r_458__5_, r_458__4_, r_458__3_, r_458__2_, r_458__1_, r_458__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N915)? data_i : 1'b0;
  assign N914 = sel_i[914];
  assign N915 = N3313;
  assign { r_n_458__63_, r_n_458__62_, r_n_458__61_, r_n_458__60_, r_n_458__59_, r_n_458__58_, r_n_458__57_, r_n_458__56_, r_n_458__55_, r_n_458__54_, r_n_458__53_, r_n_458__52_, r_n_458__51_, r_n_458__50_, r_n_458__49_, r_n_458__48_, r_n_458__47_, r_n_458__46_, r_n_458__45_, r_n_458__44_, r_n_458__43_, r_n_458__42_, r_n_458__41_, r_n_458__40_, r_n_458__39_, r_n_458__38_, r_n_458__37_, r_n_458__36_, r_n_458__35_, r_n_458__34_, r_n_458__33_, r_n_458__32_, r_n_458__31_, r_n_458__30_, r_n_458__29_, r_n_458__28_, r_n_458__27_, r_n_458__26_, r_n_458__25_, r_n_458__24_, r_n_458__23_, r_n_458__22_, r_n_458__21_, r_n_458__20_, r_n_458__19_, r_n_458__18_, r_n_458__17_, r_n_458__16_, r_n_458__15_, r_n_458__14_, r_n_458__13_, r_n_458__12_, r_n_458__11_, r_n_458__10_, r_n_458__9_, r_n_458__8_, r_n_458__7_, r_n_458__6_, r_n_458__5_, r_n_458__4_, r_n_458__3_, r_n_458__2_, r_n_458__1_, r_n_458__0_ } = (N916)? { r_459__63_, r_459__62_, r_459__61_, r_459__60_, r_459__59_, r_459__58_, r_459__57_, r_459__56_, r_459__55_, r_459__54_, r_459__53_, r_459__52_, r_459__51_, r_459__50_, r_459__49_, r_459__48_, r_459__47_, r_459__46_, r_459__45_, r_459__44_, r_459__43_, r_459__42_, r_459__41_, r_459__40_, r_459__39_, r_459__38_, r_459__37_, r_459__36_, r_459__35_, r_459__34_, r_459__33_, r_459__32_, r_459__31_, r_459__30_, r_459__29_, r_459__28_, r_459__27_, r_459__26_, r_459__25_, r_459__24_, r_459__23_, r_459__22_, r_459__21_, r_459__20_, r_459__19_, r_459__18_, r_459__17_, r_459__16_, r_459__15_, r_459__14_, r_459__13_, r_459__12_, r_459__11_, r_459__10_, r_459__9_, r_459__8_, r_459__7_, r_459__6_, r_459__5_, r_459__4_, r_459__3_, r_459__2_, r_459__1_, r_459__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N917)? data_i : 1'b0;
  assign N916 = sel_i[916];
  assign N917 = N3318;
  assign { r_n_459__63_, r_n_459__62_, r_n_459__61_, r_n_459__60_, r_n_459__59_, r_n_459__58_, r_n_459__57_, r_n_459__56_, r_n_459__55_, r_n_459__54_, r_n_459__53_, r_n_459__52_, r_n_459__51_, r_n_459__50_, r_n_459__49_, r_n_459__48_, r_n_459__47_, r_n_459__46_, r_n_459__45_, r_n_459__44_, r_n_459__43_, r_n_459__42_, r_n_459__41_, r_n_459__40_, r_n_459__39_, r_n_459__38_, r_n_459__37_, r_n_459__36_, r_n_459__35_, r_n_459__34_, r_n_459__33_, r_n_459__32_, r_n_459__31_, r_n_459__30_, r_n_459__29_, r_n_459__28_, r_n_459__27_, r_n_459__26_, r_n_459__25_, r_n_459__24_, r_n_459__23_, r_n_459__22_, r_n_459__21_, r_n_459__20_, r_n_459__19_, r_n_459__18_, r_n_459__17_, r_n_459__16_, r_n_459__15_, r_n_459__14_, r_n_459__13_, r_n_459__12_, r_n_459__11_, r_n_459__10_, r_n_459__9_, r_n_459__8_, r_n_459__7_, r_n_459__6_, r_n_459__5_, r_n_459__4_, r_n_459__3_, r_n_459__2_, r_n_459__1_, r_n_459__0_ } = (N918)? { r_460__63_, r_460__62_, r_460__61_, r_460__60_, r_460__59_, r_460__58_, r_460__57_, r_460__56_, r_460__55_, r_460__54_, r_460__53_, r_460__52_, r_460__51_, r_460__50_, r_460__49_, r_460__48_, r_460__47_, r_460__46_, r_460__45_, r_460__44_, r_460__43_, r_460__42_, r_460__41_, r_460__40_, r_460__39_, r_460__38_, r_460__37_, r_460__36_, r_460__35_, r_460__34_, r_460__33_, r_460__32_, r_460__31_, r_460__30_, r_460__29_, r_460__28_, r_460__27_, r_460__26_, r_460__25_, r_460__24_, r_460__23_, r_460__22_, r_460__21_, r_460__20_, r_460__19_, r_460__18_, r_460__17_, r_460__16_, r_460__15_, r_460__14_, r_460__13_, r_460__12_, r_460__11_, r_460__10_, r_460__9_, r_460__8_, r_460__7_, r_460__6_, r_460__5_, r_460__4_, r_460__3_, r_460__2_, r_460__1_, r_460__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N919)? data_i : 1'b0;
  assign N918 = sel_i[918];
  assign N919 = N3323;
  assign { r_n_460__63_, r_n_460__62_, r_n_460__61_, r_n_460__60_, r_n_460__59_, r_n_460__58_, r_n_460__57_, r_n_460__56_, r_n_460__55_, r_n_460__54_, r_n_460__53_, r_n_460__52_, r_n_460__51_, r_n_460__50_, r_n_460__49_, r_n_460__48_, r_n_460__47_, r_n_460__46_, r_n_460__45_, r_n_460__44_, r_n_460__43_, r_n_460__42_, r_n_460__41_, r_n_460__40_, r_n_460__39_, r_n_460__38_, r_n_460__37_, r_n_460__36_, r_n_460__35_, r_n_460__34_, r_n_460__33_, r_n_460__32_, r_n_460__31_, r_n_460__30_, r_n_460__29_, r_n_460__28_, r_n_460__27_, r_n_460__26_, r_n_460__25_, r_n_460__24_, r_n_460__23_, r_n_460__22_, r_n_460__21_, r_n_460__20_, r_n_460__19_, r_n_460__18_, r_n_460__17_, r_n_460__16_, r_n_460__15_, r_n_460__14_, r_n_460__13_, r_n_460__12_, r_n_460__11_, r_n_460__10_, r_n_460__9_, r_n_460__8_, r_n_460__7_, r_n_460__6_, r_n_460__5_, r_n_460__4_, r_n_460__3_, r_n_460__2_, r_n_460__1_, r_n_460__0_ } = (N920)? { r_461__63_, r_461__62_, r_461__61_, r_461__60_, r_461__59_, r_461__58_, r_461__57_, r_461__56_, r_461__55_, r_461__54_, r_461__53_, r_461__52_, r_461__51_, r_461__50_, r_461__49_, r_461__48_, r_461__47_, r_461__46_, r_461__45_, r_461__44_, r_461__43_, r_461__42_, r_461__41_, r_461__40_, r_461__39_, r_461__38_, r_461__37_, r_461__36_, r_461__35_, r_461__34_, r_461__33_, r_461__32_, r_461__31_, r_461__30_, r_461__29_, r_461__28_, r_461__27_, r_461__26_, r_461__25_, r_461__24_, r_461__23_, r_461__22_, r_461__21_, r_461__20_, r_461__19_, r_461__18_, r_461__17_, r_461__16_, r_461__15_, r_461__14_, r_461__13_, r_461__12_, r_461__11_, r_461__10_, r_461__9_, r_461__8_, r_461__7_, r_461__6_, r_461__5_, r_461__4_, r_461__3_, r_461__2_, r_461__1_, r_461__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N921)? data_i : 1'b0;
  assign N920 = sel_i[920];
  assign N921 = N3328;
  assign { r_n_461__63_, r_n_461__62_, r_n_461__61_, r_n_461__60_, r_n_461__59_, r_n_461__58_, r_n_461__57_, r_n_461__56_, r_n_461__55_, r_n_461__54_, r_n_461__53_, r_n_461__52_, r_n_461__51_, r_n_461__50_, r_n_461__49_, r_n_461__48_, r_n_461__47_, r_n_461__46_, r_n_461__45_, r_n_461__44_, r_n_461__43_, r_n_461__42_, r_n_461__41_, r_n_461__40_, r_n_461__39_, r_n_461__38_, r_n_461__37_, r_n_461__36_, r_n_461__35_, r_n_461__34_, r_n_461__33_, r_n_461__32_, r_n_461__31_, r_n_461__30_, r_n_461__29_, r_n_461__28_, r_n_461__27_, r_n_461__26_, r_n_461__25_, r_n_461__24_, r_n_461__23_, r_n_461__22_, r_n_461__21_, r_n_461__20_, r_n_461__19_, r_n_461__18_, r_n_461__17_, r_n_461__16_, r_n_461__15_, r_n_461__14_, r_n_461__13_, r_n_461__12_, r_n_461__11_, r_n_461__10_, r_n_461__9_, r_n_461__8_, r_n_461__7_, r_n_461__6_, r_n_461__5_, r_n_461__4_, r_n_461__3_, r_n_461__2_, r_n_461__1_, r_n_461__0_ } = (N922)? { r_462__63_, r_462__62_, r_462__61_, r_462__60_, r_462__59_, r_462__58_, r_462__57_, r_462__56_, r_462__55_, r_462__54_, r_462__53_, r_462__52_, r_462__51_, r_462__50_, r_462__49_, r_462__48_, r_462__47_, r_462__46_, r_462__45_, r_462__44_, r_462__43_, r_462__42_, r_462__41_, r_462__40_, r_462__39_, r_462__38_, r_462__37_, r_462__36_, r_462__35_, r_462__34_, r_462__33_, r_462__32_, r_462__31_, r_462__30_, r_462__29_, r_462__28_, r_462__27_, r_462__26_, r_462__25_, r_462__24_, r_462__23_, r_462__22_, r_462__21_, r_462__20_, r_462__19_, r_462__18_, r_462__17_, r_462__16_, r_462__15_, r_462__14_, r_462__13_, r_462__12_, r_462__11_, r_462__10_, r_462__9_, r_462__8_, r_462__7_, r_462__6_, r_462__5_, r_462__4_, r_462__3_, r_462__2_, r_462__1_, r_462__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N923)? data_i : 1'b0;
  assign N922 = sel_i[922];
  assign N923 = N3333;
  assign { r_n_462__63_, r_n_462__62_, r_n_462__61_, r_n_462__60_, r_n_462__59_, r_n_462__58_, r_n_462__57_, r_n_462__56_, r_n_462__55_, r_n_462__54_, r_n_462__53_, r_n_462__52_, r_n_462__51_, r_n_462__50_, r_n_462__49_, r_n_462__48_, r_n_462__47_, r_n_462__46_, r_n_462__45_, r_n_462__44_, r_n_462__43_, r_n_462__42_, r_n_462__41_, r_n_462__40_, r_n_462__39_, r_n_462__38_, r_n_462__37_, r_n_462__36_, r_n_462__35_, r_n_462__34_, r_n_462__33_, r_n_462__32_, r_n_462__31_, r_n_462__30_, r_n_462__29_, r_n_462__28_, r_n_462__27_, r_n_462__26_, r_n_462__25_, r_n_462__24_, r_n_462__23_, r_n_462__22_, r_n_462__21_, r_n_462__20_, r_n_462__19_, r_n_462__18_, r_n_462__17_, r_n_462__16_, r_n_462__15_, r_n_462__14_, r_n_462__13_, r_n_462__12_, r_n_462__11_, r_n_462__10_, r_n_462__9_, r_n_462__8_, r_n_462__7_, r_n_462__6_, r_n_462__5_, r_n_462__4_, r_n_462__3_, r_n_462__2_, r_n_462__1_, r_n_462__0_ } = (N924)? { r_463__63_, r_463__62_, r_463__61_, r_463__60_, r_463__59_, r_463__58_, r_463__57_, r_463__56_, r_463__55_, r_463__54_, r_463__53_, r_463__52_, r_463__51_, r_463__50_, r_463__49_, r_463__48_, r_463__47_, r_463__46_, r_463__45_, r_463__44_, r_463__43_, r_463__42_, r_463__41_, r_463__40_, r_463__39_, r_463__38_, r_463__37_, r_463__36_, r_463__35_, r_463__34_, r_463__33_, r_463__32_, r_463__31_, r_463__30_, r_463__29_, r_463__28_, r_463__27_, r_463__26_, r_463__25_, r_463__24_, r_463__23_, r_463__22_, r_463__21_, r_463__20_, r_463__19_, r_463__18_, r_463__17_, r_463__16_, r_463__15_, r_463__14_, r_463__13_, r_463__12_, r_463__11_, r_463__10_, r_463__9_, r_463__8_, r_463__7_, r_463__6_, r_463__5_, r_463__4_, r_463__3_, r_463__2_, r_463__1_, r_463__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N925)? data_i : 1'b0;
  assign N924 = sel_i[924];
  assign N925 = N3338;
  assign { r_n_463__63_, r_n_463__62_, r_n_463__61_, r_n_463__60_, r_n_463__59_, r_n_463__58_, r_n_463__57_, r_n_463__56_, r_n_463__55_, r_n_463__54_, r_n_463__53_, r_n_463__52_, r_n_463__51_, r_n_463__50_, r_n_463__49_, r_n_463__48_, r_n_463__47_, r_n_463__46_, r_n_463__45_, r_n_463__44_, r_n_463__43_, r_n_463__42_, r_n_463__41_, r_n_463__40_, r_n_463__39_, r_n_463__38_, r_n_463__37_, r_n_463__36_, r_n_463__35_, r_n_463__34_, r_n_463__33_, r_n_463__32_, r_n_463__31_, r_n_463__30_, r_n_463__29_, r_n_463__28_, r_n_463__27_, r_n_463__26_, r_n_463__25_, r_n_463__24_, r_n_463__23_, r_n_463__22_, r_n_463__21_, r_n_463__20_, r_n_463__19_, r_n_463__18_, r_n_463__17_, r_n_463__16_, r_n_463__15_, r_n_463__14_, r_n_463__13_, r_n_463__12_, r_n_463__11_, r_n_463__10_, r_n_463__9_, r_n_463__8_, r_n_463__7_, r_n_463__6_, r_n_463__5_, r_n_463__4_, r_n_463__3_, r_n_463__2_, r_n_463__1_, r_n_463__0_ } = (N926)? { r_464__63_, r_464__62_, r_464__61_, r_464__60_, r_464__59_, r_464__58_, r_464__57_, r_464__56_, r_464__55_, r_464__54_, r_464__53_, r_464__52_, r_464__51_, r_464__50_, r_464__49_, r_464__48_, r_464__47_, r_464__46_, r_464__45_, r_464__44_, r_464__43_, r_464__42_, r_464__41_, r_464__40_, r_464__39_, r_464__38_, r_464__37_, r_464__36_, r_464__35_, r_464__34_, r_464__33_, r_464__32_, r_464__31_, r_464__30_, r_464__29_, r_464__28_, r_464__27_, r_464__26_, r_464__25_, r_464__24_, r_464__23_, r_464__22_, r_464__21_, r_464__20_, r_464__19_, r_464__18_, r_464__17_, r_464__16_, r_464__15_, r_464__14_, r_464__13_, r_464__12_, r_464__11_, r_464__10_, r_464__9_, r_464__8_, r_464__7_, r_464__6_, r_464__5_, r_464__4_, r_464__3_, r_464__2_, r_464__1_, r_464__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N927)? data_i : 1'b0;
  assign N926 = sel_i[926];
  assign N927 = N3343;
  assign { r_n_464__63_, r_n_464__62_, r_n_464__61_, r_n_464__60_, r_n_464__59_, r_n_464__58_, r_n_464__57_, r_n_464__56_, r_n_464__55_, r_n_464__54_, r_n_464__53_, r_n_464__52_, r_n_464__51_, r_n_464__50_, r_n_464__49_, r_n_464__48_, r_n_464__47_, r_n_464__46_, r_n_464__45_, r_n_464__44_, r_n_464__43_, r_n_464__42_, r_n_464__41_, r_n_464__40_, r_n_464__39_, r_n_464__38_, r_n_464__37_, r_n_464__36_, r_n_464__35_, r_n_464__34_, r_n_464__33_, r_n_464__32_, r_n_464__31_, r_n_464__30_, r_n_464__29_, r_n_464__28_, r_n_464__27_, r_n_464__26_, r_n_464__25_, r_n_464__24_, r_n_464__23_, r_n_464__22_, r_n_464__21_, r_n_464__20_, r_n_464__19_, r_n_464__18_, r_n_464__17_, r_n_464__16_, r_n_464__15_, r_n_464__14_, r_n_464__13_, r_n_464__12_, r_n_464__11_, r_n_464__10_, r_n_464__9_, r_n_464__8_, r_n_464__7_, r_n_464__6_, r_n_464__5_, r_n_464__4_, r_n_464__3_, r_n_464__2_, r_n_464__1_, r_n_464__0_ } = (N928)? { r_465__63_, r_465__62_, r_465__61_, r_465__60_, r_465__59_, r_465__58_, r_465__57_, r_465__56_, r_465__55_, r_465__54_, r_465__53_, r_465__52_, r_465__51_, r_465__50_, r_465__49_, r_465__48_, r_465__47_, r_465__46_, r_465__45_, r_465__44_, r_465__43_, r_465__42_, r_465__41_, r_465__40_, r_465__39_, r_465__38_, r_465__37_, r_465__36_, r_465__35_, r_465__34_, r_465__33_, r_465__32_, r_465__31_, r_465__30_, r_465__29_, r_465__28_, r_465__27_, r_465__26_, r_465__25_, r_465__24_, r_465__23_, r_465__22_, r_465__21_, r_465__20_, r_465__19_, r_465__18_, r_465__17_, r_465__16_, r_465__15_, r_465__14_, r_465__13_, r_465__12_, r_465__11_, r_465__10_, r_465__9_, r_465__8_, r_465__7_, r_465__6_, r_465__5_, r_465__4_, r_465__3_, r_465__2_, r_465__1_, r_465__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N929)? data_i : 1'b0;
  assign N928 = sel_i[928];
  assign N929 = N3348;
  assign { r_n_465__63_, r_n_465__62_, r_n_465__61_, r_n_465__60_, r_n_465__59_, r_n_465__58_, r_n_465__57_, r_n_465__56_, r_n_465__55_, r_n_465__54_, r_n_465__53_, r_n_465__52_, r_n_465__51_, r_n_465__50_, r_n_465__49_, r_n_465__48_, r_n_465__47_, r_n_465__46_, r_n_465__45_, r_n_465__44_, r_n_465__43_, r_n_465__42_, r_n_465__41_, r_n_465__40_, r_n_465__39_, r_n_465__38_, r_n_465__37_, r_n_465__36_, r_n_465__35_, r_n_465__34_, r_n_465__33_, r_n_465__32_, r_n_465__31_, r_n_465__30_, r_n_465__29_, r_n_465__28_, r_n_465__27_, r_n_465__26_, r_n_465__25_, r_n_465__24_, r_n_465__23_, r_n_465__22_, r_n_465__21_, r_n_465__20_, r_n_465__19_, r_n_465__18_, r_n_465__17_, r_n_465__16_, r_n_465__15_, r_n_465__14_, r_n_465__13_, r_n_465__12_, r_n_465__11_, r_n_465__10_, r_n_465__9_, r_n_465__8_, r_n_465__7_, r_n_465__6_, r_n_465__5_, r_n_465__4_, r_n_465__3_, r_n_465__2_, r_n_465__1_, r_n_465__0_ } = (N930)? { r_466__63_, r_466__62_, r_466__61_, r_466__60_, r_466__59_, r_466__58_, r_466__57_, r_466__56_, r_466__55_, r_466__54_, r_466__53_, r_466__52_, r_466__51_, r_466__50_, r_466__49_, r_466__48_, r_466__47_, r_466__46_, r_466__45_, r_466__44_, r_466__43_, r_466__42_, r_466__41_, r_466__40_, r_466__39_, r_466__38_, r_466__37_, r_466__36_, r_466__35_, r_466__34_, r_466__33_, r_466__32_, r_466__31_, r_466__30_, r_466__29_, r_466__28_, r_466__27_, r_466__26_, r_466__25_, r_466__24_, r_466__23_, r_466__22_, r_466__21_, r_466__20_, r_466__19_, r_466__18_, r_466__17_, r_466__16_, r_466__15_, r_466__14_, r_466__13_, r_466__12_, r_466__11_, r_466__10_, r_466__9_, r_466__8_, r_466__7_, r_466__6_, r_466__5_, r_466__4_, r_466__3_, r_466__2_, r_466__1_, r_466__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N931)? data_i : 1'b0;
  assign N930 = sel_i[930];
  assign N931 = N3353;
  assign { r_n_466__63_, r_n_466__62_, r_n_466__61_, r_n_466__60_, r_n_466__59_, r_n_466__58_, r_n_466__57_, r_n_466__56_, r_n_466__55_, r_n_466__54_, r_n_466__53_, r_n_466__52_, r_n_466__51_, r_n_466__50_, r_n_466__49_, r_n_466__48_, r_n_466__47_, r_n_466__46_, r_n_466__45_, r_n_466__44_, r_n_466__43_, r_n_466__42_, r_n_466__41_, r_n_466__40_, r_n_466__39_, r_n_466__38_, r_n_466__37_, r_n_466__36_, r_n_466__35_, r_n_466__34_, r_n_466__33_, r_n_466__32_, r_n_466__31_, r_n_466__30_, r_n_466__29_, r_n_466__28_, r_n_466__27_, r_n_466__26_, r_n_466__25_, r_n_466__24_, r_n_466__23_, r_n_466__22_, r_n_466__21_, r_n_466__20_, r_n_466__19_, r_n_466__18_, r_n_466__17_, r_n_466__16_, r_n_466__15_, r_n_466__14_, r_n_466__13_, r_n_466__12_, r_n_466__11_, r_n_466__10_, r_n_466__9_, r_n_466__8_, r_n_466__7_, r_n_466__6_, r_n_466__5_, r_n_466__4_, r_n_466__3_, r_n_466__2_, r_n_466__1_, r_n_466__0_ } = (N932)? { r_467__63_, r_467__62_, r_467__61_, r_467__60_, r_467__59_, r_467__58_, r_467__57_, r_467__56_, r_467__55_, r_467__54_, r_467__53_, r_467__52_, r_467__51_, r_467__50_, r_467__49_, r_467__48_, r_467__47_, r_467__46_, r_467__45_, r_467__44_, r_467__43_, r_467__42_, r_467__41_, r_467__40_, r_467__39_, r_467__38_, r_467__37_, r_467__36_, r_467__35_, r_467__34_, r_467__33_, r_467__32_, r_467__31_, r_467__30_, r_467__29_, r_467__28_, r_467__27_, r_467__26_, r_467__25_, r_467__24_, r_467__23_, r_467__22_, r_467__21_, r_467__20_, r_467__19_, r_467__18_, r_467__17_, r_467__16_, r_467__15_, r_467__14_, r_467__13_, r_467__12_, r_467__11_, r_467__10_, r_467__9_, r_467__8_, r_467__7_, r_467__6_, r_467__5_, r_467__4_, r_467__3_, r_467__2_, r_467__1_, r_467__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N933)? data_i : 1'b0;
  assign N932 = sel_i[932];
  assign N933 = N3358;
  assign { r_n_467__63_, r_n_467__62_, r_n_467__61_, r_n_467__60_, r_n_467__59_, r_n_467__58_, r_n_467__57_, r_n_467__56_, r_n_467__55_, r_n_467__54_, r_n_467__53_, r_n_467__52_, r_n_467__51_, r_n_467__50_, r_n_467__49_, r_n_467__48_, r_n_467__47_, r_n_467__46_, r_n_467__45_, r_n_467__44_, r_n_467__43_, r_n_467__42_, r_n_467__41_, r_n_467__40_, r_n_467__39_, r_n_467__38_, r_n_467__37_, r_n_467__36_, r_n_467__35_, r_n_467__34_, r_n_467__33_, r_n_467__32_, r_n_467__31_, r_n_467__30_, r_n_467__29_, r_n_467__28_, r_n_467__27_, r_n_467__26_, r_n_467__25_, r_n_467__24_, r_n_467__23_, r_n_467__22_, r_n_467__21_, r_n_467__20_, r_n_467__19_, r_n_467__18_, r_n_467__17_, r_n_467__16_, r_n_467__15_, r_n_467__14_, r_n_467__13_, r_n_467__12_, r_n_467__11_, r_n_467__10_, r_n_467__9_, r_n_467__8_, r_n_467__7_, r_n_467__6_, r_n_467__5_, r_n_467__4_, r_n_467__3_, r_n_467__2_, r_n_467__1_, r_n_467__0_ } = (N934)? { r_468__63_, r_468__62_, r_468__61_, r_468__60_, r_468__59_, r_468__58_, r_468__57_, r_468__56_, r_468__55_, r_468__54_, r_468__53_, r_468__52_, r_468__51_, r_468__50_, r_468__49_, r_468__48_, r_468__47_, r_468__46_, r_468__45_, r_468__44_, r_468__43_, r_468__42_, r_468__41_, r_468__40_, r_468__39_, r_468__38_, r_468__37_, r_468__36_, r_468__35_, r_468__34_, r_468__33_, r_468__32_, r_468__31_, r_468__30_, r_468__29_, r_468__28_, r_468__27_, r_468__26_, r_468__25_, r_468__24_, r_468__23_, r_468__22_, r_468__21_, r_468__20_, r_468__19_, r_468__18_, r_468__17_, r_468__16_, r_468__15_, r_468__14_, r_468__13_, r_468__12_, r_468__11_, r_468__10_, r_468__9_, r_468__8_, r_468__7_, r_468__6_, r_468__5_, r_468__4_, r_468__3_, r_468__2_, r_468__1_, r_468__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N935)? data_i : 1'b0;
  assign N934 = sel_i[934];
  assign N935 = N3363;
  assign { r_n_468__63_, r_n_468__62_, r_n_468__61_, r_n_468__60_, r_n_468__59_, r_n_468__58_, r_n_468__57_, r_n_468__56_, r_n_468__55_, r_n_468__54_, r_n_468__53_, r_n_468__52_, r_n_468__51_, r_n_468__50_, r_n_468__49_, r_n_468__48_, r_n_468__47_, r_n_468__46_, r_n_468__45_, r_n_468__44_, r_n_468__43_, r_n_468__42_, r_n_468__41_, r_n_468__40_, r_n_468__39_, r_n_468__38_, r_n_468__37_, r_n_468__36_, r_n_468__35_, r_n_468__34_, r_n_468__33_, r_n_468__32_, r_n_468__31_, r_n_468__30_, r_n_468__29_, r_n_468__28_, r_n_468__27_, r_n_468__26_, r_n_468__25_, r_n_468__24_, r_n_468__23_, r_n_468__22_, r_n_468__21_, r_n_468__20_, r_n_468__19_, r_n_468__18_, r_n_468__17_, r_n_468__16_, r_n_468__15_, r_n_468__14_, r_n_468__13_, r_n_468__12_, r_n_468__11_, r_n_468__10_, r_n_468__9_, r_n_468__8_, r_n_468__7_, r_n_468__6_, r_n_468__5_, r_n_468__4_, r_n_468__3_, r_n_468__2_, r_n_468__1_, r_n_468__0_ } = (N936)? { r_469__63_, r_469__62_, r_469__61_, r_469__60_, r_469__59_, r_469__58_, r_469__57_, r_469__56_, r_469__55_, r_469__54_, r_469__53_, r_469__52_, r_469__51_, r_469__50_, r_469__49_, r_469__48_, r_469__47_, r_469__46_, r_469__45_, r_469__44_, r_469__43_, r_469__42_, r_469__41_, r_469__40_, r_469__39_, r_469__38_, r_469__37_, r_469__36_, r_469__35_, r_469__34_, r_469__33_, r_469__32_, r_469__31_, r_469__30_, r_469__29_, r_469__28_, r_469__27_, r_469__26_, r_469__25_, r_469__24_, r_469__23_, r_469__22_, r_469__21_, r_469__20_, r_469__19_, r_469__18_, r_469__17_, r_469__16_, r_469__15_, r_469__14_, r_469__13_, r_469__12_, r_469__11_, r_469__10_, r_469__9_, r_469__8_, r_469__7_, r_469__6_, r_469__5_, r_469__4_, r_469__3_, r_469__2_, r_469__1_, r_469__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N937)? data_i : 1'b0;
  assign N936 = sel_i[936];
  assign N937 = N3368;
  assign { r_n_469__63_, r_n_469__62_, r_n_469__61_, r_n_469__60_, r_n_469__59_, r_n_469__58_, r_n_469__57_, r_n_469__56_, r_n_469__55_, r_n_469__54_, r_n_469__53_, r_n_469__52_, r_n_469__51_, r_n_469__50_, r_n_469__49_, r_n_469__48_, r_n_469__47_, r_n_469__46_, r_n_469__45_, r_n_469__44_, r_n_469__43_, r_n_469__42_, r_n_469__41_, r_n_469__40_, r_n_469__39_, r_n_469__38_, r_n_469__37_, r_n_469__36_, r_n_469__35_, r_n_469__34_, r_n_469__33_, r_n_469__32_, r_n_469__31_, r_n_469__30_, r_n_469__29_, r_n_469__28_, r_n_469__27_, r_n_469__26_, r_n_469__25_, r_n_469__24_, r_n_469__23_, r_n_469__22_, r_n_469__21_, r_n_469__20_, r_n_469__19_, r_n_469__18_, r_n_469__17_, r_n_469__16_, r_n_469__15_, r_n_469__14_, r_n_469__13_, r_n_469__12_, r_n_469__11_, r_n_469__10_, r_n_469__9_, r_n_469__8_, r_n_469__7_, r_n_469__6_, r_n_469__5_, r_n_469__4_, r_n_469__3_, r_n_469__2_, r_n_469__1_, r_n_469__0_ } = (N938)? { r_470__63_, r_470__62_, r_470__61_, r_470__60_, r_470__59_, r_470__58_, r_470__57_, r_470__56_, r_470__55_, r_470__54_, r_470__53_, r_470__52_, r_470__51_, r_470__50_, r_470__49_, r_470__48_, r_470__47_, r_470__46_, r_470__45_, r_470__44_, r_470__43_, r_470__42_, r_470__41_, r_470__40_, r_470__39_, r_470__38_, r_470__37_, r_470__36_, r_470__35_, r_470__34_, r_470__33_, r_470__32_, r_470__31_, r_470__30_, r_470__29_, r_470__28_, r_470__27_, r_470__26_, r_470__25_, r_470__24_, r_470__23_, r_470__22_, r_470__21_, r_470__20_, r_470__19_, r_470__18_, r_470__17_, r_470__16_, r_470__15_, r_470__14_, r_470__13_, r_470__12_, r_470__11_, r_470__10_, r_470__9_, r_470__8_, r_470__7_, r_470__6_, r_470__5_, r_470__4_, r_470__3_, r_470__2_, r_470__1_, r_470__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N939)? data_i : 1'b0;
  assign N938 = sel_i[938];
  assign N939 = N3373;
  assign { r_n_470__63_, r_n_470__62_, r_n_470__61_, r_n_470__60_, r_n_470__59_, r_n_470__58_, r_n_470__57_, r_n_470__56_, r_n_470__55_, r_n_470__54_, r_n_470__53_, r_n_470__52_, r_n_470__51_, r_n_470__50_, r_n_470__49_, r_n_470__48_, r_n_470__47_, r_n_470__46_, r_n_470__45_, r_n_470__44_, r_n_470__43_, r_n_470__42_, r_n_470__41_, r_n_470__40_, r_n_470__39_, r_n_470__38_, r_n_470__37_, r_n_470__36_, r_n_470__35_, r_n_470__34_, r_n_470__33_, r_n_470__32_, r_n_470__31_, r_n_470__30_, r_n_470__29_, r_n_470__28_, r_n_470__27_, r_n_470__26_, r_n_470__25_, r_n_470__24_, r_n_470__23_, r_n_470__22_, r_n_470__21_, r_n_470__20_, r_n_470__19_, r_n_470__18_, r_n_470__17_, r_n_470__16_, r_n_470__15_, r_n_470__14_, r_n_470__13_, r_n_470__12_, r_n_470__11_, r_n_470__10_, r_n_470__9_, r_n_470__8_, r_n_470__7_, r_n_470__6_, r_n_470__5_, r_n_470__4_, r_n_470__3_, r_n_470__2_, r_n_470__1_, r_n_470__0_ } = (N940)? { r_471__63_, r_471__62_, r_471__61_, r_471__60_, r_471__59_, r_471__58_, r_471__57_, r_471__56_, r_471__55_, r_471__54_, r_471__53_, r_471__52_, r_471__51_, r_471__50_, r_471__49_, r_471__48_, r_471__47_, r_471__46_, r_471__45_, r_471__44_, r_471__43_, r_471__42_, r_471__41_, r_471__40_, r_471__39_, r_471__38_, r_471__37_, r_471__36_, r_471__35_, r_471__34_, r_471__33_, r_471__32_, r_471__31_, r_471__30_, r_471__29_, r_471__28_, r_471__27_, r_471__26_, r_471__25_, r_471__24_, r_471__23_, r_471__22_, r_471__21_, r_471__20_, r_471__19_, r_471__18_, r_471__17_, r_471__16_, r_471__15_, r_471__14_, r_471__13_, r_471__12_, r_471__11_, r_471__10_, r_471__9_, r_471__8_, r_471__7_, r_471__6_, r_471__5_, r_471__4_, r_471__3_, r_471__2_, r_471__1_, r_471__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N941)? data_i : 1'b0;
  assign N940 = sel_i[940];
  assign N941 = N3378;
  assign { r_n_471__63_, r_n_471__62_, r_n_471__61_, r_n_471__60_, r_n_471__59_, r_n_471__58_, r_n_471__57_, r_n_471__56_, r_n_471__55_, r_n_471__54_, r_n_471__53_, r_n_471__52_, r_n_471__51_, r_n_471__50_, r_n_471__49_, r_n_471__48_, r_n_471__47_, r_n_471__46_, r_n_471__45_, r_n_471__44_, r_n_471__43_, r_n_471__42_, r_n_471__41_, r_n_471__40_, r_n_471__39_, r_n_471__38_, r_n_471__37_, r_n_471__36_, r_n_471__35_, r_n_471__34_, r_n_471__33_, r_n_471__32_, r_n_471__31_, r_n_471__30_, r_n_471__29_, r_n_471__28_, r_n_471__27_, r_n_471__26_, r_n_471__25_, r_n_471__24_, r_n_471__23_, r_n_471__22_, r_n_471__21_, r_n_471__20_, r_n_471__19_, r_n_471__18_, r_n_471__17_, r_n_471__16_, r_n_471__15_, r_n_471__14_, r_n_471__13_, r_n_471__12_, r_n_471__11_, r_n_471__10_, r_n_471__9_, r_n_471__8_, r_n_471__7_, r_n_471__6_, r_n_471__5_, r_n_471__4_, r_n_471__3_, r_n_471__2_, r_n_471__1_, r_n_471__0_ } = (N942)? { r_472__63_, r_472__62_, r_472__61_, r_472__60_, r_472__59_, r_472__58_, r_472__57_, r_472__56_, r_472__55_, r_472__54_, r_472__53_, r_472__52_, r_472__51_, r_472__50_, r_472__49_, r_472__48_, r_472__47_, r_472__46_, r_472__45_, r_472__44_, r_472__43_, r_472__42_, r_472__41_, r_472__40_, r_472__39_, r_472__38_, r_472__37_, r_472__36_, r_472__35_, r_472__34_, r_472__33_, r_472__32_, r_472__31_, r_472__30_, r_472__29_, r_472__28_, r_472__27_, r_472__26_, r_472__25_, r_472__24_, r_472__23_, r_472__22_, r_472__21_, r_472__20_, r_472__19_, r_472__18_, r_472__17_, r_472__16_, r_472__15_, r_472__14_, r_472__13_, r_472__12_, r_472__11_, r_472__10_, r_472__9_, r_472__8_, r_472__7_, r_472__6_, r_472__5_, r_472__4_, r_472__3_, r_472__2_, r_472__1_, r_472__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N943)? data_i : 1'b0;
  assign N942 = sel_i[942];
  assign N943 = N3383;
  assign { r_n_472__63_, r_n_472__62_, r_n_472__61_, r_n_472__60_, r_n_472__59_, r_n_472__58_, r_n_472__57_, r_n_472__56_, r_n_472__55_, r_n_472__54_, r_n_472__53_, r_n_472__52_, r_n_472__51_, r_n_472__50_, r_n_472__49_, r_n_472__48_, r_n_472__47_, r_n_472__46_, r_n_472__45_, r_n_472__44_, r_n_472__43_, r_n_472__42_, r_n_472__41_, r_n_472__40_, r_n_472__39_, r_n_472__38_, r_n_472__37_, r_n_472__36_, r_n_472__35_, r_n_472__34_, r_n_472__33_, r_n_472__32_, r_n_472__31_, r_n_472__30_, r_n_472__29_, r_n_472__28_, r_n_472__27_, r_n_472__26_, r_n_472__25_, r_n_472__24_, r_n_472__23_, r_n_472__22_, r_n_472__21_, r_n_472__20_, r_n_472__19_, r_n_472__18_, r_n_472__17_, r_n_472__16_, r_n_472__15_, r_n_472__14_, r_n_472__13_, r_n_472__12_, r_n_472__11_, r_n_472__10_, r_n_472__9_, r_n_472__8_, r_n_472__7_, r_n_472__6_, r_n_472__5_, r_n_472__4_, r_n_472__3_, r_n_472__2_, r_n_472__1_, r_n_472__0_ } = (N944)? { r_473__63_, r_473__62_, r_473__61_, r_473__60_, r_473__59_, r_473__58_, r_473__57_, r_473__56_, r_473__55_, r_473__54_, r_473__53_, r_473__52_, r_473__51_, r_473__50_, r_473__49_, r_473__48_, r_473__47_, r_473__46_, r_473__45_, r_473__44_, r_473__43_, r_473__42_, r_473__41_, r_473__40_, r_473__39_, r_473__38_, r_473__37_, r_473__36_, r_473__35_, r_473__34_, r_473__33_, r_473__32_, r_473__31_, r_473__30_, r_473__29_, r_473__28_, r_473__27_, r_473__26_, r_473__25_, r_473__24_, r_473__23_, r_473__22_, r_473__21_, r_473__20_, r_473__19_, r_473__18_, r_473__17_, r_473__16_, r_473__15_, r_473__14_, r_473__13_, r_473__12_, r_473__11_, r_473__10_, r_473__9_, r_473__8_, r_473__7_, r_473__6_, r_473__5_, r_473__4_, r_473__3_, r_473__2_, r_473__1_, r_473__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N945)? data_i : 1'b0;
  assign N944 = sel_i[944];
  assign N945 = N3388;
  assign { r_n_473__63_, r_n_473__62_, r_n_473__61_, r_n_473__60_, r_n_473__59_, r_n_473__58_, r_n_473__57_, r_n_473__56_, r_n_473__55_, r_n_473__54_, r_n_473__53_, r_n_473__52_, r_n_473__51_, r_n_473__50_, r_n_473__49_, r_n_473__48_, r_n_473__47_, r_n_473__46_, r_n_473__45_, r_n_473__44_, r_n_473__43_, r_n_473__42_, r_n_473__41_, r_n_473__40_, r_n_473__39_, r_n_473__38_, r_n_473__37_, r_n_473__36_, r_n_473__35_, r_n_473__34_, r_n_473__33_, r_n_473__32_, r_n_473__31_, r_n_473__30_, r_n_473__29_, r_n_473__28_, r_n_473__27_, r_n_473__26_, r_n_473__25_, r_n_473__24_, r_n_473__23_, r_n_473__22_, r_n_473__21_, r_n_473__20_, r_n_473__19_, r_n_473__18_, r_n_473__17_, r_n_473__16_, r_n_473__15_, r_n_473__14_, r_n_473__13_, r_n_473__12_, r_n_473__11_, r_n_473__10_, r_n_473__9_, r_n_473__8_, r_n_473__7_, r_n_473__6_, r_n_473__5_, r_n_473__4_, r_n_473__3_, r_n_473__2_, r_n_473__1_, r_n_473__0_ } = (N946)? { r_474__63_, r_474__62_, r_474__61_, r_474__60_, r_474__59_, r_474__58_, r_474__57_, r_474__56_, r_474__55_, r_474__54_, r_474__53_, r_474__52_, r_474__51_, r_474__50_, r_474__49_, r_474__48_, r_474__47_, r_474__46_, r_474__45_, r_474__44_, r_474__43_, r_474__42_, r_474__41_, r_474__40_, r_474__39_, r_474__38_, r_474__37_, r_474__36_, r_474__35_, r_474__34_, r_474__33_, r_474__32_, r_474__31_, r_474__30_, r_474__29_, r_474__28_, r_474__27_, r_474__26_, r_474__25_, r_474__24_, r_474__23_, r_474__22_, r_474__21_, r_474__20_, r_474__19_, r_474__18_, r_474__17_, r_474__16_, r_474__15_, r_474__14_, r_474__13_, r_474__12_, r_474__11_, r_474__10_, r_474__9_, r_474__8_, r_474__7_, r_474__6_, r_474__5_, r_474__4_, r_474__3_, r_474__2_, r_474__1_, r_474__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N947)? data_i : 1'b0;
  assign N946 = sel_i[946];
  assign N947 = N3393;
  assign { r_n_474__63_, r_n_474__62_, r_n_474__61_, r_n_474__60_, r_n_474__59_, r_n_474__58_, r_n_474__57_, r_n_474__56_, r_n_474__55_, r_n_474__54_, r_n_474__53_, r_n_474__52_, r_n_474__51_, r_n_474__50_, r_n_474__49_, r_n_474__48_, r_n_474__47_, r_n_474__46_, r_n_474__45_, r_n_474__44_, r_n_474__43_, r_n_474__42_, r_n_474__41_, r_n_474__40_, r_n_474__39_, r_n_474__38_, r_n_474__37_, r_n_474__36_, r_n_474__35_, r_n_474__34_, r_n_474__33_, r_n_474__32_, r_n_474__31_, r_n_474__30_, r_n_474__29_, r_n_474__28_, r_n_474__27_, r_n_474__26_, r_n_474__25_, r_n_474__24_, r_n_474__23_, r_n_474__22_, r_n_474__21_, r_n_474__20_, r_n_474__19_, r_n_474__18_, r_n_474__17_, r_n_474__16_, r_n_474__15_, r_n_474__14_, r_n_474__13_, r_n_474__12_, r_n_474__11_, r_n_474__10_, r_n_474__9_, r_n_474__8_, r_n_474__7_, r_n_474__6_, r_n_474__5_, r_n_474__4_, r_n_474__3_, r_n_474__2_, r_n_474__1_, r_n_474__0_ } = (N948)? { r_475__63_, r_475__62_, r_475__61_, r_475__60_, r_475__59_, r_475__58_, r_475__57_, r_475__56_, r_475__55_, r_475__54_, r_475__53_, r_475__52_, r_475__51_, r_475__50_, r_475__49_, r_475__48_, r_475__47_, r_475__46_, r_475__45_, r_475__44_, r_475__43_, r_475__42_, r_475__41_, r_475__40_, r_475__39_, r_475__38_, r_475__37_, r_475__36_, r_475__35_, r_475__34_, r_475__33_, r_475__32_, r_475__31_, r_475__30_, r_475__29_, r_475__28_, r_475__27_, r_475__26_, r_475__25_, r_475__24_, r_475__23_, r_475__22_, r_475__21_, r_475__20_, r_475__19_, r_475__18_, r_475__17_, r_475__16_, r_475__15_, r_475__14_, r_475__13_, r_475__12_, r_475__11_, r_475__10_, r_475__9_, r_475__8_, r_475__7_, r_475__6_, r_475__5_, r_475__4_, r_475__3_, r_475__2_, r_475__1_, r_475__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N949)? data_i : 1'b0;
  assign N948 = sel_i[948];
  assign N949 = N3398;
  assign { r_n_475__63_, r_n_475__62_, r_n_475__61_, r_n_475__60_, r_n_475__59_, r_n_475__58_, r_n_475__57_, r_n_475__56_, r_n_475__55_, r_n_475__54_, r_n_475__53_, r_n_475__52_, r_n_475__51_, r_n_475__50_, r_n_475__49_, r_n_475__48_, r_n_475__47_, r_n_475__46_, r_n_475__45_, r_n_475__44_, r_n_475__43_, r_n_475__42_, r_n_475__41_, r_n_475__40_, r_n_475__39_, r_n_475__38_, r_n_475__37_, r_n_475__36_, r_n_475__35_, r_n_475__34_, r_n_475__33_, r_n_475__32_, r_n_475__31_, r_n_475__30_, r_n_475__29_, r_n_475__28_, r_n_475__27_, r_n_475__26_, r_n_475__25_, r_n_475__24_, r_n_475__23_, r_n_475__22_, r_n_475__21_, r_n_475__20_, r_n_475__19_, r_n_475__18_, r_n_475__17_, r_n_475__16_, r_n_475__15_, r_n_475__14_, r_n_475__13_, r_n_475__12_, r_n_475__11_, r_n_475__10_, r_n_475__9_, r_n_475__8_, r_n_475__7_, r_n_475__6_, r_n_475__5_, r_n_475__4_, r_n_475__3_, r_n_475__2_, r_n_475__1_, r_n_475__0_ } = (N950)? { r_476__63_, r_476__62_, r_476__61_, r_476__60_, r_476__59_, r_476__58_, r_476__57_, r_476__56_, r_476__55_, r_476__54_, r_476__53_, r_476__52_, r_476__51_, r_476__50_, r_476__49_, r_476__48_, r_476__47_, r_476__46_, r_476__45_, r_476__44_, r_476__43_, r_476__42_, r_476__41_, r_476__40_, r_476__39_, r_476__38_, r_476__37_, r_476__36_, r_476__35_, r_476__34_, r_476__33_, r_476__32_, r_476__31_, r_476__30_, r_476__29_, r_476__28_, r_476__27_, r_476__26_, r_476__25_, r_476__24_, r_476__23_, r_476__22_, r_476__21_, r_476__20_, r_476__19_, r_476__18_, r_476__17_, r_476__16_, r_476__15_, r_476__14_, r_476__13_, r_476__12_, r_476__11_, r_476__10_, r_476__9_, r_476__8_, r_476__7_, r_476__6_, r_476__5_, r_476__4_, r_476__3_, r_476__2_, r_476__1_, r_476__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N951)? data_i : 1'b0;
  assign N950 = sel_i[950];
  assign N951 = N3403;
  assign { r_n_476__63_, r_n_476__62_, r_n_476__61_, r_n_476__60_, r_n_476__59_, r_n_476__58_, r_n_476__57_, r_n_476__56_, r_n_476__55_, r_n_476__54_, r_n_476__53_, r_n_476__52_, r_n_476__51_, r_n_476__50_, r_n_476__49_, r_n_476__48_, r_n_476__47_, r_n_476__46_, r_n_476__45_, r_n_476__44_, r_n_476__43_, r_n_476__42_, r_n_476__41_, r_n_476__40_, r_n_476__39_, r_n_476__38_, r_n_476__37_, r_n_476__36_, r_n_476__35_, r_n_476__34_, r_n_476__33_, r_n_476__32_, r_n_476__31_, r_n_476__30_, r_n_476__29_, r_n_476__28_, r_n_476__27_, r_n_476__26_, r_n_476__25_, r_n_476__24_, r_n_476__23_, r_n_476__22_, r_n_476__21_, r_n_476__20_, r_n_476__19_, r_n_476__18_, r_n_476__17_, r_n_476__16_, r_n_476__15_, r_n_476__14_, r_n_476__13_, r_n_476__12_, r_n_476__11_, r_n_476__10_, r_n_476__9_, r_n_476__8_, r_n_476__7_, r_n_476__6_, r_n_476__5_, r_n_476__4_, r_n_476__3_, r_n_476__2_, r_n_476__1_, r_n_476__0_ } = (N952)? { r_477__63_, r_477__62_, r_477__61_, r_477__60_, r_477__59_, r_477__58_, r_477__57_, r_477__56_, r_477__55_, r_477__54_, r_477__53_, r_477__52_, r_477__51_, r_477__50_, r_477__49_, r_477__48_, r_477__47_, r_477__46_, r_477__45_, r_477__44_, r_477__43_, r_477__42_, r_477__41_, r_477__40_, r_477__39_, r_477__38_, r_477__37_, r_477__36_, r_477__35_, r_477__34_, r_477__33_, r_477__32_, r_477__31_, r_477__30_, r_477__29_, r_477__28_, r_477__27_, r_477__26_, r_477__25_, r_477__24_, r_477__23_, r_477__22_, r_477__21_, r_477__20_, r_477__19_, r_477__18_, r_477__17_, r_477__16_, r_477__15_, r_477__14_, r_477__13_, r_477__12_, r_477__11_, r_477__10_, r_477__9_, r_477__8_, r_477__7_, r_477__6_, r_477__5_, r_477__4_, r_477__3_, r_477__2_, r_477__1_, r_477__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N953)? data_i : 1'b0;
  assign N952 = sel_i[952];
  assign N953 = N3408;
  assign { r_n_477__63_, r_n_477__62_, r_n_477__61_, r_n_477__60_, r_n_477__59_, r_n_477__58_, r_n_477__57_, r_n_477__56_, r_n_477__55_, r_n_477__54_, r_n_477__53_, r_n_477__52_, r_n_477__51_, r_n_477__50_, r_n_477__49_, r_n_477__48_, r_n_477__47_, r_n_477__46_, r_n_477__45_, r_n_477__44_, r_n_477__43_, r_n_477__42_, r_n_477__41_, r_n_477__40_, r_n_477__39_, r_n_477__38_, r_n_477__37_, r_n_477__36_, r_n_477__35_, r_n_477__34_, r_n_477__33_, r_n_477__32_, r_n_477__31_, r_n_477__30_, r_n_477__29_, r_n_477__28_, r_n_477__27_, r_n_477__26_, r_n_477__25_, r_n_477__24_, r_n_477__23_, r_n_477__22_, r_n_477__21_, r_n_477__20_, r_n_477__19_, r_n_477__18_, r_n_477__17_, r_n_477__16_, r_n_477__15_, r_n_477__14_, r_n_477__13_, r_n_477__12_, r_n_477__11_, r_n_477__10_, r_n_477__9_, r_n_477__8_, r_n_477__7_, r_n_477__6_, r_n_477__5_, r_n_477__4_, r_n_477__3_, r_n_477__2_, r_n_477__1_, r_n_477__0_ } = (N954)? { r_478__63_, r_478__62_, r_478__61_, r_478__60_, r_478__59_, r_478__58_, r_478__57_, r_478__56_, r_478__55_, r_478__54_, r_478__53_, r_478__52_, r_478__51_, r_478__50_, r_478__49_, r_478__48_, r_478__47_, r_478__46_, r_478__45_, r_478__44_, r_478__43_, r_478__42_, r_478__41_, r_478__40_, r_478__39_, r_478__38_, r_478__37_, r_478__36_, r_478__35_, r_478__34_, r_478__33_, r_478__32_, r_478__31_, r_478__30_, r_478__29_, r_478__28_, r_478__27_, r_478__26_, r_478__25_, r_478__24_, r_478__23_, r_478__22_, r_478__21_, r_478__20_, r_478__19_, r_478__18_, r_478__17_, r_478__16_, r_478__15_, r_478__14_, r_478__13_, r_478__12_, r_478__11_, r_478__10_, r_478__9_, r_478__8_, r_478__7_, r_478__6_, r_478__5_, r_478__4_, r_478__3_, r_478__2_, r_478__1_, r_478__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N955)? data_i : 1'b0;
  assign N954 = sel_i[954];
  assign N955 = N3413;
  assign { r_n_478__63_, r_n_478__62_, r_n_478__61_, r_n_478__60_, r_n_478__59_, r_n_478__58_, r_n_478__57_, r_n_478__56_, r_n_478__55_, r_n_478__54_, r_n_478__53_, r_n_478__52_, r_n_478__51_, r_n_478__50_, r_n_478__49_, r_n_478__48_, r_n_478__47_, r_n_478__46_, r_n_478__45_, r_n_478__44_, r_n_478__43_, r_n_478__42_, r_n_478__41_, r_n_478__40_, r_n_478__39_, r_n_478__38_, r_n_478__37_, r_n_478__36_, r_n_478__35_, r_n_478__34_, r_n_478__33_, r_n_478__32_, r_n_478__31_, r_n_478__30_, r_n_478__29_, r_n_478__28_, r_n_478__27_, r_n_478__26_, r_n_478__25_, r_n_478__24_, r_n_478__23_, r_n_478__22_, r_n_478__21_, r_n_478__20_, r_n_478__19_, r_n_478__18_, r_n_478__17_, r_n_478__16_, r_n_478__15_, r_n_478__14_, r_n_478__13_, r_n_478__12_, r_n_478__11_, r_n_478__10_, r_n_478__9_, r_n_478__8_, r_n_478__7_, r_n_478__6_, r_n_478__5_, r_n_478__4_, r_n_478__3_, r_n_478__2_, r_n_478__1_, r_n_478__0_ } = (N956)? { r_479__63_, r_479__62_, r_479__61_, r_479__60_, r_479__59_, r_479__58_, r_479__57_, r_479__56_, r_479__55_, r_479__54_, r_479__53_, r_479__52_, r_479__51_, r_479__50_, r_479__49_, r_479__48_, r_479__47_, r_479__46_, r_479__45_, r_479__44_, r_479__43_, r_479__42_, r_479__41_, r_479__40_, r_479__39_, r_479__38_, r_479__37_, r_479__36_, r_479__35_, r_479__34_, r_479__33_, r_479__32_, r_479__31_, r_479__30_, r_479__29_, r_479__28_, r_479__27_, r_479__26_, r_479__25_, r_479__24_, r_479__23_, r_479__22_, r_479__21_, r_479__20_, r_479__19_, r_479__18_, r_479__17_, r_479__16_, r_479__15_, r_479__14_, r_479__13_, r_479__12_, r_479__11_, r_479__10_, r_479__9_, r_479__8_, r_479__7_, r_479__6_, r_479__5_, r_479__4_, r_479__3_, r_479__2_, r_479__1_, r_479__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N957)? data_i : 1'b0;
  assign N956 = sel_i[956];
  assign N957 = N3418;
  assign { r_n_479__63_, r_n_479__62_, r_n_479__61_, r_n_479__60_, r_n_479__59_, r_n_479__58_, r_n_479__57_, r_n_479__56_, r_n_479__55_, r_n_479__54_, r_n_479__53_, r_n_479__52_, r_n_479__51_, r_n_479__50_, r_n_479__49_, r_n_479__48_, r_n_479__47_, r_n_479__46_, r_n_479__45_, r_n_479__44_, r_n_479__43_, r_n_479__42_, r_n_479__41_, r_n_479__40_, r_n_479__39_, r_n_479__38_, r_n_479__37_, r_n_479__36_, r_n_479__35_, r_n_479__34_, r_n_479__33_, r_n_479__32_, r_n_479__31_, r_n_479__30_, r_n_479__29_, r_n_479__28_, r_n_479__27_, r_n_479__26_, r_n_479__25_, r_n_479__24_, r_n_479__23_, r_n_479__22_, r_n_479__21_, r_n_479__20_, r_n_479__19_, r_n_479__18_, r_n_479__17_, r_n_479__16_, r_n_479__15_, r_n_479__14_, r_n_479__13_, r_n_479__12_, r_n_479__11_, r_n_479__10_, r_n_479__9_, r_n_479__8_, r_n_479__7_, r_n_479__6_, r_n_479__5_, r_n_479__4_, r_n_479__3_, r_n_479__2_, r_n_479__1_, r_n_479__0_ } = (N958)? { r_480__63_, r_480__62_, r_480__61_, r_480__60_, r_480__59_, r_480__58_, r_480__57_, r_480__56_, r_480__55_, r_480__54_, r_480__53_, r_480__52_, r_480__51_, r_480__50_, r_480__49_, r_480__48_, r_480__47_, r_480__46_, r_480__45_, r_480__44_, r_480__43_, r_480__42_, r_480__41_, r_480__40_, r_480__39_, r_480__38_, r_480__37_, r_480__36_, r_480__35_, r_480__34_, r_480__33_, r_480__32_, r_480__31_, r_480__30_, r_480__29_, r_480__28_, r_480__27_, r_480__26_, r_480__25_, r_480__24_, r_480__23_, r_480__22_, r_480__21_, r_480__20_, r_480__19_, r_480__18_, r_480__17_, r_480__16_, r_480__15_, r_480__14_, r_480__13_, r_480__12_, r_480__11_, r_480__10_, r_480__9_, r_480__8_, r_480__7_, r_480__6_, r_480__5_, r_480__4_, r_480__3_, r_480__2_, r_480__1_, r_480__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N959)? data_i : 1'b0;
  assign N958 = sel_i[958];
  assign N959 = N3423;
  assign { r_n_480__63_, r_n_480__62_, r_n_480__61_, r_n_480__60_, r_n_480__59_, r_n_480__58_, r_n_480__57_, r_n_480__56_, r_n_480__55_, r_n_480__54_, r_n_480__53_, r_n_480__52_, r_n_480__51_, r_n_480__50_, r_n_480__49_, r_n_480__48_, r_n_480__47_, r_n_480__46_, r_n_480__45_, r_n_480__44_, r_n_480__43_, r_n_480__42_, r_n_480__41_, r_n_480__40_, r_n_480__39_, r_n_480__38_, r_n_480__37_, r_n_480__36_, r_n_480__35_, r_n_480__34_, r_n_480__33_, r_n_480__32_, r_n_480__31_, r_n_480__30_, r_n_480__29_, r_n_480__28_, r_n_480__27_, r_n_480__26_, r_n_480__25_, r_n_480__24_, r_n_480__23_, r_n_480__22_, r_n_480__21_, r_n_480__20_, r_n_480__19_, r_n_480__18_, r_n_480__17_, r_n_480__16_, r_n_480__15_, r_n_480__14_, r_n_480__13_, r_n_480__12_, r_n_480__11_, r_n_480__10_, r_n_480__9_, r_n_480__8_, r_n_480__7_, r_n_480__6_, r_n_480__5_, r_n_480__4_, r_n_480__3_, r_n_480__2_, r_n_480__1_, r_n_480__0_ } = (N960)? { r_481__63_, r_481__62_, r_481__61_, r_481__60_, r_481__59_, r_481__58_, r_481__57_, r_481__56_, r_481__55_, r_481__54_, r_481__53_, r_481__52_, r_481__51_, r_481__50_, r_481__49_, r_481__48_, r_481__47_, r_481__46_, r_481__45_, r_481__44_, r_481__43_, r_481__42_, r_481__41_, r_481__40_, r_481__39_, r_481__38_, r_481__37_, r_481__36_, r_481__35_, r_481__34_, r_481__33_, r_481__32_, r_481__31_, r_481__30_, r_481__29_, r_481__28_, r_481__27_, r_481__26_, r_481__25_, r_481__24_, r_481__23_, r_481__22_, r_481__21_, r_481__20_, r_481__19_, r_481__18_, r_481__17_, r_481__16_, r_481__15_, r_481__14_, r_481__13_, r_481__12_, r_481__11_, r_481__10_, r_481__9_, r_481__8_, r_481__7_, r_481__6_, r_481__5_, r_481__4_, r_481__3_, r_481__2_, r_481__1_, r_481__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N961)? data_i : 1'b0;
  assign N960 = sel_i[960];
  assign N961 = N3428;
  assign { r_n_481__63_, r_n_481__62_, r_n_481__61_, r_n_481__60_, r_n_481__59_, r_n_481__58_, r_n_481__57_, r_n_481__56_, r_n_481__55_, r_n_481__54_, r_n_481__53_, r_n_481__52_, r_n_481__51_, r_n_481__50_, r_n_481__49_, r_n_481__48_, r_n_481__47_, r_n_481__46_, r_n_481__45_, r_n_481__44_, r_n_481__43_, r_n_481__42_, r_n_481__41_, r_n_481__40_, r_n_481__39_, r_n_481__38_, r_n_481__37_, r_n_481__36_, r_n_481__35_, r_n_481__34_, r_n_481__33_, r_n_481__32_, r_n_481__31_, r_n_481__30_, r_n_481__29_, r_n_481__28_, r_n_481__27_, r_n_481__26_, r_n_481__25_, r_n_481__24_, r_n_481__23_, r_n_481__22_, r_n_481__21_, r_n_481__20_, r_n_481__19_, r_n_481__18_, r_n_481__17_, r_n_481__16_, r_n_481__15_, r_n_481__14_, r_n_481__13_, r_n_481__12_, r_n_481__11_, r_n_481__10_, r_n_481__9_, r_n_481__8_, r_n_481__7_, r_n_481__6_, r_n_481__5_, r_n_481__4_, r_n_481__3_, r_n_481__2_, r_n_481__1_, r_n_481__0_ } = (N962)? { r_482__63_, r_482__62_, r_482__61_, r_482__60_, r_482__59_, r_482__58_, r_482__57_, r_482__56_, r_482__55_, r_482__54_, r_482__53_, r_482__52_, r_482__51_, r_482__50_, r_482__49_, r_482__48_, r_482__47_, r_482__46_, r_482__45_, r_482__44_, r_482__43_, r_482__42_, r_482__41_, r_482__40_, r_482__39_, r_482__38_, r_482__37_, r_482__36_, r_482__35_, r_482__34_, r_482__33_, r_482__32_, r_482__31_, r_482__30_, r_482__29_, r_482__28_, r_482__27_, r_482__26_, r_482__25_, r_482__24_, r_482__23_, r_482__22_, r_482__21_, r_482__20_, r_482__19_, r_482__18_, r_482__17_, r_482__16_, r_482__15_, r_482__14_, r_482__13_, r_482__12_, r_482__11_, r_482__10_, r_482__9_, r_482__8_, r_482__7_, r_482__6_, r_482__5_, r_482__4_, r_482__3_, r_482__2_, r_482__1_, r_482__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N963)? data_i : 1'b0;
  assign N962 = sel_i[962];
  assign N963 = N3433;
  assign { r_n_482__63_, r_n_482__62_, r_n_482__61_, r_n_482__60_, r_n_482__59_, r_n_482__58_, r_n_482__57_, r_n_482__56_, r_n_482__55_, r_n_482__54_, r_n_482__53_, r_n_482__52_, r_n_482__51_, r_n_482__50_, r_n_482__49_, r_n_482__48_, r_n_482__47_, r_n_482__46_, r_n_482__45_, r_n_482__44_, r_n_482__43_, r_n_482__42_, r_n_482__41_, r_n_482__40_, r_n_482__39_, r_n_482__38_, r_n_482__37_, r_n_482__36_, r_n_482__35_, r_n_482__34_, r_n_482__33_, r_n_482__32_, r_n_482__31_, r_n_482__30_, r_n_482__29_, r_n_482__28_, r_n_482__27_, r_n_482__26_, r_n_482__25_, r_n_482__24_, r_n_482__23_, r_n_482__22_, r_n_482__21_, r_n_482__20_, r_n_482__19_, r_n_482__18_, r_n_482__17_, r_n_482__16_, r_n_482__15_, r_n_482__14_, r_n_482__13_, r_n_482__12_, r_n_482__11_, r_n_482__10_, r_n_482__9_, r_n_482__8_, r_n_482__7_, r_n_482__6_, r_n_482__5_, r_n_482__4_, r_n_482__3_, r_n_482__2_, r_n_482__1_, r_n_482__0_ } = (N964)? { r_483__63_, r_483__62_, r_483__61_, r_483__60_, r_483__59_, r_483__58_, r_483__57_, r_483__56_, r_483__55_, r_483__54_, r_483__53_, r_483__52_, r_483__51_, r_483__50_, r_483__49_, r_483__48_, r_483__47_, r_483__46_, r_483__45_, r_483__44_, r_483__43_, r_483__42_, r_483__41_, r_483__40_, r_483__39_, r_483__38_, r_483__37_, r_483__36_, r_483__35_, r_483__34_, r_483__33_, r_483__32_, r_483__31_, r_483__30_, r_483__29_, r_483__28_, r_483__27_, r_483__26_, r_483__25_, r_483__24_, r_483__23_, r_483__22_, r_483__21_, r_483__20_, r_483__19_, r_483__18_, r_483__17_, r_483__16_, r_483__15_, r_483__14_, r_483__13_, r_483__12_, r_483__11_, r_483__10_, r_483__9_, r_483__8_, r_483__7_, r_483__6_, r_483__5_, r_483__4_, r_483__3_, r_483__2_, r_483__1_, r_483__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N965)? data_i : 1'b0;
  assign N964 = sel_i[964];
  assign N965 = N3438;
  assign { r_n_483__63_, r_n_483__62_, r_n_483__61_, r_n_483__60_, r_n_483__59_, r_n_483__58_, r_n_483__57_, r_n_483__56_, r_n_483__55_, r_n_483__54_, r_n_483__53_, r_n_483__52_, r_n_483__51_, r_n_483__50_, r_n_483__49_, r_n_483__48_, r_n_483__47_, r_n_483__46_, r_n_483__45_, r_n_483__44_, r_n_483__43_, r_n_483__42_, r_n_483__41_, r_n_483__40_, r_n_483__39_, r_n_483__38_, r_n_483__37_, r_n_483__36_, r_n_483__35_, r_n_483__34_, r_n_483__33_, r_n_483__32_, r_n_483__31_, r_n_483__30_, r_n_483__29_, r_n_483__28_, r_n_483__27_, r_n_483__26_, r_n_483__25_, r_n_483__24_, r_n_483__23_, r_n_483__22_, r_n_483__21_, r_n_483__20_, r_n_483__19_, r_n_483__18_, r_n_483__17_, r_n_483__16_, r_n_483__15_, r_n_483__14_, r_n_483__13_, r_n_483__12_, r_n_483__11_, r_n_483__10_, r_n_483__9_, r_n_483__8_, r_n_483__7_, r_n_483__6_, r_n_483__5_, r_n_483__4_, r_n_483__3_, r_n_483__2_, r_n_483__1_, r_n_483__0_ } = (N966)? { r_484__63_, r_484__62_, r_484__61_, r_484__60_, r_484__59_, r_484__58_, r_484__57_, r_484__56_, r_484__55_, r_484__54_, r_484__53_, r_484__52_, r_484__51_, r_484__50_, r_484__49_, r_484__48_, r_484__47_, r_484__46_, r_484__45_, r_484__44_, r_484__43_, r_484__42_, r_484__41_, r_484__40_, r_484__39_, r_484__38_, r_484__37_, r_484__36_, r_484__35_, r_484__34_, r_484__33_, r_484__32_, r_484__31_, r_484__30_, r_484__29_, r_484__28_, r_484__27_, r_484__26_, r_484__25_, r_484__24_, r_484__23_, r_484__22_, r_484__21_, r_484__20_, r_484__19_, r_484__18_, r_484__17_, r_484__16_, r_484__15_, r_484__14_, r_484__13_, r_484__12_, r_484__11_, r_484__10_, r_484__9_, r_484__8_, r_484__7_, r_484__6_, r_484__5_, r_484__4_, r_484__3_, r_484__2_, r_484__1_, r_484__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N967)? data_i : 1'b0;
  assign N966 = sel_i[966];
  assign N967 = N3443;
  assign { r_n_484__63_, r_n_484__62_, r_n_484__61_, r_n_484__60_, r_n_484__59_, r_n_484__58_, r_n_484__57_, r_n_484__56_, r_n_484__55_, r_n_484__54_, r_n_484__53_, r_n_484__52_, r_n_484__51_, r_n_484__50_, r_n_484__49_, r_n_484__48_, r_n_484__47_, r_n_484__46_, r_n_484__45_, r_n_484__44_, r_n_484__43_, r_n_484__42_, r_n_484__41_, r_n_484__40_, r_n_484__39_, r_n_484__38_, r_n_484__37_, r_n_484__36_, r_n_484__35_, r_n_484__34_, r_n_484__33_, r_n_484__32_, r_n_484__31_, r_n_484__30_, r_n_484__29_, r_n_484__28_, r_n_484__27_, r_n_484__26_, r_n_484__25_, r_n_484__24_, r_n_484__23_, r_n_484__22_, r_n_484__21_, r_n_484__20_, r_n_484__19_, r_n_484__18_, r_n_484__17_, r_n_484__16_, r_n_484__15_, r_n_484__14_, r_n_484__13_, r_n_484__12_, r_n_484__11_, r_n_484__10_, r_n_484__9_, r_n_484__8_, r_n_484__7_, r_n_484__6_, r_n_484__5_, r_n_484__4_, r_n_484__3_, r_n_484__2_, r_n_484__1_, r_n_484__0_ } = (N968)? { r_485__63_, r_485__62_, r_485__61_, r_485__60_, r_485__59_, r_485__58_, r_485__57_, r_485__56_, r_485__55_, r_485__54_, r_485__53_, r_485__52_, r_485__51_, r_485__50_, r_485__49_, r_485__48_, r_485__47_, r_485__46_, r_485__45_, r_485__44_, r_485__43_, r_485__42_, r_485__41_, r_485__40_, r_485__39_, r_485__38_, r_485__37_, r_485__36_, r_485__35_, r_485__34_, r_485__33_, r_485__32_, r_485__31_, r_485__30_, r_485__29_, r_485__28_, r_485__27_, r_485__26_, r_485__25_, r_485__24_, r_485__23_, r_485__22_, r_485__21_, r_485__20_, r_485__19_, r_485__18_, r_485__17_, r_485__16_, r_485__15_, r_485__14_, r_485__13_, r_485__12_, r_485__11_, r_485__10_, r_485__9_, r_485__8_, r_485__7_, r_485__6_, r_485__5_, r_485__4_, r_485__3_, r_485__2_, r_485__1_, r_485__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N969)? data_i : 1'b0;
  assign N968 = sel_i[968];
  assign N969 = N3448;
  assign { r_n_485__63_, r_n_485__62_, r_n_485__61_, r_n_485__60_, r_n_485__59_, r_n_485__58_, r_n_485__57_, r_n_485__56_, r_n_485__55_, r_n_485__54_, r_n_485__53_, r_n_485__52_, r_n_485__51_, r_n_485__50_, r_n_485__49_, r_n_485__48_, r_n_485__47_, r_n_485__46_, r_n_485__45_, r_n_485__44_, r_n_485__43_, r_n_485__42_, r_n_485__41_, r_n_485__40_, r_n_485__39_, r_n_485__38_, r_n_485__37_, r_n_485__36_, r_n_485__35_, r_n_485__34_, r_n_485__33_, r_n_485__32_, r_n_485__31_, r_n_485__30_, r_n_485__29_, r_n_485__28_, r_n_485__27_, r_n_485__26_, r_n_485__25_, r_n_485__24_, r_n_485__23_, r_n_485__22_, r_n_485__21_, r_n_485__20_, r_n_485__19_, r_n_485__18_, r_n_485__17_, r_n_485__16_, r_n_485__15_, r_n_485__14_, r_n_485__13_, r_n_485__12_, r_n_485__11_, r_n_485__10_, r_n_485__9_, r_n_485__8_, r_n_485__7_, r_n_485__6_, r_n_485__5_, r_n_485__4_, r_n_485__3_, r_n_485__2_, r_n_485__1_, r_n_485__0_ } = (N970)? { r_486__63_, r_486__62_, r_486__61_, r_486__60_, r_486__59_, r_486__58_, r_486__57_, r_486__56_, r_486__55_, r_486__54_, r_486__53_, r_486__52_, r_486__51_, r_486__50_, r_486__49_, r_486__48_, r_486__47_, r_486__46_, r_486__45_, r_486__44_, r_486__43_, r_486__42_, r_486__41_, r_486__40_, r_486__39_, r_486__38_, r_486__37_, r_486__36_, r_486__35_, r_486__34_, r_486__33_, r_486__32_, r_486__31_, r_486__30_, r_486__29_, r_486__28_, r_486__27_, r_486__26_, r_486__25_, r_486__24_, r_486__23_, r_486__22_, r_486__21_, r_486__20_, r_486__19_, r_486__18_, r_486__17_, r_486__16_, r_486__15_, r_486__14_, r_486__13_, r_486__12_, r_486__11_, r_486__10_, r_486__9_, r_486__8_, r_486__7_, r_486__6_, r_486__5_, r_486__4_, r_486__3_, r_486__2_, r_486__1_, r_486__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N971)? data_i : 1'b0;
  assign N970 = sel_i[970];
  assign N971 = N3453;
  assign { r_n_486__63_, r_n_486__62_, r_n_486__61_, r_n_486__60_, r_n_486__59_, r_n_486__58_, r_n_486__57_, r_n_486__56_, r_n_486__55_, r_n_486__54_, r_n_486__53_, r_n_486__52_, r_n_486__51_, r_n_486__50_, r_n_486__49_, r_n_486__48_, r_n_486__47_, r_n_486__46_, r_n_486__45_, r_n_486__44_, r_n_486__43_, r_n_486__42_, r_n_486__41_, r_n_486__40_, r_n_486__39_, r_n_486__38_, r_n_486__37_, r_n_486__36_, r_n_486__35_, r_n_486__34_, r_n_486__33_, r_n_486__32_, r_n_486__31_, r_n_486__30_, r_n_486__29_, r_n_486__28_, r_n_486__27_, r_n_486__26_, r_n_486__25_, r_n_486__24_, r_n_486__23_, r_n_486__22_, r_n_486__21_, r_n_486__20_, r_n_486__19_, r_n_486__18_, r_n_486__17_, r_n_486__16_, r_n_486__15_, r_n_486__14_, r_n_486__13_, r_n_486__12_, r_n_486__11_, r_n_486__10_, r_n_486__9_, r_n_486__8_, r_n_486__7_, r_n_486__6_, r_n_486__5_, r_n_486__4_, r_n_486__3_, r_n_486__2_, r_n_486__1_, r_n_486__0_ } = (N972)? { r_487__63_, r_487__62_, r_487__61_, r_487__60_, r_487__59_, r_487__58_, r_487__57_, r_487__56_, r_487__55_, r_487__54_, r_487__53_, r_487__52_, r_487__51_, r_487__50_, r_487__49_, r_487__48_, r_487__47_, r_487__46_, r_487__45_, r_487__44_, r_487__43_, r_487__42_, r_487__41_, r_487__40_, r_487__39_, r_487__38_, r_487__37_, r_487__36_, r_487__35_, r_487__34_, r_487__33_, r_487__32_, r_487__31_, r_487__30_, r_487__29_, r_487__28_, r_487__27_, r_487__26_, r_487__25_, r_487__24_, r_487__23_, r_487__22_, r_487__21_, r_487__20_, r_487__19_, r_487__18_, r_487__17_, r_487__16_, r_487__15_, r_487__14_, r_487__13_, r_487__12_, r_487__11_, r_487__10_, r_487__9_, r_487__8_, r_487__7_, r_487__6_, r_487__5_, r_487__4_, r_487__3_, r_487__2_, r_487__1_, r_487__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N973)? data_i : 1'b0;
  assign N972 = sel_i[972];
  assign N973 = N3458;
  assign { r_n_487__63_, r_n_487__62_, r_n_487__61_, r_n_487__60_, r_n_487__59_, r_n_487__58_, r_n_487__57_, r_n_487__56_, r_n_487__55_, r_n_487__54_, r_n_487__53_, r_n_487__52_, r_n_487__51_, r_n_487__50_, r_n_487__49_, r_n_487__48_, r_n_487__47_, r_n_487__46_, r_n_487__45_, r_n_487__44_, r_n_487__43_, r_n_487__42_, r_n_487__41_, r_n_487__40_, r_n_487__39_, r_n_487__38_, r_n_487__37_, r_n_487__36_, r_n_487__35_, r_n_487__34_, r_n_487__33_, r_n_487__32_, r_n_487__31_, r_n_487__30_, r_n_487__29_, r_n_487__28_, r_n_487__27_, r_n_487__26_, r_n_487__25_, r_n_487__24_, r_n_487__23_, r_n_487__22_, r_n_487__21_, r_n_487__20_, r_n_487__19_, r_n_487__18_, r_n_487__17_, r_n_487__16_, r_n_487__15_, r_n_487__14_, r_n_487__13_, r_n_487__12_, r_n_487__11_, r_n_487__10_, r_n_487__9_, r_n_487__8_, r_n_487__7_, r_n_487__6_, r_n_487__5_, r_n_487__4_, r_n_487__3_, r_n_487__2_, r_n_487__1_, r_n_487__0_ } = (N974)? { r_488__63_, r_488__62_, r_488__61_, r_488__60_, r_488__59_, r_488__58_, r_488__57_, r_488__56_, r_488__55_, r_488__54_, r_488__53_, r_488__52_, r_488__51_, r_488__50_, r_488__49_, r_488__48_, r_488__47_, r_488__46_, r_488__45_, r_488__44_, r_488__43_, r_488__42_, r_488__41_, r_488__40_, r_488__39_, r_488__38_, r_488__37_, r_488__36_, r_488__35_, r_488__34_, r_488__33_, r_488__32_, r_488__31_, r_488__30_, r_488__29_, r_488__28_, r_488__27_, r_488__26_, r_488__25_, r_488__24_, r_488__23_, r_488__22_, r_488__21_, r_488__20_, r_488__19_, r_488__18_, r_488__17_, r_488__16_, r_488__15_, r_488__14_, r_488__13_, r_488__12_, r_488__11_, r_488__10_, r_488__9_, r_488__8_, r_488__7_, r_488__6_, r_488__5_, r_488__4_, r_488__3_, r_488__2_, r_488__1_, r_488__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N975)? data_i : 1'b0;
  assign N974 = sel_i[974];
  assign N975 = N3463;
  assign { r_n_488__63_, r_n_488__62_, r_n_488__61_, r_n_488__60_, r_n_488__59_, r_n_488__58_, r_n_488__57_, r_n_488__56_, r_n_488__55_, r_n_488__54_, r_n_488__53_, r_n_488__52_, r_n_488__51_, r_n_488__50_, r_n_488__49_, r_n_488__48_, r_n_488__47_, r_n_488__46_, r_n_488__45_, r_n_488__44_, r_n_488__43_, r_n_488__42_, r_n_488__41_, r_n_488__40_, r_n_488__39_, r_n_488__38_, r_n_488__37_, r_n_488__36_, r_n_488__35_, r_n_488__34_, r_n_488__33_, r_n_488__32_, r_n_488__31_, r_n_488__30_, r_n_488__29_, r_n_488__28_, r_n_488__27_, r_n_488__26_, r_n_488__25_, r_n_488__24_, r_n_488__23_, r_n_488__22_, r_n_488__21_, r_n_488__20_, r_n_488__19_, r_n_488__18_, r_n_488__17_, r_n_488__16_, r_n_488__15_, r_n_488__14_, r_n_488__13_, r_n_488__12_, r_n_488__11_, r_n_488__10_, r_n_488__9_, r_n_488__8_, r_n_488__7_, r_n_488__6_, r_n_488__5_, r_n_488__4_, r_n_488__3_, r_n_488__2_, r_n_488__1_, r_n_488__0_ } = (N976)? { r_489__63_, r_489__62_, r_489__61_, r_489__60_, r_489__59_, r_489__58_, r_489__57_, r_489__56_, r_489__55_, r_489__54_, r_489__53_, r_489__52_, r_489__51_, r_489__50_, r_489__49_, r_489__48_, r_489__47_, r_489__46_, r_489__45_, r_489__44_, r_489__43_, r_489__42_, r_489__41_, r_489__40_, r_489__39_, r_489__38_, r_489__37_, r_489__36_, r_489__35_, r_489__34_, r_489__33_, r_489__32_, r_489__31_, r_489__30_, r_489__29_, r_489__28_, r_489__27_, r_489__26_, r_489__25_, r_489__24_, r_489__23_, r_489__22_, r_489__21_, r_489__20_, r_489__19_, r_489__18_, r_489__17_, r_489__16_, r_489__15_, r_489__14_, r_489__13_, r_489__12_, r_489__11_, r_489__10_, r_489__9_, r_489__8_, r_489__7_, r_489__6_, r_489__5_, r_489__4_, r_489__3_, r_489__2_, r_489__1_, r_489__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N977)? data_i : 1'b0;
  assign N976 = sel_i[976];
  assign N977 = N3468;
  assign { r_n_489__63_, r_n_489__62_, r_n_489__61_, r_n_489__60_, r_n_489__59_, r_n_489__58_, r_n_489__57_, r_n_489__56_, r_n_489__55_, r_n_489__54_, r_n_489__53_, r_n_489__52_, r_n_489__51_, r_n_489__50_, r_n_489__49_, r_n_489__48_, r_n_489__47_, r_n_489__46_, r_n_489__45_, r_n_489__44_, r_n_489__43_, r_n_489__42_, r_n_489__41_, r_n_489__40_, r_n_489__39_, r_n_489__38_, r_n_489__37_, r_n_489__36_, r_n_489__35_, r_n_489__34_, r_n_489__33_, r_n_489__32_, r_n_489__31_, r_n_489__30_, r_n_489__29_, r_n_489__28_, r_n_489__27_, r_n_489__26_, r_n_489__25_, r_n_489__24_, r_n_489__23_, r_n_489__22_, r_n_489__21_, r_n_489__20_, r_n_489__19_, r_n_489__18_, r_n_489__17_, r_n_489__16_, r_n_489__15_, r_n_489__14_, r_n_489__13_, r_n_489__12_, r_n_489__11_, r_n_489__10_, r_n_489__9_, r_n_489__8_, r_n_489__7_, r_n_489__6_, r_n_489__5_, r_n_489__4_, r_n_489__3_, r_n_489__2_, r_n_489__1_, r_n_489__0_ } = (N978)? { r_490__63_, r_490__62_, r_490__61_, r_490__60_, r_490__59_, r_490__58_, r_490__57_, r_490__56_, r_490__55_, r_490__54_, r_490__53_, r_490__52_, r_490__51_, r_490__50_, r_490__49_, r_490__48_, r_490__47_, r_490__46_, r_490__45_, r_490__44_, r_490__43_, r_490__42_, r_490__41_, r_490__40_, r_490__39_, r_490__38_, r_490__37_, r_490__36_, r_490__35_, r_490__34_, r_490__33_, r_490__32_, r_490__31_, r_490__30_, r_490__29_, r_490__28_, r_490__27_, r_490__26_, r_490__25_, r_490__24_, r_490__23_, r_490__22_, r_490__21_, r_490__20_, r_490__19_, r_490__18_, r_490__17_, r_490__16_, r_490__15_, r_490__14_, r_490__13_, r_490__12_, r_490__11_, r_490__10_, r_490__9_, r_490__8_, r_490__7_, r_490__6_, r_490__5_, r_490__4_, r_490__3_, r_490__2_, r_490__1_, r_490__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N979)? data_i : 1'b0;
  assign N978 = sel_i[978];
  assign N979 = N3473;
  assign { r_n_490__63_, r_n_490__62_, r_n_490__61_, r_n_490__60_, r_n_490__59_, r_n_490__58_, r_n_490__57_, r_n_490__56_, r_n_490__55_, r_n_490__54_, r_n_490__53_, r_n_490__52_, r_n_490__51_, r_n_490__50_, r_n_490__49_, r_n_490__48_, r_n_490__47_, r_n_490__46_, r_n_490__45_, r_n_490__44_, r_n_490__43_, r_n_490__42_, r_n_490__41_, r_n_490__40_, r_n_490__39_, r_n_490__38_, r_n_490__37_, r_n_490__36_, r_n_490__35_, r_n_490__34_, r_n_490__33_, r_n_490__32_, r_n_490__31_, r_n_490__30_, r_n_490__29_, r_n_490__28_, r_n_490__27_, r_n_490__26_, r_n_490__25_, r_n_490__24_, r_n_490__23_, r_n_490__22_, r_n_490__21_, r_n_490__20_, r_n_490__19_, r_n_490__18_, r_n_490__17_, r_n_490__16_, r_n_490__15_, r_n_490__14_, r_n_490__13_, r_n_490__12_, r_n_490__11_, r_n_490__10_, r_n_490__9_, r_n_490__8_, r_n_490__7_, r_n_490__6_, r_n_490__5_, r_n_490__4_, r_n_490__3_, r_n_490__2_, r_n_490__1_, r_n_490__0_ } = (N980)? { r_491__63_, r_491__62_, r_491__61_, r_491__60_, r_491__59_, r_491__58_, r_491__57_, r_491__56_, r_491__55_, r_491__54_, r_491__53_, r_491__52_, r_491__51_, r_491__50_, r_491__49_, r_491__48_, r_491__47_, r_491__46_, r_491__45_, r_491__44_, r_491__43_, r_491__42_, r_491__41_, r_491__40_, r_491__39_, r_491__38_, r_491__37_, r_491__36_, r_491__35_, r_491__34_, r_491__33_, r_491__32_, r_491__31_, r_491__30_, r_491__29_, r_491__28_, r_491__27_, r_491__26_, r_491__25_, r_491__24_, r_491__23_, r_491__22_, r_491__21_, r_491__20_, r_491__19_, r_491__18_, r_491__17_, r_491__16_, r_491__15_, r_491__14_, r_491__13_, r_491__12_, r_491__11_, r_491__10_, r_491__9_, r_491__8_, r_491__7_, r_491__6_, r_491__5_, r_491__4_, r_491__3_, r_491__2_, r_491__1_, r_491__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N981)? data_i : 1'b0;
  assign N980 = sel_i[980];
  assign N981 = N3478;
  assign { r_n_491__63_, r_n_491__62_, r_n_491__61_, r_n_491__60_, r_n_491__59_, r_n_491__58_, r_n_491__57_, r_n_491__56_, r_n_491__55_, r_n_491__54_, r_n_491__53_, r_n_491__52_, r_n_491__51_, r_n_491__50_, r_n_491__49_, r_n_491__48_, r_n_491__47_, r_n_491__46_, r_n_491__45_, r_n_491__44_, r_n_491__43_, r_n_491__42_, r_n_491__41_, r_n_491__40_, r_n_491__39_, r_n_491__38_, r_n_491__37_, r_n_491__36_, r_n_491__35_, r_n_491__34_, r_n_491__33_, r_n_491__32_, r_n_491__31_, r_n_491__30_, r_n_491__29_, r_n_491__28_, r_n_491__27_, r_n_491__26_, r_n_491__25_, r_n_491__24_, r_n_491__23_, r_n_491__22_, r_n_491__21_, r_n_491__20_, r_n_491__19_, r_n_491__18_, r_n_491__17_, r_n_491__16_, r_n_491__15_, r_n_491__14_, r_n_491__13_, r_n_491__12_, r_n_491__11_, r_n_491__10_, r_n_491__9_, r_n_491__8_, r_n_491__7_, r_n_491__6_, r_n_491__5_, r_n_491__4_, r_n_491__3_, r_n_491__2_, r_n_491__1_, r_n_491__0_ } = (N982)? { r_492__63_, r_492__62_, r_492__61_, r_492__60_, r_492__59_, r_492__58_, r_492__57_, r_492__56_, r_492__55_, r_492__54_, r_492__53_, r_492__52_, r_492__51_, r_492__50_, r_492__49_, r_492__48_, r_492__47_, r_492__46_, r_492__45_, r_492__44_, r_492__43_, r_492__42_, r_492__41_, r_492__40_, r_492__39_, r_492__38_, r_492__37_, r_492__36_, r_492__35_, r_492__34_, r_492__33_, r_492__32_, r_492__31_, r_492__30_, r_492__29_, r_492__28_, r_492__27_, r_492__26_, r_492__25_, r_492__24_, r_492__23_, r_492__22_, r_492__21_, r_492__20_, r_492__19_, r_492__18_, r_492__17_, r_492__16_, r_492__15_, r_492__14_, r_492__13_, r_492__12_, r_492__11_, r_492__10_, r_492__9_, r_492__8_, r_492__7_, r_492__6_, r_492__5_, r_492__4_, r_492__3_, r_492__2_, r_492__1_, r_492__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N983)? data_i : 1'b0;
  assign N982 = sel_i[982];
  assign N983 = N3483;
  assign { r_n_492__63_, r_n_492__62_, r_n_492__61_, r_n_492__60_, r_n_492__59_, r_n_492__58_, r_n_492__57_, r_n_492__56_, r_n_492__55_, r_n_492__54_, r_n_492__53_, r_n_492__52_, r_n_492__51_, r_n_492__50_, r_n_492__49_, r_n_492__48_, r_n_492__47_, r_n_492__46_, r_n_492__45_, r_n_492__44_, r_n_492__43_, r_n_492__42_, r_n_492__41_, r_n_492__40_, r_n_492__39_, r_n_492__38_, r_n_492__37_, r_n_492__36_, r_n_492__35_, r_n_492__34_, r_n_492__33_, r_n_492__32_, r_n_492__31_, r_n_492__30_, r_n_492__29_, r_n_492__28_, r_n_492__27_, r_n_492__26_, r_n_492__25_, r_n_492__24_, r_n_492__23_, r_n_492__22_, r_n_492__21_, r_n_492__20_, r_n_492__19_, r_n_492__18_, r_n_492__17_, r_n_492__16_, r_n_492__15_, r_n_492__14_, r_n_492__13_, r_n_492__12_, r_n_492__11_, r_n_492__10_, r_n_492__9_, r_n_492__8_, r_n_492__7_, r_n_492__6_, r_n_492__5_, r_n_492__4_, r_n_492__3_, r_n_492__2_, r_n_492__1_, r_n_492__0_ } = (N984)? { r_493__63_, r_493__62_, r_493__61_, r_493__60_, r_493__59_, r_493__58_, r_493__57_, r_493__56_, r_493__55_, r_493__54_, r_493__53_, r_493__52_, r_493__51_, r_493__50_, r_493__49_, r_493__48_, r_493__47_, r_493__46_, r_493__45_, r_493__44_, r_493__43_, r_493__42_, r_493__41_, r_493__40_, r_493__39_, r_493__38_, r_493__37_, r_493__36_, r_493__35_, r_493__34_, r_493__33_, r_493__32_, r_493__31_, r_493__30_, r_493__29_, r_493__28_, r_493__27_, r_493__26_, r_493__25_, r_493__24_, r_493__23_, r_493__22_, r_493__21_, r_493__20_, r_493__19_, r_493__18_, r_493__17_, r_493__16_, r_493__15_, r_493__14_, r_493__13_, r_493__12_, r_493__11_, r_493__10_, r_493__9_, r_493__8_, r_493__7_, r_493__6_, r_493__5_, r_493__4_, r_493__3_, r_493__2_, r_493__1_, r_493__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N985)? data_i : 1'b0;
  assign N984 = sel_i[984];
  assign N985 = N3488;
  assign { r_n_493__63_, r_n_493__62_, r_n_493__61_, r_n_493__60_, r_n_493__59_, r_n_493__58_, r_n_493__57_, r_n_493__56_, r_n_493__55_, r_n_493__54_, r_n_493__53_, r_n_493__52_, r_n_493__51_, r_n_493__50_, r_n_493__49_, r_n_493__48_, r_n_493__47_, r_n_493__46_, r_n_493__45_, r_n_493__44_, r_n_493__43_, r_n_493__42_, r_n_493__41_, r_n_493__40_, r_n_493__39_, r_n_493__38_, r_n_493__37_, r_n_493__36_, r_n_493__35_, r_n_493__34_, r_n_493__33_, r_n_493__32_, r_n_493__31_, r_n_493__30_, r_n_493__29_, r_n_493__28_, r_n_493__27_, r_n_493__26_, r_n_493__25_, r_n_493__24_, r_n_493__23_, r_n_493__22_, r_n_493__21_, r_n_493__20_, r_n_493__19_, r_n_493__18_, r_n_493__17_, r_n_493__16_, r_n_493__15_, r_n_493__14_, r_n_493__13_, r_n_493__12_, r_n_493__11_, r_n_493__10_, r_n_493__9_, r_n_493__8_, r_n_493__7_, r_n_493__6_, r_n_493__5_, r_n_493__4_, r_n_493__3_, r_n_493__2_, r_n_493__1_, r_n_493__0_ } = (N986)? { r_494__63_, r_494__62_, r_494__61_, r_494__60_, r_494__59_, r_494__58_, r_494__57_, r_494__56_, r_494__55_, r_494__54_, r_494__53_, r_494__52_, r_494__51_, r_494__50_, r_494__49_, r_494__48_, r_494__47_, r_494__46_, r_494__45_, r_494__44_, r_494__43_, r_494__42_, r_494__41_, r_494__40_, r_494__39_, r_494__38_, r_494__37_, r_494__36_, r_494__35_, r_494__34_, r_494__33_, r_494__32_, r_494__31_, r_494__30_, r_494__29_, r_494__28_, r_494__27_, r_494__26_, r_494__25_, r_494__24_, r_494__23_, r_494__22_, r_494__21_, r_494__20_, r_494__19_, r_494__18_, r_494__17_, r_494__16_, r_494__15_, r_494__14_, r_494__13_, r_494__12_, r_494__11_, r_494__10_, r_494__9_, r_494__8_, r_494__7_, r_494__6_, r_494__5_, r_494__4_, r_494__3_, r_494__2_, r_494__1_, r_494__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N987)? data_i : 1'b0;
  assign N986 = sel_i[986];
  assign N987 = N3493;
  assign { r_n_494__63_, r_n_494__62_, r_n_494__61_, r_n_494__60_, r_n_494__59_, r_n_494__58_, r_n_494__57_, r_n_494__56_, r_n_494__55_, r_n_494__54_, r_n_494__53_, r_n_494__52_, r_n_494__51_, r_n_494__50_, r_n_494__49_, r_n_494__48_, r_n_494__47_, r_n_494__46_, r_n_494__45_, r_n_494__44_, r_n_494__43_, r_n_494__42_, r_n_494__41_, r_n_494__40_, r_n_494__39_, r_n_494__38_, r_n_494__37_, r_n_494__36_, r_n_494__35_, r_n_494__34_, r_n_494__33_, r_n_494__32_, r_n_494__31_, r_n_494__30_, r_n_494__29_, r_n_494__28_, r_n_494__27_, r_n_494__26_, r_n_494__25_, r_n_494__24_, r_n_494__23_, r_n_494__22_, r_n_494__21_, r_n_494__20_, r_n_494__19_, r_n_494__18_, r_n_494__17_, r_n_494__16_, r_n_494__15_, r_n_494__14_, r_n_494__13_, r_n_494__12_, r_n_494__11_, r_n_494__10_, r_n_494__9_, r_n_494__8_, r_n_494__7_, r_n_494__6_, r_n_494__5_, r_n_494__4_, r_n_494__3_, r_n_494__2_, r_n_494__1_, r_n_494__0_ } = (N988)? { r_495__63_, r_495__62_, r_495__61_, r_495__60_, r_495__59_, r_495__58_, r_495__57_, r_495__56_, r_495__55_, r_495__54_, r_495__53_, r_495__52_, r_495__51_, r_495__50_, r_495__49_, r_495__48_, r_495__47_, r_495__46_, r_495__45_, r_495__44_, r_495__43_, r_495__42_, r_495__41_, r_495__40_, r_495__39_, r_495__38_, r_495__37_, r_495__36_, r_495__35_, r_495__34_, r_495__33_, r_495__32_, r_495__31_, r_495__30_, r_495__29_, r_495__28_, r_495__27_, r_495__26_, r_495__25_, r_495__24_, r_495__23_, r_495__22_, r_495__21_, r_495__20_, r_495__19_, r_495__18_, r_495__17_, r_495__16_, r_495__15_, r_495__14_, r_495__13_, r_495__12_, r_495__11_, r_495__10_, r_495__9_, r_495__8_, r_495__7_, r_495__6_, r_495__5_, r_495__4_, r_495__3_, r_495__2_, r_495__1_, r_495__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N989)? data_i : 1'b0;
  assign N988 = sel_i[988];
  assign N989 = N3498;
  assign { r_n_495__63_, r_n_495__62_, r_n_495__61_, r_n_495__60_, r_n_495__59_, r_n_495__58_, r_n_495__57_, r_n_495__56_, r_n_495__55_, r_n_495__54_, r_n_495__53_, r_n_495__52_, r_n_495__51_, r_n_495__50_, r_n_495__49_, r_n_495__48_, r_n_495__47_, r_n_495__46_, r_n_495__45_, r_n_495__44_, r_n_495__43_, r_n_495__42_, r_n_495__41_, r_n_495__40_, r_n_495__39_, r_n_495__38_, r_n_495__37_, r_n_495__36_, r_n_495__35_, r_n_495__34_, r_n_495__33_, r_n_495__32_, r_n_495__31_, r_n_495__30_, r_n_495__29_, r_n_495__28_, r_n_495__27_, r_n_495__26_, r_n_495__25_, r_n_495__24_, r_n_495__23_, r_n_495__22_, r_n_495__21_, r_n_495__20_, r_n_495__19_, r_n_495__18_, r_n_495__17_, r_n_495__16_, r_n_495__15_, r_n_495__14_, r_n_495__13_, r_n_495__12_, r_n_495__11_, r_n_495__10_, r_n_495__9_, r_n_495__8_, r_n_495__7_, r_n_495__6_, r_n_495__5_, r_n_495__4_, r_n_495__3_, r_n_495__2_, r_n_495__1_, r_n_495__0_ } = (N990)? { r_496__63_, r_496__62_, r_496__61_, r_496__60_, r_496__59_, r_496__58_, r_496__57_, r_496__56_, r_496__55_, r_496__54_, r_496__53_, r_496__52_, r_496__51_, r_496__50_, r_496__49_, r_496__48_, r_496__47_, r_496__46_, r_496__45_, r_496__44_, r_496__43_, r_496__42_, r_496__41_, r_496__40_, r_496__39_, r_496__38_, r_496__37_, r_496__36_, r_496__35_, r_496__34_, r_496__33_, r_496__32_, r_496__31_, r_496__30_, r_496__29_, r_496__28_, r_496__27_, r_496__26_, r_496__25_, r_496__24_, r_496__23_, r_496__22_, r_496__21_, r_496__20_, r_496__19_, r_496__18_, r_496__17_, r_496__16_, r_496__15_, r_496__14_, r_496__13_, r_496__12_, r_496__11_, r_496__10_, r_496__9_, r_496__8_, r_496__7_, r_496__6_, r_496__5_, r_496__4_, r_496__3_, r_496__2_, r_496__1_, r_496__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N991)? data_i : 1'b0;
  assign N990 = sel_i[990];
  assign N991 = N3503;
  assign { r_n_496__63_, r_n_496__62_, r_n_496__61_, r_n_496__60_, r_n_496__59_, r_n_496__58_, r_n_496__57_, r_n_496__56_, r_n_496__55_, r_n_496__54_, r_n_496__53_, r_n_496__52_, r_n_496__51_, r_n_496__50_, r_n_496__49_, r_n_496__48_, r_n_496__47_, r_n_496__46_, r_n_496__45_, r_n_496__44_, r_n_496__43_, r_n_496__42_, r_n_496__41_, r_n_496__40_, r_n_496__39_, r_n_496__38_, r_n_496__37_, r_n_496__36_, r_n_496__35_, r_n_496__34_, r_n_496__33_, r_n_496__32_, r_n_496__31_, r_n_496__30_, r_n_496__29_, r_n_496__28_, r_n_496__27_, r_n_496__26_, r_n_496__25_, r_n_496__24_, r_n_496__23_, r_n_496__22_, r_n_496__21_, r_n_496__20_, r_n_496__19_, r_n_496__18_, r_n_496__17_, r_n_496__16_, r_n_496__15_, r_n_496__14_, r_n_496__13_, r_n_496__12_, r_n_496__11_, r_n_496__10_, r_n_496__9_, r_n_496__8_, r_n_496__7_, r_n_496__6_, r_n_496__5_, r_n_496__4_, r_n_496__3_, r_n_496__2_, r_n_496__1_, r_n_496__0_ } = (N992)? { r_497__63_, r_497__62_, r_497__61_, r_497__60_, r_497__59_, r_497__58_, r_497__57_, r_497__56_, r_497__55_, r_497__54_, r_497__53_, r_497__52_, r_497__51_, r_497__50_, r_497__49_, r_497__48_, r_497__47_, r_497__46_, r_497__45_, r_497__44_, r_497__43_, r_497__42_, r_497__41_, r_497__40_, r_497__39_, r_497__38_, r_497__37_, r_497__36_, r_497__35_, r_497__34_, r_497__33_, r_497__32_, r_497__31_, r_497__30_, r_497__29_, r_497__28_, r_497__27_, r_497__26_, r_497__25_, r_497__24_, r_497__23_, r_497__22_, r_497__21_, r_497__20_, r_497__19_, r_497__18_, r_497__17_, r_497__16_, r_497__15_, r_497__14_, r_497__13_, r_497__12_, r_497__11_, r_497__10_, r_497__9_, r_497__8_, r_497__7_, r_497__6_, r_497__5_, r_497__4_, r_497__3_, r_497__2_, r_497__1_, r_497__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N993)? data_i : 1'b0;
  assign N992 = sel_i[992];
  assign N993 = N3508;
  assign { r_n_497__63_, r_n_497__62_, r_n_497__61_, r_n_497__60_, r_n_497__59_, r_n_497__58_, r_n_497__57_, r_n_497__56_, r_n_497__55_, r_n_497__54_, r_n_497__53_, r_n_497__52_, r_n_497__51_, r_n_497__50_, r_n_497__49_, r_n_497__48_, r_n_497__47_, r_n_497__46_, r_n_497__45_, r_n_497__44_, r_n_497__43_, r_n_497__42_, r_n_497__41_, r_n_497__40_, r_n_497__39_, r_n_497__38_, r_n_497__37_, r_n_497__36_, r_n_497__35_, r_n_497__34_, r_n_497__33_, r_n_497__32_, r_n_497__31_, r_n_497__30_, r_n_497__29_, r_n_497__28_, r_n_497__27_, r_n_497__26_, r_n_497__25_, r_n_497__24_, r_n_497__23_, r_n_497__22_, r_n_497__21_, r_n_497__20_, r_n_497__19_, r_n_497__18_, r_n_497__17_, r_n_497__16_, r_n_497__15_, r_n_497__14_, r_n_497__13_, r_n_497__12_, r_n_497__11_, r_n_497__10_, r_n_497__9_, r_n_497__8_, r_n_497__7_, r_n_497__6_, r_n_497__5_, r_n_497__4_, r_n_497__3_, r_n_497__2_, r_n_497__1_, r_n_497__0_ } = (N994)? { r_498__63_, r_498__62_, r_498__61_, r_498__60_, r_498__59_, r_498__58_, r_498__57_, r_498__56_, r_498__55_, r_498__54_, r_498__53_, r_498__52_, r_498__51_, r_498__50_, r_498__49_, r_498__48_, r_498__47_, r_498__46_, r_498__45_, r_498__44_, r_498__43_, r_498__42_, r_498__41_, r_498__40_, r_498__39_, r_498__38_, r_498__37_, r_498__36_, r_498__35_, r_498__34_, r_498__33_, r_498__32_, r_498__31_, r_498__30_, r_498__29_, r_498__28_, r_498__27_, r_498__26_, r_498__25_, r_498__24_, r_498__23_, r_498__22_, r_498__21_, r_498__20_, r_498__19_, r_498__18_, r_498__17_, r_498__16_, r_498__15_, r_498__14_, r_498__13_, r_498__12_, r_498__11_, r_498__10_, r_498__9_, r_498__8_, r_498__7_, r_498__6_, r_498__5_, r_498__4_, r_498__3_, r_498__2_, r_498__1_, r_498__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N995)? data_i : 1'b0;
  assign N994 = sel_i[994];
  assign N995 = N3513;
  assign { r_n_498__63_, r_n_498__62_, r_n_498__61_, r_n_498__60_, r_n_498__59_, r_n_498__58_, r_n_498__57_, r_n_498__56_, r_n_498__55_, r_n_498__54_, r_n_498__53_, r_n_498__52_, r_n_498__51_, r_n_498__50_, r_n_498__49_, r_n_498__48_, r_n_498__47_, r_n_498__46_, r_n_498__45_, r_n_498__44_, r_n_498__43_, r_n_498__42_, r_n_498__41_, r_n_498__40_, r_n_498__39_, r_n_498__38_, r_n_498__37_, r_n_498__36_, r_n_498__35_, r_n_498__34_, r_n_498__33_, r_n_498__32_, r_n_498__31_, r_n_498__30_, r_n_498__29_, r_n_498__28_, r_n_498__27_, r_n_498__26_, r_n_498__25_, r_n_498__24_, r_n_498__23_, r_n_498__22_, r_n_498__21_, r_n_498__20_, r_n_498__19_, r_n_498__18_, r_n_498__17_, r_n_498__16_, r_n_498__15_, r_n_498__14_, r_n_498__13_, r_n_498__12_, r_n_498__11_, r_n_498__10_, r_n_498__9_, r_n_498__8_, r_n_498__7_, r_n_498__6_, r_n_498__5_, r_n_498__4_, r_n_498__3_, r_n_498__2_, r_n_498__1_, r_n_498__0_ } = (N996)? { r_499__63_, r_499__62_, r_499__61_, r_499__60_, r_499__59_, r_499__58_, r_499__57_, r_499__56_, r_499__55_, r_499__54_, r_499__53_, r_499__52_, r_499__51_, r_499__50_, r_499__49_, r_499__48_, r_499__47_, r_499__46_, r_499__45_, r_499__44_, r_499__43_, r_499__42_, r_499__41_, r_499__40_, r_499__39_, r_499__38_, r_499__37_, r_499__36_, r_499__35_, r_499__34_, r_499__33_, r_499__32_, r_499__31_, r_499__30_, r_499__29_, r_499__28_, r_499__27_, r_499__26_, r_499__25_, r_499__24_, r_499__23_, r_499__22_, r_499__21_, r_499__20_, r_499__19_, r_499__18_, r_499__17_, r_499__16_, r_499__15_, r_499__14_, r_499__13_, r_499__12_, r_499__11_, r_499__10_, r_499__9_, r_499__8_, r_499__7_, r_499__6_, r_499__5_, r_499__4_, r_499__3_, r_499__2_, r_499__1_, r_499__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N997)? data_i : 1'b0;
  assign N996 = sel_i[996];
  assign N997 = N3518;
  assign { r_n_499__63_, r_n_499__62_, r_n_499__61_, r_n_499__60_, r_n_499__59_, r_n_499__58_, r_n_499__57_, r_n_499__56_, r_n_499__55_, r_n_499__54_, r_n_499__53_, r_n_499__52_, r_n_499__51_, r_n_499__50_, r_n_499__49_, r_n_499__48_, r_n_499__47_, r_n_499__46_, r_n_499__45_, r_n_499__44_, r_n_499__43_, r_n_499__42_, r_n_499__41_, r_n_499__40_, r_n_499__39_, r_n_499__38_, r_n_499__37_, r_n_499__36_, r_n_499__35_, r_n_499__34_, r_n_499__33_, r_n_499__32_, r_n_499__31_, r_n_499__30_, r_n_499__29_, r_n_499__28_, r_n_499__27_, r_n_499__26_, r_n_499__25_, r_n_499__24_, r_n_499__23_, r_n_499__22_, r_n_499__21_, r_n_499__20_, r_n_499__19_, r_n_499__18_, r_n_499__17_, r_n_499__16_, r_n_499__15_, r_n_499__14_, r_n_499__13_, r_n_499__12_, r_n_499__11_, r_n_499__10_, r_n_499__9_, r_n_499__8_, r_n_499__7_, r_n_499__6_, r_n_499__5_, r_n_499__4_, r_n_499__3_, r_n_499__2_, r_n_499__1_, r_n_499__0_ } = (N998)? { r_500__63_, r_500__62_, r_500__61_, r_500__60_, r_500__59_, r_500__58_, r_500__57_, r_500__56_, r_500__55_, r_500__54_, r_500__53_, r_500__52_, r_500__51_, r_500__50_, r_500__49_, r_500__48_, r_500__47_, r_500__46_, r_500__45_, r_500__44_, r_500__43_, r_500__42_, r_500__41_, r_500__40_, r_500__39_, r_500__38_, r_500__37_, r_500__36_, r_500__35_, r_500__34_, r_500__33_, r_500__32_, r_500__31_, r_500__30_, r_500__29_, r_500__28_, r_500__27_, r_500__26_, r_500__25_, r_500__24_, r_500__23_, r_500__22_, r_500__21_, r_500__20_, r_500__19_, r_500__18_, r_500__17_, r_500__16_, r_500__15_, r_500__14_, r_500__13_, r_500__12_, r_500__11_, r_500__10_, r_500__9_, r_500__8_, r_500__7_, r_500__6_, r_500__5_, r_500__4_, r_500__3_, r_500__2_, r_500__1_, r_500__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N999)? data_i : 1'b0;
  assign N998 = sel_i[998];
  assign N999 = N3523;
  assign { r_n_500__63_, r_n_500__62_, r_n_500__61_, r_n_500__60_, r_n_500__59_, r_n_500__58_, r_n_500__57_, r_n_500__56_, r_n_500__55_, r_n_500__54_, r_n_500__53_, r_n_500__52_, r_n_500__51_, r_n_500__50_, r_n_500__49_, r_n_500__48_, r_n_500__47_, r_n_500__46_, r_n_500__45_, r_n_500__44_, r_n_500__43_, r_n_500__42_, r_n_500__41_, r_n_500__40_, r_n_500__39_, r_n_500__38_, r_n_500__37_, r_n_500__36_, r_n_500__35_, r_n_500__34_, r_n_500__33_, r_n_500__32_, r_n_500__31_, r_n_500__30_, r_n_500__29_, r_n_500__28_, r_n_500__27_, r_n_500__26_, r_n_500__25_, r_n_500__24_, r_n_500__23_, r_n_500__22_, r_n_500__21_, r_n_500__20_, r_n_500__19_, r_n_500__18_, r_n_500__17_, r_n_500__16_, r_n_500__15_, r_n_500__14_, r_n_500__13_, r_n_500__12_, r_n_500__11_, r_n_500__10_, r_n_500__9_, r_n_500__8_, r_n_500__7_, r_n_500__6_, r_n_500__5_, r_n_500__4_, r_n_500__3_, r_n_500__2_, r_n_500__1_, r_n_500__0_ } = (N1000)? { r_501__63_, r_501__62_, r_501__61_, r_501__60_, r_501__59_, r_501__58_, r_501__57_, r_501__56_, r_501__55_, r_501__54_, r_501__53_, r_501__52_, r_501__51_, r_501__50_, r_501__49_, r_501__48_, r_501__47_, r_501__46_, r_501__45_, r_501__44_, r_501__43_, r_501__42_, r_501__41_, r_501__40_, r_501__39_, r_501__38_, r_501__37_, r_501__36_, r_501__35_, r_501__34_, r_501__33_, r_501__32_, r_501__31_, r_501__30_, r_501__29_, r_501__28_, r_501__27_, r_501__26_, r_501__25_, r_501__24_, r_501__23_, r_501__22_, r_501__21_, r_501__20_, r_501__19_, r_501__18_, r_501__17_, r_501__16_, r_501__15_, r_501__14_, r_501__13_, r_501__12_, r_501__11_, r_501__10_, r_501__9_, r_501__8_, r_501__7_, r_501__6_, r_501__5_, r_501__4_, r_501__3_, r_501__2_, r_501__1_, r_501__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N1001)? data_i : 1'b0;
  assign N1000 = sel_i[1000];
  assign N1001 = N3528;
  assign { r_n_501__63_, r_n_501__62_, r_n_501__61_, r_n_501__60_, r_n_501__59_, r_n_501__58_, r_n_501__57_, r_n_501__56_, r_n_501__55_, r_n_501__54_, r_n_501__53_, r_n_501__52_, r_n_501__51_, r_n_501__50_, r_n_501__49_, r_n_501__48_, r_n_501__47_, r_n_501__46_, r_n_501__45_, r_n_501__44_, r_n_501__43_, r_n_501__42_, r_n_501__41_, r_n_501__40_, r_n_501__39_, r_n_501__38_, r_n_501__37_, r_n_501__36_, r_n_501__35_, r_n_501__34_, r_n_501__33_, r_n_501__32_, r_n_501__31_, r_n_501__30_, r_n_501__29_, r_n_501__28_, r_n_501__27_, r_n_501__26_, r_n_501__25_, r_n_501__24_, r_n_501__23_, r_n_501__22_, r_n_501__21_, r_n_501__20_, r_n_501__19_, r_n_501__18_, r_n_501__17_, r_n_501__16_, r_n_501__15_, r_n_501__14_, r_n_501__13_, r_n_501__12_, r_n_501__11_, r_n_501__10_, r_n_501__9_, r_n_501__8_, r_n_501__7_, r_n_501__6_, r_n_501__5_, r_n_501__4_, r_n_501__3_, r_n_501__2_, r_n_501__1_, r_n_501__0_ } = (N1002)? { r_502__63_, r_502__62_, r_502__61_, r_502__60_, r_502__59_, r_502__58_, r_502__57_, r_502__56_, r_502__55_, r_502__54_, r_502__53_, r_502__52_, r_502__51_, r_502__50_, r_502__49_, r_502__48_, r_502__47_, r_502__46_, r_502__45_, r_502__44_, r_502__43_, r_502__42_, r_502__41_, r_502__40_, r_502__39_, r_502__38_, r_502__37_, r_502__36_, r_502__35_, r_502__34_, r_502__33_, r_502__32_, r_502__31_, r_502__30_, r_502__29_, r_502__28_, r_502__27_, r_502__26_, r_502__25_, r_502__24_, r_502__23_, r_502__22_, r_502__21_, r_502__20_, r_502__19_, r_502__18_, r_502__17_, r_502__16_, r_502__15_, r_502__14_, r_502__13_, r_502__12_, r_502__11_, r_502__10_, r_502__9_, r_502__8_, r_502__7_, r_502__6_, r_502__5_, r_502__4_, r_502__3_, r_502__2_, r_502__1_, r_502__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N1003)? data_i : 1'b0;
  assign N1002 = sel_i[1002];
  assign N1003 = N3533;
  assign { r_n_502__63_, r_n_502__62_, r_n_502__61_, r_n_502__60_, r_n_502__59_, r_n_502__58_, r_n_502__57_, r_n_502__56_, r_n_502__55_, r_n_502__54_, r_n_502__53_, r_n_502__52_, r_n_502__51_, r_n_502__50_, r_n_502__49_, r_n_502__48_, r_n_502__47_, r_n_502__46_, r_n_502__45_, r_n_502__44_, r_n_502__43_, r_n_502__42_, r_n_502__41_, r_n_502__40_, r_n_502__39_, r_n_502__38_, r_n_502__37_, r_n_502__36_, r_n_502__35_, r_n_502__34_, r_n_502__33_, r_n_502__32_, r_n_502__31_, r_n_502__30_, r_n_502__29_, r_n_502__28_, r_n_502__27_, r_n_502__26_, r_n_502__25_, r_n_502__24_, r_n_502__23_, r_n_502__22_, r_n_502__21_, r_n_502__20_, r_n_502__19_, r_n_502__18_, r_n_502__17_, r_n_502__16_, r_n_502__15_, r_n_502__14_, r_n_502__13_, r_n_502__12_, r_n_502__11_, r_n_502__10_, r_n_502__9_, r_n_502__8_, r_n_502__7_, r_n_502__6_, r_n_502__5_, r_n_502__4_, r_n_502__3_, r_n_502__2_, r_n_502__1_, r_n_502__0_ } = (N1004)? { r_503__63_, r_503__62_, r_503__61_, r_503__60_, r_503__59_, r_503__58_, r_503__57_, r_503__56_, r_503__55_, r_503__54_, r_503__53_, r_503__52_, r_503__51_, r_503__50_, r_503__49_, r_503__48_, r_503__47_, r_503__46_, r_503__45_, r_503__44_, r_503__43_, r_503__42_, r_503__41_, r_503__40_, r_503__39_, r_503__38_, r_503__37_, r_503__36_, r_503__35_, r_503__34_, r_503__33_, r_503__32_, r_503__31_, r_503__30_, r_503__29_, r_503__28_, r_503__27_, r_503__26_, r_503__25_, r_503__24_, r_503__23_, r_503__22_, r_503__21_, r_503__20_, r_503__19_, r_503__18_, r_503__17_, r_503__16_, r_503__15_, r_503__14_, r_503__13_, r_503__12_, r_503__11_, r_503__10_, r_503__9_, r_503__8_, r_503__7_, r_503__6_, r_503__5_, r_503__4_, r_503__3_, r_503__2_, r_503__1_, r_503__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N1005)? data_i : 1'b0;
  assign N1004 = sel_i[1004];
  assign N1005 = N3538;
  assign { r_n_503__63_, r_n_503__62_, r_n_503__61_, r_n_503__60_, r_n_503__59_, r_n_503__58_, r_n_503__57_, r_n_503__56_, r_n_503__55_, r_n_503__54_, r_n_503__53_, r_n_503__52_, r_n_503__51_, r_n_503__50_, r_n_503__49_, r_n_503__48_, r_n_503__47_, r_n_503__46_, r_n_503__45_, r_n_503__44_, r_n_503__43_, r_n_503__42_, r_n_503__41_, r_n_503__40_, r_n_503__39_, r_n_503__38_, r_n_503__37_, r_n_503__36_, r_n_503__35_, r_n_503__34_, r_n_503__33_, r_n_503__32_, r_n_503__31_, r_n_503__30_, r_n_503__29_, r_n_503__28_, r_n_503__27_, r_n_503__26_, r_n_503__25_, r_n_503__24_, r_n_503__23_, r_n_503__22_, r_n_503__21_, r_n_503__20_, r_n_503__19_, r_n_503__18_, r_n_503__17_, r_n_503__16_, r_n_503__15_, r_n_503__14_, r_n_503__13_, r_n_503__12_, r_n_503__11_, r_n_503__10_, r_n_503__9_, r_n_503__8_, r_n_503__7_, r_n_503__6_, r_n_503__5_, r_n_503__4_, r_n_503__3_, r_n_503__2_, r_n_503__1_, r_n_503__0_ } = (N1006)? { r_504__63_, r_504__62_, r_504__61_, r_504__60_, r_504__59_, r_504__58_, r_504__57_, r_504__56_, r_504__55_, r_504__54_, r_504__53_, r_504__52_, r_504__51_, r_504__50_, r_504__49_, r_504__48_, r_504__47_, r_504__46_, r_504__45_, r_504__44_, r_504__43_, r_504__42_, r_504__41_, r_504__40_, r_504__39_, r_504__38_, r_504__37_, r_504__36_, r_504__35_, r_504__34_, r_504__33_, r_504__32_, r_504__31_, r_504__30_, r_504__29_, r_504__28_, r_504__27_, r_504__26_, r_504__25_, r_504__24_, r_504__23_, r_504__22_, r_504__21_, r_504__20_, r_504__19_, r_504__18_, r_504__17_, r_504__16_, r_504__15_, r_504__14_, r_504__13_, r_504__12_, r_504__11_, r_504__10_, r_504__9_, r_504__8_, r_504__7_, r_504__6_, r_504__5_, r_504__4_, r_504__3_, r_504__2_, r_504__1_, r_504__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N1007)? data_i : 1'b0;
  assign N1006 = sel_i[1006];
  assign N1007 = N3543;
  assign { r_n_504__63_, r_n_504__62_, r_n_504__61_, r_n_504__60_, r_n_504__59_, r_n_504__58_, r_n_504__57_, r_n_504__56_, r_n_504__55_, r_n_504__54_, r_n_504__53_, r_n_504__52_, r_n_504__51_, r_n_504__50_, r_n_504__49_, r_n_504__48_, r_n_504__47_, r_n_504__46_, r_n_504__45_, r_n_504__44_, r_n_504__43_, r_n_504__42_, r_n_504__41_, r_n_504__40_, r_n_504__39_, r_n_504__38_, r_n_504__37_, r_n_504__36_, r_n_504__35_, r_n_504__34_, r_n_504__33_, r_n_504__32_, r_n_504__31_, r_n_504__30_, r_n_504__29_, r_n_504__28_, r_n_504__27_, r_n_504__26_, r_n_504__25_, r_n_504__24_, r_n_504__23_, r_n_504__22_, r_n_504__21_, r_n_504__20_, r_n_504__19_, r_n_504__18_, r_n_504__17_, r_n_504__16_, r_n_504__15_, r_n_504__14_, r_n_504__13_, r_n_504__12_, r_n_504__11_, r_n_504__10_, r_n_504__9_, r_n_504__8_, r_n_504__7_, r_n_504__6_, r_n_504__5_, r_n_504__4_, r_n_504__3_, r_n_504__2_, r_n_504__1_, r_n_504__0_ } = (N1008)? { r_505__63_, r_505__62_, r_505__61_, r_505__60_, r_505__59_, r_505__58_, r_505__57_, r_505__56_, r_505__55_, r_505__54_, r_505__53_, r_505__52_, r_505__51_, r_505__50_, r_505__49_, r_505__48_, r_505__47_, r_505__46_, r_505__45_, r_505__44_, r_505__43_, r_505__42_, r_505__41_, r_505__40_, r_505__39_, r_505__38_, r_505__37_, r_505__36_, r_505__35_, r_505__34_, r_505__33_, r_505__32_, r_505__31_, r_505__30_, r_505__29_, r_505__28_, r_505__27_, r_505__26_, r_505__25_, r_505__24_, r_505__23_, r_505__22_, r_505__21_, r_505__20_, r_505__19_, r_505__18_, r_505__17_, r_505__16_, r_505__15_, r_505__14_, r_505__13_, r_505__12_, r_505__11_, r_505__10_, r_505__9_, r_505__8_, r_505__7_, r_505__6_, r_505__5_, r_505__4_, r_505__3_, r_505__2_, r_505__1_, r_505__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N1009)? data_i : 1'b0;
  assign N1008 = sel_i[1008];
  assign N1009 = N3548;
  assign { r_n_505__63_, r_n_505__62_, r_n_505__61_, r_n_505__60_, r_n_505__59_, r_n_505__58_, r_n_505__57_, r_n_505__56_, r_n_505__55_, r_n_505__54_, r_n_505__53_, r_n_505__52_, r_n_505__51_, r_n_505__50_, r_n_505__49_, r_n_505__48_, r_n_505__47_, r_n_505__46_, r_n_505__45_, r_n_505__44_, r_n_505__43_, r_n_505__42_, r_n_505__41_, r_n_505__40_, r_n_505__39_, r_n_505__38_, r_n_505__37_, r_n_505__36_, r_n_505__35_, r_n_505__34_, r_n_505__33_, r_n_505__32_, r_n_505__31_, r_n_505__30_, r_n_505__29_, r_n_505__28_, r_n_505__27_, r_n_505__26_, r_n_505__25_, r_n_505__24_, r_n_505__23_, r_n_505__22_, r_n_505__21_, r_n_505__20_, r_n_505__19_, r_n_505__18_, r_n_505__17_, r_n_505__16_, r_n_505__15_, r_n_505__14_, r_n_505__13_, r_n_505__12_, r_n_505__11_, r_n_505__10_, r_n_505__9_, r_n_505__8_, r_n_505__7_, r_n_505__6_, r_n_505__5_, r_n_505__4_, r_n_505__3_, r_n_505__2_, r_n_505__1_, r_n_505__0_ } = (N1010)? { r_506__63_, r_506__62_, r_506__61_, r_506__60_, r_506__59_, r_506__58_, r_506__57_, r_506__56_, r_506__55_, r_506__54_, r_506__53_, r_506__52_, r_506__51_, r_506__50_, r_506__49_, r_506__48_, r_506__47_, r_506__46_, r_506__45_, r_506__44_, r_506__43_, r_506__42_, r_506__41_, r_506__40_, r_506__39_, r_506__38_, r_506__37_, r_506__36_, r_506__35_, r_506__34_, r_506__33_, r_506__32_, r_506__31_, r_506__30_, r_506__29_, r_506__28_, r_506__27_, r_506__26_, r_506__25_, r_506__24_, r_506__23_, r_506__22_, r_506__21_, r_506__20_, r_506__19_, r_506__18_, r_506__17_, r_506__16_, r_506__15_, r_506__14_, r_506__13_, r_506__12_, r_506__11_, r_506__10_, r_506__9_, r_506__8_, r_506__7_, r_506__6_, r_506__5_, r_506__4_, r_506__3_, r_506__2_, r_506__1_, r_506__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N1011)? data_i : 1'b0;
  assign N1010 = sel_i[1010];
  assign N1011 = N3553;
  assign { r_n_506__63_, r_n_506__62_, r_n_506__61_, r_n_506__60_, r_n_506__59_, r_n_506__58_, r_n_506__57_, r_n_506__56_, r_n_506__55_, r_n_506__54_, r_n_506__53_, r_n_506__52_, r_n_506__51_, r_n_506__50_, r_n_506__49_, r_n_506__48_, r_n_506__47_, r_n_506__46_, r_n_506__45_, r_n_506__44_, r_n_506__43_, r_n_506__42_, r_n_506__41_, r_n_506__40_, r_n_506__39_, r_n_506__38_, r_n_506__37_, r_n_506__36_, r_n_506__35_, r_n_506__34_, r_n_506__33_, r_n_506__32_, r_n_506__31_, r_n_506__30_, r_n_506__29_, r_n_506__28_, r_n_506__27_, r_n_506__26_, r_n_506__25_, r_n_506__24_, r_n_506__23_, r_n_506__22_, r_n_506__21_, r_n_506__20_, r_n_506__19_, r_n_506__18_, r_n_506__17_, r_n_506__16_, r_n_506__15_, r_n_506__14_, r_n_506__13_, r_n_506__12_, r_n_506__11_, r_n_506__10_, r_n_506__9_, r_n_506__8_, r_n_506__7_, r_n_506__6_, r_n_506__5_, r_n_506__4_, r_n_506__3_, r_n_506__2_, r_n_506__1_, r_n_506__0_ } = (N1012)? { r_507__63_, r_507__62_, r_507__61_, r_507__60_, r_507__59_, r_507__58_, r_507__57_, r_507__56_, r_507__55_, r_507__54_, r_507__53_, r_507__52_, r_507__51_, r_507__50_, r_507__49_, r_507__48_, r_507__47_, r_507__46_, r_507__45_, r_507__44_, r_507__43_, r_507__42_, r_507__41_, r_507__40_, r_507__39_, r_507__38_, r_507__37_, r_507__36_, r_507__35_, r_507__34_, r_507__33_, r_507__32_, r_507__31_, r_507__30_, r_507__29_, r_507__28_, r_507__27_, r_507__26_, r_507__25_, r_507__24_, r_507__23_, r_507__22_, r_507__21_, r_507__20_, r_507__19_, r_507__18_, r_507__17_, r_507__16_, r_507__15_, r_507__14_, r_507__13_, r_507__12_, r_507__11_, r_507__10_, r_507__9_, r_507__8_, r_507__7_, r_507__6_, r_507__5_, r_507__4_, r_507__3_, r_507__2_, r_507__1_, r_507__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N1013)? data_i : 1'b0;
  assign N1012 = sel_i[1012];
  assign N1013 = N3558;
  assign { r_n_507__63_, r_n_507__62_, r_n_507__61_, r_n_507__60_, r_n_507__59_, r_n_507__58_, r_n_507__57_, r_n_507__56_, r_n_507__55_, r_n_507__54_, r_n_507__53_, r_n_507__52_, r_n_507__51_, r_n_507__50_, r_n_507__49_, r_n_507__48_, r_n_507__47_, r_n_507__46_, r_n_507__45_, r_n_507__44_, r_n_507__43_, r_n_507__42_, r_n_507__41_, r_n_507__40_, r_n_507__39_, r_n_507__38_, r_n_507__37_, r_n_507__36_, r_n_507__35_, r_n_507__34_, r_n_507__33_, r_n_507__32_, r_n_507__31_, r_n_507__30_, r_n_507__29_, r_n_507__28_, r_n_507__27_, r_n_507__26_, r_n_507__25_, r_n_507__24_, r_n_507__23_, r_n_507__22_, r_n_507__21_, r_n_507__20_, r_n_507__19_, r_n_507__18_, r_n_507__17_, r_n_507__16_, r_n_507__15_, r_n_507__14_, r_n_507__13_, r_n_507__12_, r_n_507__11_, r_n_507__10_, r_n_507__9_, r_n_507__8_, r_n_507__7_, r_n_507__6_, r_n_507__5_, r_n_507__4_, r_n_507__3_, r_n_507__2_, r_n_507__1_, r_n_507__0_ } = (N1014)? { r_508__63_, r_508__62_, r_508__61_, r_508__60_, r_508__59_, r_508__58_, r_508__57_, r_508__56_, r_508__55_, r_508__54_, r_508__53_, r_508__52_, r_508__51_, r_508__50_, r_508__49_, r_508__48_, r_508__47_, r_508__46_, r_508__45_, r_508__44_, r_508__43_, r_508__42_, r_508__41_, r_508__40_, r_508__39_, r_508__38_, r_508__37_, r_508__36_, r_508__35_, r_508__34_, r_508__33_, r_508__32_, r_508__31_, r_508__30_, r_508__29_, r_508__28_, r_508__27_, r_508__26_, r_508__25_, r_508__24_, r_508__23_, r_508__22_, r_508__21_, r_508__20_, r_508__19_, r_508__18_, r_508__17_, r_508__16_, r_508__15_, r_508__14_, r_508__13_, r_508__12_, r_508__11_, r_508__10_, r_508__9_, r_508__8_, r_508__7_, r_508__6_, r_508__5_, r_508__4_, r_508__3_, r_508__2_, r_508__1_, r_508__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N1015)? data_i : 1'b0;
  assign N1014 = sel_i[1014];
  assign N1015 = N3563;
  assign { r_n_508__63_, r_n_508__62_, r_n_508__61_, r_n_508__60_, r_n_508__59_, r_n_508__58_, r_n_508__57_, r_n_508__56_, r_n_508__55_, r_n_508__54_, r_n_508__53_, r_n_508__52_, r_n_508__51_, r_n_508__50_, r_n_508__49_, r_n_508__48_, r_n_508__47_, r_n_508__46_, r_n_508__45_, r_n_508__44_, r_n_508__43_, r_n_508__42_, r_n_508__41_, r_n_508__40_, r_n_508__39_, r_n_508__38_, r_n_508__37_, r_n_508__36_, r_n_508__35_, r_n_508__34_, r_n_508__33_, r_n_508__32_, r_n_508__31_, r_n_508__30_, r_n_508__29_, r_n_508__28_, r_n_508__27_, r_n_508__26_, r_n_508__25_, r_n_508__24_, r_n_508__23_, r_n_508__22_, r_n_508__21_, r_n_508__20_, r_n_508__19_, r_n_508__18_, r_n_508__17_, r_n_508__16_, r_n_508__15_, r_n_508__14_, r_n_508__13_, r_n_508__12_, r_n_508__11_, r_n_508__10_, r_n_508__9_, r_n_508__8_, r_n_508__7_, r_n_508__6_, r_n_508__5_, r_n_508__4_, r_n_508__3_, r_n_508__2_, r_n_508__1_, r_n_508__0_ } = (N1016)? { r_509__63_, r_509__62_, r_509__61_, r_509__60_, r_509__59_, r_509__58_, r_509__57_, r_509__56_, r_509__55_, r_509__54_, r_509__53_, r_509__52_, r_509__51_, r_509__50_, r_509__49_, r_509__48_, r_509__47_, r_509__46_, r_509__45_, r_509__44_, r_509__43_, r_509__42_, r_509__41_, r_509__40_, r_509__39_, r_509__38_, r_509__37_, r_509__36_, r_509__35_, r_509__34_, r_509__33_, r_509__32_, r_509__31_, r_509__30_, r_509__29_, r_509__28_, r_509__27_, r_509__26_, r_509__25_, r_509__24_, r_509__23_, r_509__22_, r_509__21_, r_509__20_, r_509__19_, r_509__18_, r_509__17_, r_509__16_, r_509__15_, r_509__14_, r_509__13_, r_509__12_, r_509__11_, r_509__10_, r_509__9_, r_509__8_, r_509__7_, r_509__6_, r_509__5_, r_509__4_, r_509__3_, r_509__2_, r_509__1_, r_509__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N1017)? data_i : 1'b0;
  assign N1016 = sel_i[1016];
  assign N1017 = N3568;
  assign { r_n_509__63_, r_n_509__62_, r_n_509__61_, r_n_509__60_, r_n_509__59_, r_n_509__58_, r_n_509__57_, r_n_509__56_, r_n_509__55_, r_n_509__54_, r_n_509__53_, r_n_509__52_, r_n_509__51_, r_n_509__50_, r_n_509__49_, r_n_509__48_, r_n_509__47_, r_n_509__46_, r_n_509__45_, r_n_509__44_, r_n_509__43_, r_n_509__42_, r_n_509__41_, r_n_509__40_, r_n_509__39_, r_n_509__38_, r_n_509__37_, r_n_509__36_, r_n_509__35_, r_n_509__34_, r_n_509__33_, r_n_509__32_, r_n_509__31_, r_n_509__30_, r_n_509__29_, r_n_509__28_, r_n_509__27_, r_n_509__26_, r_n_509__25_, r_n_509__24_, r_n_509__23_, r_n_509__22_, r_n_509__21_, r_n_509__20_, r_n_509__19_, r_n_509__18_, r_n_509__17_, r_n_509__16_, r_n_509__15_, r_n_509__14_, r_n_509__13_, r_n_509__12_, r_n_509__11_, r_n_509__10_, r_n_509__9_, r_n_509__8_, r_n_509__7_, r_n_509__6_, r_n_509__5_, r_n_509__4_, r_n_509__3_, r_n_509__2_, r_n_509__1_, r_n_509__0_ } = (N1018)? { r_510__63_, r_510__62_, r_510__61_, r_510__60_, r_510__59_, r_510__58_, r_510__57_, r_510__56_, r_510__55_, r_510__54_, r_510__53_, r_510__52_, r_510__51_, r_510__50_, r_510__49_, r_510__48_, r_510__47_, r_510__46_, r_510__45_, r_510__44_, r_510__43_, r_510__42_, r_510__41_, r_510__40_, r_510__39_, r_510__38_, r_510__37_, r_510__36_, r_510__35_, r_510__34_, r_510__33_, r_510__32_, r_510__31_, r_510__30_, r_510__29_, r_510__28_, r_510__27_, r_510__26_, r_510__25_, r_510__24_, r_510__23_, r_510__22_, r_510__21_, r_510__20_, r_510__19_, r_510__18_, r_510__17_, r_510__16_, r_510__15_, r_510__14_, r_510__13_, r_510__12_, r_510__11_, r_510__10_, r_510__9_, r_510__8_, r_510__7_, r_510__6_, r_510__5_, r_510__4_, r_510__3_, r_510__2_, r_510__1_, r_510__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N1019)? data_i : 1'b0;
  assign N1018 = sel_i[1018];
  assign N1019 = N3573;
  assign { r_n_510__63_, r_n_510__62_, r_n_510__61_, r_n_510__60_, r_n_510__59_, r_n_510__58_, r_n_510__57_, r_n_510__56_, r_n_510__55_, r_n_510__54_, r_n_510__53_, r_n_510__52_, r_n_510__51_, r_n_510__50_, r_n_510__49_, r_n_510__48_, r_n_510__47_, r_n_510__46_, r_n_510__45_, r_n_510__44_, r_n_510__43_, r_n_510__42_, r_n_510__41_, r_n_510__40_, r_n_510__39_, r_n_510__38_, r_n_510__37_, r_n_510__36_, r_n_510__35_, r_n_510__34_, r_n_510__33_, r_n_510__32_, r_n_510__31_, r_n_510__30_, r_n_510__29_, r_n_510__28_, r_n_510__27_, r_n_510__26_, r_n_510__25_, r_n_510__24_, r_n_510__23_, r_n_510__22_, r_n_510__21_, r_n_510__20_, r_n_510__19_, r_n_510__18_, r_n_510__17_, r_n_510__16_, r_n_510__15_, r_n_510__14_, r_n_510__13_, r_n_510__12_, r_n_510__11_, r_n_510__10_, r_n_510__9_, r_n_510__8_, r_n_510__7_, r_n_510__6_, r_n_510__5_, r_n_510__4_, r_n_510__3_, r_n_510__2_, r_n_510__1_, r_n_510__0_ } = (N1020)? { r_511__63_, r_511__62_, r_511__61_, r_511__60_, r_511__59_, r_511__58_, r_511__57_, r_511__56_, r_511__55_, r_511__54_, r_511__53_, r_511__52_, r_511__51_, r_511__50_, r_511__49_, r_511__48_, r_511__47_, r_511__46_, r_511__45_, r_511__44_, r_511__43_, r_511__42_, r_511__41_, r_511__40_, r_511__39_, r_511__38_, r_511__37_, r_511__36_, r_511__35_, r_511__34_, r_511__33_, r_511__32_, r_511__31_, r_511__30_, r_511__29_, r_511__28_, r_511__27_, r_511__26_, r_511__25_, r_511__24_, r_511__23_, r_511__22_, r_511__21_, r_511__20_, r_511__19_, r_511__18_, r_511__17_, r_511__16_, r_511__15_, r_511__14_, r_511__13_, r_511__12_, r_511__11_, r_511__10_, r_511__9_, r_511__8_, r_511__7_, r_511__6_, r_511__5_, r_511__4_, r_511__3_, r_511__2_, r_511__1_, r_511__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N1021)? data_i : 1'b0;
  assign N1020 = sel_i[1020];
  assign N1021 = N3578;
  assign { r_n_511__63_, r_n_511__62_, r_n_511__61_, r_n_511__60_, r_n_511__59_, r_n_511__58_, r_n_511__57_, r_n_511__56_, r_n_511__55_, r_n_511__54_, r_n_511__53_, r_n_511__52_, r_n_511__51_, r_n_511__50_, r_n_511__49_, r_n_511__48_, r_n_511__47_, r_n_511__46_, r_n_511__45_, r_n_511__44_, r_n_511__43_, r_n_511__42_, r_n_511__41_, r_n_511__40_, r_n_511__39_, r_n_511__38_, r_n_511__37_, r_n_511__36_, r_n_511__35_, r_n_511__34_, r_n_511__33_, r_n_511__32_, r_n_511__31_, r_n_511__30_, r_n_511__29_, r_n_511__28_, r_n_511__27_, r_n_511__26_, r_n_511__25_, r_n_511__24_, r_n_511__23_, r_n_511__22_, r_n_511__21_, r_n_511__20_, r_n_511__19_, r_n_511__18_, r_n_511__17_, r_n_511__16_, r_n_511__15_, r_n_511__14_, r_n_511__13_, r_n_511__12_, r_n_511__11_, r_n_511__10_, r_n_511__9_, r_n_511__8_, r_n_511__7_, r_n_511__6_, r_n_511__5_, r_n_511__4_, r_n_511__3_, r_n_511__2_, r_n_511__1_, r_n_511__0_ } = (N1022)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N1023)? data_i : 1'b0;
  assign N1022 = sel_i[1022];
  assign N1023 = N3583;
  assign N1025 = ~sel_i[1];
  assign N1027 = N1024 | N1026;
  assign N1030 = ~sel_i[3];
  assign N1032 = N1029 | N1031;
  assign N1035 = ~sel_i[5];
  assign N1037 = N1034 | N1036;
  assign N1040 = ~sel_i[7];
  assign N1042 = N1039 | N1041;
  assign N1045 = ~sel_i[9];
  assign N1047 = N1044 | N1046;
  assign N1050 = ~sel_i[11];
  assign N1052 = N1049 | N1051;
  assign N1055 = ~sel_i[13];
  assign N1057 = N1054 | N1056;
  assign N1060 = ~sel_i[15];
  assign N1062 = N1059 | N1061;
  assign N1065 = ~sel_i[17];
  assign N1067 = N1064 | N1066;
  assign N1070 = ~sel_i[19];
  assign N1072 = N1069 | N1071;
  assign N1075 = ~sel_i[21];
  assign N1077 = N1074 | N1076;
  assign N1080 = ~sel_i[23];
  assign N1082 = N1079 | N1081;
  assign N1085 = ~sel_i[25];
  assign N1087 = N1084 | N1086;
  assign N1090 = ~sel_i[27];
  assign N1092 = N1089 | N1091;
  assign N1095 = ~sel_i[29];
  assign N1097 = N1094 | N1096;
  assign N1100 = ~sel_i[31];
  assign N1102 = N1099 | N1101;
  assign N1105 = ~sel_i[33];
  assign N1107 = N1104 | N1106;
  assign N1110 = ~sel_i[35];
  assign N1112 = N1109 | N1111;
  assign N1115 = ~sel_i[37];
  assign N1117 = N1114 | N1116;
  assign N1120 = ~sel_i[39];
  assign N1122 = N1119 | N1121;
  assign N1125 = ~sel_i[41];
  assign N1127 = N1124 | N1126;
  assign N1130 = ~sel_i[43];
  assign N1132 = N1129 | N1131;
  assign N1135 = ~sel_i[45];
  assign N1137 = N1134 | N1136;
  assign N1140 = ~sel_i[47];
  assign N1142 = N1139 | N1141;
  assign N1145 = ~sel_i[49];
  assign N1147 = N1144 | N1146;
  assign N1150 = ~sel_i[51];
  assign N1152 = N1149 | N1151;
  assign N1155 = ~sel_i[53];
  assign N1157 = N1154 | N1156;
  assign N1160 = ~sel_i[55];
  assign N1162 = N1159 | N1161;
  assign N1165 = ~sel_i[57];
  assign N1167 = N1164 | N1166;
  assign N1170 = ~sel_i[59];
  assign N1172 = N1169 | N1171;
  assign N1175 = ~sel_i[61];
  assign N1177 = N1174 | N1176;
  assign N1180 = ~sel_i[63];
  assign N1182 = N1179 | N1181;
  assign N1185 = ~sel_i[65];
  assign N1187 = N1184 | N1186;
  assign N1190 = ~sel_i[67];
  assign N1192 = N1189 | N1191;
  assign N1195 = ~sel_i[69];
  assign N1197 = N1194 | N1196;
  assign N1200 = ~sel_i[71];
  assign N1202 = N1199 | N1201;
  assign N1205 = ~sel_i[73];
  assign N1207 = N1204 | N1206;
  assign N1210 = ~sel_i[75];
  assign N1212 = N1209 | N1211;
  assign N1215 = ~sel_i[77];
  assign N1217 = N1214 | N1216;
  assign N1220 = ~sel_i[79];
  assign N1222 = N1219 | N1221;
  assign N1225 = ~sel_i[81];
  assign N1227 = N1224 | N1226;
  assign N1230 = ~sel_i[83];
  assign N1232 = N1229 | N1231;
  assign N1235 = ~sel_i[85];
  assign N1237 = N1234 | N1236;
  assign N1240 = ~sel_i[87];
  assign N1242 = N1239 | N1241;
  assign N1245 = ~sel_i[89];
  assign N1247 = N1244 | N1246;
  assign N1250 = ~sel_i[91];
  assign N1252 = N1249 | N1251;
  assign N1255 = ~sel_i[93];
  assign N1257 = N1254 | N1256;
  assign N1260 = ~sel_i[95];
  assign N1262 = N1259 | N1261;
  assign N1265 = ~sel_i[97];
  assign N1267 = N1264 | N1266;
  assign N1270 = ~sel_i[99];
  assign N1272 = N1269 | N1271;
  assign N1275 = ~sel_i[101];
  assign N1277 = N1274 | N1276;
  assign N1280 = ~sel_i[103];
  assign N1282 = N1279 | N1281;
  assign N1285 = ~sel_i[105];
  assign N1287 = N1284 | N1286;
  assign N1290 = ~sel_i[107];
  assign N1292 = N1289 | N1291;
  assign N1295 = ~sel_i[109];
  assign N1297 = N1294 | N1296;
  assign N1300 = ~sel_i[111];
  assign N1302 = N1299 | N1301;
  assign N1305 = ~sel_i[113];
  assign N1307 = N1304 | N1306;
  assign N1310 = ~sel_i[115];
  assign N1312 = N1309 | N1311;
  assign N1315 = ~sel_i[117];
  assign N1317 = N1314 | N1316;
  assign N1320 = ~sel_i[119];
  assign N1322 = N1319 | N1321;
  assign N1325 = ~sel_i[121];
  assign N1327 = N1324 | N1326;
  assign N1330 = ~sel_i[123];
  assign N1332 = N1329 | N1331;
  assign N1335 = ~sel_i[125];
  assign N1337 = N1334 | N1336;
  assign N1340 = ~sel_i[127];
  assign N1342 = N1339 | N1341;
  assign N1345 = ~sel_i[129];
  assign N1347 = N1344 | N1346;
  assign N1350 = ~sel_i[131];
  assign N1352 = N1349 | N1351;
  assign N1355 = ~sel_i[133];
  assign N1357 = N1354 | N1356;
  assign N1360 = ~sel_i[135];
  assign N1362 = N1359 | N1361;
  assign N1365 = ~sel_i[137];
  assign N1367 = N1364 | N1366;
  assign N1370 = ~sel_i[139];
  assign N1372 = N1369 | N1371;
  assign N1375 = ~sel_i[141];
  assign N1377 = N1374 | N1376;
  assign N1380 = ~sel_i[143];
  assign N1382 = N1379 | N1381;
  assign N1385 = ~sel_i[145];
  assign N1387 = N1384 | N1386;
  assign N1390 = ~sel_i[147];
  assign N1392 = N1389 | N1391;
  assign N1395 = ~sel_i[149];
  assign N1397 = N1394 | N1396;
  assign N1400 = ~sel_i[151];
  assign N1402 = N1399 | N1401;
  assign N1405 = ~sel_i[153];
  assign N1407 = N1404 | N1406;
  assign N1410 = ~sel_i[155];
  assign N1412 = N1409 | N1411;
  assign N1415 = ~sel_i[157];
  assign N1417 = N1414 | N1416;
  assign N1420 = ~sel_i[159];
  assign N1422 = N1419 | N1421;
  assign N1425 = ~sel_i[161];
  assign N1427 = N1424 | N1426;
  assign N1430 = ~sel_i[163];
  assign N1432 = N1429 | N1431;
  assign N1435 = ~sel_i[165];
  assign N1437 = N1434 | N1436;
  assign N1440 = ~sel_i[167];
  assign N1442 = N1439 | N1441;
  assign N1445 = ~sel_i[169];
  assign N1447 = N1444 | N1446;
  assign N1450 = ~sel_i[171];
  assign N1452 = N1449 | N1451;
  assign N1455 = ~sel_i[173];
  assign N1457 = N1454 | N1456;
  assign N1460 = ~sel_i[175];
  assign N1462 = N1459 | N1461;
  assign N1465 = ~sel_i[177];
  assign N1467 = N1464 | N1466;
  assign N1470 = ~sel_i[179];
  assign N1472 = N1469 | N1471;
  assign N1475 = ~sel_i[181];
  assign N1477 = N1474 | N1476;
  assign N1480 = ~sel_i[183];
  assign N1482 = N1479 | N1481;
  assign N1485 = ~sel_i[185];
  assign N1487 = N1484 | N1486;
  assign N1490 = ~sel_i[187];
  assign N1492 = N1489 | N1491;
  assign N1495 = ~sel_i[189];
  assign N1497 = N1494 | N1496;
  assign N1500 = ~sel_i[191];
  assign N1502 = N1499 | N1501;
  assign N1505 = ~sel_i[193];
  assign N1507 = N1504 | N1506;
  assign N1510 = ~sel_i[195];
  assign N1512 = N1509 | N1511;
  assign N1515 = ~sel_i[197];
  assign N1517 = N1514 | N1516;
  assign N1520 = ~sel_i[199];
  assign N1522 = N1519 | N1521;
  assign N1525 = ~sel_i[201];
  assign N1527 = N1524 | N1526;
  assign N1530 = ~sel_i[203];
  assign N1532 = N1529 | N1531;
  assign N1535 = ~sel_i[205];
  assign N1537 = N1534 | N1536;
  assign N1540 = ~sel_i[207];
  assign N1542 = N1539 | N1541;
  assign N1545 = ~sel_i[209];
  assign N1547 = N1544 | N1546;
  assign N1550 = ~sel_i[211];
  assign N1552 = N1549 | N1551;
  assign N1555 = ~sel_i[213];
  assign N1557 = N1554 | N1556;
  assign N1560 = ~sel_i[215];
  assign N1562 = N1559 | N1561;
  assign N1565 = ~sel_i[217];
  assign N1567 = N1564 | N1566;
  assign N1570 = ~sel_i[219];
  assign N1572 = N1569 | N1571;
  assign N1575 = ~sel_i[221];
  assign N1577 = N1574 | N1576;
  assign N1580 = ~sel_i[223];
  assign N1582 = N1579 | N1581;
  assign N1585 = ~sel_i[225];
  assign N1587 = N1584 | N1586;
  assign N1590 = ~sel_i[227];
  assign N1592 = N1589 | N1591;
  assign N1595 = ~sel_i[229];
  assign N1597 = N1594 | N1596;
  assign N1600 = ~sel_i[231];
  assign N1602 = N1599 | N1601;
  assign N1605 = ~sel_i[233];
  assign N1607 = N1604 | N1606;
  assign N1610 = ~sel_i[235];
  assign N1612 = N1609 | N1611;
  assign N1615 = ~sel_i[237];
  assign N1617 = N1614 | N1616;
  assign N1620 = ~sel_i[239];
  assign N1622 = N1619 | N1621;
  assign N1625 = ~sel_i[241];
  assign N1627 = N1624 | N1626;
  assign N1630 = ~sel_i[243];
  assign N1632 = N1629 | N1631;
  assign N1635 = ~sel_i[245];
  assign N1637 = N1634 | N1636;
  assign N1640 = ~sel_i[247];
  assign N1642 = N1639 | N1641;
  assign N1645 = ~sel_i[249];
  assign N1647 = N1644 | N1646;
  assign N1650 = ~sel_i[251];
  assign N1652 = N1649 | N1651;
  assign N1655 = ~sel_i[253];
  assign N1657 = N1654 | N1656;
  assign N1660 = ~sel_i[255];
  assign N1662 = N1659 | N1661;
  assign N1665 = ~sel_i[257];
  assign N1667 = N1664 | N1666;
  assign N1670 = ~sel_i[259];
  assign N1672 = N1669 | N1671;
  assign N1675 = ~sel_i[261];
  assign N1677 = N1674 | N1676;
  assign N1680 = ~sel_i[263];
  assign N1682 = N1679 | N1681;
  assign N1685 = ~sel_i[265];
  assign N1687 = N1684 | N1686;
  assign N1690 = ~sel_i[267];
  assign N1692 = N1689 | N1691;
  assign N1695 = ~sel_i[269];
  assign N1697 = N1694 | N1696;
  assign N1700 = ~sel_i[271];
  assign N1702 = N1699 | N1701;
  assign N1705 = ~sel_i[273];
  assign N1707 = N1704 | N1706;
  assign N1710 = ~sel_i[275];
  assign N1712 = N1709 | N1711;
  assign N1715 = ~sel_i[277];
  assign N1717 = N1714 | N1716;
  assign N1720 = ~sel_i[279];
  assign N1722 = N1719 | N1721;
  assign N1725 = ~sel_i[281];
  assign N1727 = N1724 | N1726;
  assign N1730 = ~sel_i[283];
  assign N1732 = N1729 | N1731;
  assign N1735 = ~sel_i[285];
  assign N1737 = N1734 | N1736;
  assign N1740 = ~sel_i[287];
  assign N1742 = N1739 | N1741;
  assign N1745 = ~sel_i[289];
  assign N1747 = N1744 | N1746;
  assign N1750 = ~sel_i[291];
  assign N1752 = N1749 | N1751;
  assign N1755 = ~sel_i[293];
  assign N1757 = N1754 | N1756;
  assign N1760 = ~sel_i[295];
  assign N1762 = N1759 | N1761;
  assign N1765 = ~sel_i[297];
  assign N1767 = N1764 | N1766;
  assign N1770 = ~sel_i[299];
  assign N1772 = N1769 | N1771;
  assign N1775 = ~sel_i[301];
  assign N1777 = N1774 | N1776;
  assign N1780 = ~sel_i[303];
  assign N1782 = N1779 | N1781;
  assign N1785 = ~sel_i[305];
  assign N1787 = N1784 | N1786;
  assign N1790 = ~sel_i[307];
  assign N1792 = N1789 | N1791;
  assign N1795 = ~sel_i[309];
  assign N1797 = N1794 | N1796;
  assign N1800 = ~sel_i[311];
  assign N1802 = N1799 | N1801;
  assign N1805 = ~sel_i[313];
  assign N1807 = N1804 | N1806;
  assign N1810 = ~sel_i[315];
  assign N1812 = N1809 | N1811;
  assign N1815 = ~sel_i[317];
  assign N1817 = N1814 | N1816;
  assign N1820 = ~sel_i[319];
  assign N1822 = N1819 | N1821;
  assign N1825 = ~sel_i[321];
  assign N1827 = N1824 | N1826;
  assign N1830 = ~sel_i[323];
  assign N1832 = N1829 | N1831;
  assign N1835 = ~sel_i[325];
  assign N1837 = N1834 | N1836;
  assign N1840 = ~sel_i[327];
  assign N1842 = N1839 | N1841;
  assign N1845 = ~sel_i[329];
  assign N1847 = N1844 | N1846;
  assign N1850 = ~sel_i[331];
  assign N1852 = N1849 | N1851;
  assign N1855 = ~sel_i[333];
  assign N1857 = N1854 | N1856;
  assign N1860 = ~sel_i[335];
  assign N1862 = N1859 | N1861;
  assign N1865 = ~sel_i[337];
  assign N1867 = N1864 | N1866;
  assign N1870 = ~sel_i[339];
  assign N1872 = N1869 | N1871;
  assign N1875 = ~sel_i[341];
  assign N1877 = N1874 | N1876;
  assign N1880 = ~sel_i[343];
  assign N1882 = N1879 | N1881;
  assign N1885 = ~sel_i[345];
  assign N1887 = N1884 | N1886;
  assign N1890 = ~sel_i[347];
  assign N1892 = N1889 | N1891;
  assign N1895 = ~sel_i[349];
  assign N1897 = N1894 | N1896;
  assign N1900 = ~sel_i[351];
  assign N1902 = N1899 | N1901;
  assign N1905 = ~sel_i[353];
  assign N1907 = N1904 | N1906;
  assign N1910 = ~sel_i[355];
  assign N1912 = N1909 | N1911;
  assign N1915 = ~sel_i[357];
  assign N1917 = N1914 | N1916;
  assign N1920 = ~sel_i[359];
  assign N1922 = N1919 | N1921;
  assign N1925 = ~sel_i[361];
  assign N1927 = N1924 | N1926;
  assign N1930 = ~sel_i[363];
  assign N1932 = N1929 | N1931;
  assign N1935 = ~sel_i[365];
  assign N1937 = N1934 | N1936;
  assign N1940 = ~sel_i[367];
  assign N1942 = N1939 | N1941;
  assign N1945 = ~sel_i[369];
  assign N1947 = N1944 | N1946;
  assign N1950 = ~sel_i[371];
  assign N1952 = N1949 | N1951;
  assign N1955 = ~sel_i[373];
  assign N1957 = N1954 | N1956;
  assign N1960 = ~sel_i[375];
  assign N1962 = N1959 | N1961;
  assign N1965 = ~sel_i[377];
  assign N1967 = N1964 | N1966;
  assign N1970 = ~sel_i[379];
  assign N1972 = N1969 | N1971;
  assign N1975 = ~sel_i[381];
  assign N1977 = N1974 | N1976;
  assign N1980 = ~sel_i[383];
  assign N1982 = N1979 | N1981;
  assign N1985 = ~sel_i[385];
  assign N1987 = N1984 | N1986;
  assign N1990 = ~sel_i[387];
  assign N1992 = N1989 | N1991;
  assign N1995 = ~sel_i[389];
  assign N1997 = N1994 | N1996;
  assign N2000 = ~sel_i[391];
  assign N2002 = N1999 | N2001;
  assign N2005 = ~sel_i[393];
  assign N2007 = N2004 | N2006;
  assign N2010 = ~sel_i[395];
  assign N2012 = N2009 | N2011;
  assign N2015 = ~sel_i[397];
  assign N2017 = N2014 | N2016;
  assign N2020 = ~sel_i[399];
  assign N2022 = N2019 | N2021;
  assign N2025 = ~sel_i[401];
  assign N2027 = N2024 | N2026;
  assign N2030 = ~sel_i[403];
  assign N2032 = N2029 | N2031;
  assign N2035 = ~sel_i[405];
  assign N2037 = N2034 | N2036;
  assign N2040 = ~sel_i[407];
  assign N2042 = N2039 | N2041;
  assign N2045 = ~sel_i[409];
  assign N2047 = N2044 | N2046;
  assign N2050 = ~sel_i[411];
  assign N2052 = N2049 | N2051;
  assign N2055 = ~sel_i[413];
  assign N2057 = N2054 | N2056;
  assign N2060 = ~sel_i[415];
  assign N2062 = N2059 | N2061;
  assign N2065 = ~sel_i[417];
  assign N2067 = N2064 | N2066;
  assign N2070 = ~sel_i[419];
  assign N2072 = N2069 | N2071;
  assign N2075 = ~sel_i[421];
  assign N2077 = N2074 | N2076;
  assign N2080 = ~sel_i[423];
  assign N2082 = N2079 | N2081;
  assign N2085 = ~sel_i[425];
  assign N2087 = N2084 | N2086;
  assign N2090 = ~sel_i[427];
  assign N2092 = N2089 | N2091;
  assign N2095 = ~sel_i[429];
  assign N2097 = N2094 | N2096;
  assign N2100 = ~sel_i[431];
  assign N2102 = N2099 | N2101;
  assign N2105 = ~sel_i[433];
  assign N2107 = N2104 | N2106;
  assign N2110 = ~sel_i[435];
  assign N2112 = N2109 | N2111;
  assign N2115 = ~sel_i[437];
  assign N2117 = N2114 | N2116;
  assign N2120 = ~sel_i[439];
  assign N2122 = N2119 | N2121;
  assign N2125 = ~sel_i[441];
  assign N2127 = N2124 | N2126;
  assign N2130 = ~sel_i[443];
  assign N2132 = N2129 | N2131;
  assign N2135 = ~sel_i[445];
  assign N2137 = N2134 | N2136;
  assign N2140 = ~sel_i[447];
  assign N2142 = N2139 | N2141;
  assign N2145 = ~sel_i[449];
  assign N2147 = N2144 | N2146;
  assign N2150 = ~sel_i[451];
  assign N2152 = N2149 | N2151;
  assign N2155 = ~sel_i[453];
  assign N2157 = N2154 | N2156;
  assign N2160 = ~sel_i[455];
  assign N2162 = N2159 | N2161;
  assign N2165 = ~sel_i[457];
  assign N2167 = N2164 | N2166;
  assign N2170 = ~sel_i[459];
  assign N2172 = N2169 | N2171;
  assign N2175 = ~sel_i[461];
  assign N2177 = N2174 | N2176;
  assign N2180 = ~sel_i[463];
  assign N2182 = N2179 | N2181;
  assign N2185 = ~sel_i[465];
  assign N2187 = N2184 | N2186;
  assign N2190 = ~sel_i[467];
  assign N2192 = N2189 | N2191;
  assign N2195 = ~sel_i[469];
  assign N2197 = N2194 | N2196;
  assign N2200 = ~sel_i[471];
  assign N2202 = N2199 | N2201;
  assign N2205 = ~sel_i[473];
  assign N2207 = N2204 | N2206;
  assign N2210 = ~sel_i[475];
  assign N2212 = N2209 | N2211;
  assign N2215 = ~sel_i[477];
  assign N2217 = N2214 | N2216;
  assign N2220 = ~sel_i[479];
  assign N2222 = N2219 | N2221;
  assign N2225 = ~sel_i[481];
  assign N2227 = N2224 | N2226;
  assign N2230 = ~sel_i[483];
  assign N2232 = N2229 | N2231;
  assign N2235 = ~sel_i[485];
  assign N2237 = N2234 | N2236;
  assign N2240 = ~sel_i[487];
  assign N2242 = N2239 | N2241;
  assign N2245 = ~sel_i[489];
  assign N2247 = N2244 | N2246;
  assign N2250 = ~sel_i[491];
  assign N2252 = N2249 | N2251;
  assign N2255 = ~sel_i[493];
  assign N2257 = N2254 | N2256;
  assign N2260 = ~sel_i[495];
  assign N2262 = N2259 | N2261;
  assign N2265 = ~sel_i[497];
  assign N2267 = N2264 | N2266;
  assign N2270 = ~sel_i[499];
  assign N2272 = N2269 | N2271;
  assign N2275 = ~sel_i[501];
  assign N2277 = N2274 | N2276;
  assign N2280 = ~sel_i[503];
  assign N2282 = N2279 | N2281;
  assign N2285 = ~sel_i[505];
  assign N2287 = N2284 | N2286;
  assign N2290 = ~sel_i[507];
  assign N2292 = N2289 | N2291;
  assign N2295 = ~sel_i[509];
  assign N2297 = N2294 | N2296;
  assign N2300 = ~sel_i[511];
  assign N2302 = N2299 | N2301;
  assign N2305 = ~sel_i[513];
  assign N2307 = N2304 | N2306;
  assign N2310 = ~sel_i[515];
  assign N2312 = N2309 | N2311;
  assign N2315 = ~sel_i[517];
  assign N2317 = N2314 | N2316;
  assign N2320 = ~sel_i[519];
  assign N2322 = N2319 | N2321;
  assign N2325 = ~sel_i[521];
  assign N2327 = N2324 | N2326;
  assign N2330 = ~sel_i[523];
  assign N2332 = N2329 | N2331;
  assign N2335 = ~sel_i[525];
  assign N2337 = N2334 | N2336;
  assign N2340 = ~sel_i[527];
  assign N2342 = N2339 | N2341;
  assign N2345 = ~sel_i[529];
  assign N2347 = N2344 | N2346;
  assign N2350 = ~sel_i[531];
  assign N2352 = N2349 | N2351;
  assign N2355 = ~sel_i[533];
  assign N2357 = N2354 | N2356;
  assign N2360 = ~sel_i[535];
  assign N2362 = N2359 | N2361;
  assign N2365 = ~sel_i[537];
  assign N2367 = N2364 | N2366;
  assign N2370 = ~sel_i[539];
  assign N2372 = N2369 | N2371;
  assign N2375 = ~sel_i[541];
  assign N2377 = N2374 | N2376;
  assign N2380 = ~sel_i[543];
  assign N2382 = N2379 | N2381;
  assign N2385 = ~sel_i[545];
  assign N2387 = N2384 | N2386;
  assign N2390 = ~sel_i[547];
  assign N2392 = N2389 | N2391;
  assign N2395 = ~sel_i[549];
  assign N2397 = N2394 | N2396;
  assign N2400 = ~sel_i[551];
  assign N2402 = N2399 | N2401;
  assign N2405 = ~sel_i[553];
  assign N2407 = N2404 | N2406;
  assign N2410 = ~sel_i[555];
  assign N2412 = N2409 | N2411;
  assign N2415 = ~sel_i[557];
  assign N2417 = N2414 | N2416;
  assign N2420 = ~sel_i[559];
  assign N2422 = N2419 | N2421;
  assign N2425 = ~sel_i[561];
  assign N2427 = N2424 | N2426;
  assign N2430 = ~sel_i[563];
  assign N2432 = N2429 | N2431;
  assign N2435 = ~sel_i[565];
  assign N2437 = N2434 | N2436;
  assign N2440 = ~sel_i[567];
  assign N2442 = N2439 | N2441;
  assign N2445 = ~sel_i[569];
  assign N2447 = N2444 | N2446;
  assign N2450 = ~sel_i[571];
  assign N2452 = N2449 | N2451;
  assign N2455 = ~sel_i[573];
  assign N2457 = N2454 | N2456;
  assign N2460 = ~sel_i[575];
  assign N2462 = N2459 | N2461;
  assign N2465 = ~sel_i[577];
  assign N2467 = N2464 | N2466;
  assign N2470 = ~sel_i[579];
  assign N2472 = N2469 | N2471;
  assign N2475 = ~sel_i[581];
  assign N2477 = N2474 | N2476;
  assign N2480 = ~sel_i[583];
  assign N2482 = N2479 | N2481;
  assign N2485 = ~sel_i[585];
  assign N2487 = N2484 | N2486;
  assign N2490 = ~sel_i[587];
  assign N2492 = N2489 | N2491;
  assign N2495 = ~sel_i[589];
  assign N2497 = N2494 | N2496;
  assign N2500 = ~sel_i[591];
  assign N2502 = N2499 | N2501;
  assign N2505 = ~sel_i[593];
  assign N2507 = N2504 | N2506;
  assign N2510 = ~sel_i[595];
  assign N2512 = N2509 | N2511;
  assign N2515 = ~sel_i[597];
  assign N2517 = N2514 | N2516;
  assign N2520 = ~sel_i[599];
  assign N2522 = N2519 | N2521;
  assign N2525 = ~sel_i[601];
  assign N2527 = N2524 | N2526;
  assign N2530 = ~sel_i[603];
  assign N2532 = N2529 | N2531;
  assign N2535 = ~sel_i[605];
  assign N2537 = N2534 | N2536;
  assign N2540 = ~sel_i[607];
  assign N2542 = N2539 | N2541;
  assign N2545 = ~sel_i[609];
  assign N2547 = N2544 | N2546;
  assign N2550 = ~sel_i[611];
  assign N2552 = N2549 | N2551;
  assign N2555 = ~sel_i[613];
  assign N2557 = N2554 | N2556;
  assign N2560 = ~sel_i[615];
  assign N2562 = N2559 | N2561;
  assign N2565 = ~sel_i[617];
  assign N2567 = N2564 | N2566;
  assign N2570 = ~sel_i[619];
  assign N2572 = N2569 | N2571;
  assign N2575 = ~sel_i[621];
  assign N2577 = N2574 | N2576;
  assign N2580 = ~sel_i[623];
  assign N2582 = N2579 | N2581;
  assign N2585 = ~sel_i[625];
  assign N2587 = N2584 | N2586;
  assign N2590 = ~sel_i[627];
  assign N2592 = N2589 | N2591;
  assign N2595 = ~sel_i[629];
  assign N2597 = N2594 | N2596;
  assign N2600 = ~sel_i[631];
  assign N2602 = N2599 | N2601;
  assign N2605 = ~sel_i[633];
  assign N2607 = N2604 | N2606;
  assign N2610 = ~sel_i[635];
  assign N2612 = N2609 | N2611;
  assign N2615 = ~sel_i[637];
  assign N2617 = N2614 | N2616;
  assign N2620 = ~sel_i[639];
  assign N2622 = N2619 | N2621;
  assign N2625 = ~sel_i[641];
  assign N2627 = N2624 | N2626;
  assign N2630 = ~sel_i[643];
  assign N2632 = N2629 | N2631;
  assign N2635 = ~sel_i[645];
  assign N2637 = N2634 | N2636;
  assign N2640 = ~sel_i[647];
  assign N2642 = N2639 | N2641;
  assign N2645 = ~sel_i[649];
  assign N2647 = N2644 | N2646;
  assign N2650 = ~sel_i[651];
  assign N2652 = N2649 | N2651;
  assign N2655 = ~sel_i[653];
  assign N2657 = N2654 | N2656;
  assign N2660 = ~sel_i[655];
  assign N2662 = N2659 | N2661;
  assign N2665 = ~sel_i[657];
  assign N2667 = N2664 | N2666;
  assign N2670 = ~sel_i[659];
  assign N2672 = N2669 | N2671;
  assign N2675 = ~sel_i[661];
  assign N2677 = N2674 | N2676;
  assign N2680 = ~sel_i[663];
  assign N2682 = N2679 | N2681;
  assign N2685 = ~sel_i[665];
  assign N2687 = N2684 | N2686;
  assign N2690 = ~sel_i[667];
  assign N2692 = N2689 | N2691;
  assign N2695 = ~sel_i[669];
  assign N2697 = N2694 | N2696;
  assign N2700 = ~sel_i[671];
  assign N2702 = N2699 | N2701;
  assign N2705 = ~sel_i[673];
  assign N2707 = N2704 | N2706;
  assign N2710 = ~sel_i[675];
  assign N2712 = N2709 | N2711;
  assign N2715 = ~sel_i[677];
  assign N2717 = N2714 | N2716;
  assign N2720 = ~sel_i[679];
  assign N2722 = N2719 | N2721;
  assign N2725 = ~sel_i[681];
  assign N2727 = N2724 | N2726;
  assign N2730 = ~sel_i[683];
  assign N2732 = N2729 | N2731;
  assign N2735 = ~sel_i[685];
  assign N2737 = N2734 | N2736;
  assign N2740 = ~sel_i[687];
  assign N2742 = N2739 | N2741;
  assign N2745 = ~sel_i[689];
  assign N2747 = N2744 | N2746;
  assign N2750 = ~sel_i[691];
  assign N2752 = N2749 | N2751;
  assign N2755 = ~sel_i[693];
  assign N2757 = N2754 | N2756;
  assign N2760 = ~sel_i[695];
  assign N2762 = N2759 | N2761;
  assign N2765 = ~sel_i[697];
  assign N2767 = N2764 | N2766;
  assign N2770 = ~sel_i[699];
  assign N2772 = N2769 | N2771;
  assign N2775 = ~sel_i[701];
  assign N2777 = N2774 | N2776;
  assign N2780 = ~sel_i[703];
  assign N2782 = N2779 | N2781;
  assign N2785 = ~sel_i[705];
  assign N2787 = N2784 | N2786;
  assign N2790 = ~sel_i[707];
  assign N2792 = N2789 | N2791;
  assign N2795 = ~sel_i[709];
  assign N2797 = N2794 | N2796;
  assign N2800 = ~sel_i[711];
  assign N2802 = N2799 | N2801;
  assign N2805 = ~sel_i[713];
  assign N2807 = N2804 | N2806;
  assign N2810 = ~sel_i[715];
  assign N2812 = N2809 | N2811;
  assign N2815 = ~sel_i[717];
  assign N2817 = N2814 | N2816;
  assign N2820 = ~sel_i[719];
  assign N2822 = N2819 | N2821;
  assign N2825 = ~sel_i[721];
  assign N2827 = N2824 | N2826;
  assign N2830 = ~sel_i[723];
  assign N2832 = N2829 | N2831;
  assign N2835 = ~sel_i[725];
  assign N2837 = N2834 | N2836;
  assign N2840 = ~sel_i[727];
  assign N2842 = N2839 | N2841;
  assign N2845 = ~sel_i[729];
  assign N2847 = N2844 | N2846;
  assign N2850 = ~sel_i[731];
  assign N2852 = N2849 | N2851;
  assign N2855 = ~sel_i[733];
  assign N2857 = N2854 | N2856;
  assign N2860 = ~sel_i[735];
  assign N2862 = N2859 | N2861;
  assign N2865 = ~sel_i[737];
  assign N2867 = N2864 | N2866;
  assign N2870 = ~sel_i[739];
  assign N2872 = N2869 | N2871;
  assign N2875 = ~sel_i[741];
  assign N2877 = N2874 | N2876;
  assign N2880 = ~sel_i[743];
  assign N2882 = N2879 | N2881;
  assign N2885 = ~sel_i[745];
  assign N2887 = N2884 | N2886;
  assign N2890 = ~sel_i[747];
  assign N2892 = N2889 | N2891;
  assign N2895 = ~sel_i[749];
  assign N2897 = N2894 | N2896;
  assign N2900 = ~sel_i[751];
  assign N2902 = N2899 | N2901;
  assign N2905 = ~sel_i[753];
  assign N2907 = N2904 | N2906;
  assign N2910 = ~sel_i[755];
  assign N2912 = N2909 | N2911;
  assign N2915 = ~sel_i[757];
  assign N2917 = N2914 | N2916;
  assign N2920 = ~sel_i[759];
  assign N2922 = N2919 | N2921;
  assign N2925 = ~sel_i[761];
  assign N2927 = N2924 | N2926;
  assign N2930 = ~sel_i[763];
  assign N2932 = N2929 | N2931;
  assign N2935 = ~sel_i[765];
  assign N2937 = N2934 | N2936;
  assign N2940 = ~sel_i[767];
  assign N2942 = N2939 | N2941;
  assign N2945 = ~sel_i[769];
  assign N2947 = N2944 | N2946;
  assign N2950 = ~sel_i[771];
  assign N2952 = N2949 | N2951;
  assign N2955 = ~sel_i[773];
  assign N2957 = N2954 | N2956;
  assign N2960 = ~sel_i[775];
  assign N2962 = N2959 | N2961;
  assign N2965 = ~sel_i[777];
  assign N2967 = N2964 | N2966;
  assign N2970 = ~sel_i[779];
  assign N2972 = N2969 | N2971;
  assign N2975 = ~sel_i[781];
  assign N2977 = N2974 | N2976;
  assign N2980 = ~sel_i[783];
  assign N2982 = N2979 | N2981;
  assign N2985 = ~sel_i[785];
  assign N2987 = N2984 | N2986;
  assign N2990 = ~sel_i[787];
  assign N2992 = N2989 | N2991;
  assign N2995 = ~sel_i[789];
  assign N2997 = N2994 | N2996;
  assign N3000 = ~sel_i[791];
  assign N3002 = N2999 | N3001;
  assign N3005 = ~sel_i[793];
  assign N3007 = N3004 | N3006;
  assign N3010 = ~sel_i[795];
  assign N3012 = N3009 | N3011;
  assign N3015 = ~sel_i[797];
  assign N3017 = N3014 | N3016;
  assign N3020 = ~sel_i[799];
  assign N3022 = N3019 | N3021;
  assign N3025 = ~sel_i[801];
  assign N3027 = N3024 | N3026;
  assign N3030 = ~sel_i[803];
  assign N3032 = N3029 | N3031;
  assign N3035 = ~sel_i[805];
  assign N3037 = N3034 | N3036;
  assign N3040 = ~sel_i[807];
  assign N3042 = N3039 | N3041;
  assign N3045 = ~sel_i[809];
  assign N3047 = N3044 | N3046;
  assign N3050 = ~sel_i[811];
  assign N3052 = N3049 | N3051;
  assign N3055 = ~sel_i[813];
  assign N3057 = N3054 | N3056;
  assign N3060 = ~sel_i[815];
  assign N3062 = N3059 | N3061;
  assign N3065 = ~sel_i[817];
  assign N3067 = N3064 | N3066;
  assign N3070 = ~sel_i[819];
  assign N3072 = N3069 | N3071;
  assign N3075 = ~sel_i[821];
  assign N3077 = N3074 | N3076;
  assign N3080 = ~sel_i[823];
  assign N3082 = N3079 | N3081;
  assign N3085 = ~sel_i[825];
  assign N3087 = N3084 | N3086;
  assign N3090 = ~sel_i[827];
  assign N3092 = N3089 | N3091;
  assign N3095 = ~sel_i[829];
  assign N3097 = N3094 | N3096;
  assign N3100 = ~sel_i[831];
  assign N3102 = N3099 | N3101;
  assign N3105 = ~sel_i[833];
  assign N3107 = N3104 | N3106;
  assign N3110 = ~sel_i[835];
  assign N3112 = N3109 | N3111;
  assign N3115 = ~sel_i[837];
  assign N3117 = N3114 | N3116;
  assign N3120 = ~sel_i[839];
  assign N3122 = N3119 | N3121;
  assign N3125 = ~sel_i[841];
  assign N3127 = N3124 | N3126;
  assign N3130 = ~sel_i[843];
  assign N3132 = N3129 | N3131;
  assign N3135 = ~sel_i[845];
  assign N3137 = N3134 | N3136;
  assign N3140 = ~sel_i[847];
  assign N3142 = N3139 | N3141;
  assign N3145 = ~sel_i[849];
  assign N3147 = N3144 | N3146;
  assign N3150 = ~sel_i[851];
  assign N3152 = N3149 | N3151;
  assign N3155 = ~sel_i[853];
  assign N3157 = N3154 | N3156;
  assign N3160 = ~sel_i[855];
  assign N3162 = N3159 | N3161;
  assign N3165 = ~sel_i[857];
  assign N3167 = N3164 | N3166;
  assign N3170 = ~sel_i[859];
  assign N3172 = N3169 | N3171;
  assign N3175 = ~sel_i[861];
  assign N3177 = N3174 | N3176;
  assign N3180 = ~sel_i[863];
  assign N3182 = N3179 | N3181;
  assign N3185 = ~sel_i[865];
  assign N3187 = N3184 | N3186;
  assign N3190 = ~sel_i[867];
  assign N3192 = N3189 | N3191;
  assign N3195 = ~sel_i[869];
  assign N3197 = N3194 | N3196;
  assign N3200 = ~sel_i[871];
  assign N3202 = N3199 | N3201;
  assign N3205 = ~sel_i[873];
  assign N3207 = N3204 | N3206;
  assign N3210 = ~sel_i[875];
  assign N3212 = N3209 | N3211;
  assign N3215 = ~sel_i[877];
  assign N3217 = N3214 | N3216;
  assign N3220 = ~sel_i[879];
  assign N3222 = N3219 | N3221;
  assign N3225 = ~sel_i[881];
  assign N3227 = N3224 | N3226;
  assign N3230 = ~sel_i[883];
  assign N3232 = N3229 | N3231;
  assign N3235 = ~sel_i[885];
  assign N3237 = N3234 | N3236;
  assign N3240 = ~sel_i[887];
  assign N3242 = N3239 | N3241;
  assign N3245 = ~sel_i[889];
  assign N3247 = N3244 | N3246;
  assign N3250 = ~sel_i[891];
  assign N3252 = N3249 | N3251;
  assign N3255 = ~sel_i[893];
  assign N3257 = N3254 | N3256;
  assign N3260 = ~sel_i[895];
  assign N3262 = N3259 | N3261;
  assign N3265 = ~sel_i[897];
  assign N3267 = N3264 | N3266;
  assign N3270 = ~sel_i[899];
  assign N3272 = N3269 | N3271;
  assign N3275 = ~sel_i[901];
  assign N3277 = N3274 | N3276;
  assign N3280 = ~sel_i[903];
  assign N3282 = N3279 | N3281;
  assign N3285 = ~sel_i[905];
  assign N3287 = N3284 | N3286;
  assign N3290 = ~sel_i[907];
  assign N3292 = N3289 | N3291;
  assign N3295 = ~sel_i[909];
  assign N3297 = N3294 | N3296;
  assign N3300 = ~sel_i[911];
  assign N3302 = N3299 | N3301;
  assign N3305 = ~sel_i[913];
  assign N3307 = N3304 | N3306;
  assign N3310 = ~sel_i[915];
  assign N3312 = N3309 | N3311;
  assign N3315 = ~sel_i[917];
  assign N3317 = N3314 | N3316;
  assign N3320 = ~sel_i[919];
  assign N3322 = N3319 | N3321;
  assign N3325 = ~sel_i[921];
  assign N3327 = N3324 | N3326;
  assign N3330 = ~sel_i[923];
  assign N3332 = N3329 | N3331;
  assign N3335 = ~sel_i[925];
  assign N3337 = N3334 | N3336;
  assign N3340 = ~sel_i[927];
  assign N3342 = N3339 | N3341;
  assign N3345 = ~sel_i[929];
  assign N3347 = N3344 | N3346;
  assign N3350 = ~sel_i[931];
  assign N3352 = N3349 | N3351;
  assign N3355 = ~sel_i[933];
  assign N3357 = N3354 | N3356;
  assign N3360 = ~sel_i[935];
  assign N3362 = N3359 | N3361;
  assign N3365 = ~sel_i[937];
  assign N3367 = N3364 | N3366;
  assign N3370 = ~sel_i[939];
  assign N3372 = N3369 | N3371;
  assign N3375 = ~sel_i[941];
  assign N3377 = N3374 | N3376;
  assign N3380 = ~sel_i[943];
  assign N3382 = N3379 | N3381;
  assign N3385 = ~sel_i[945];
  assign N3387 = N3384 | N3386;
  assign N3390 = ~sel_i[947];
  assign N3392 = N3389 | N3391;
  assign N3395 = ~sel_i[949];
  assign N3397 = N3394 | N3396;
  assign N3400 = ~sel_i[951];
  assign N3402 = N3399 | N3401;
  assign N3405 = ~sel_i[953];
  assign N3407 = N3404 | N3406;
  assign N3410 = ~sel_i[955];
  assign N3412 = N3409 | N3411;
  assign N3415 = ~sel_i[957];
  assign N3417 = N3414 | N3416;
  assign N3420 = ~sel_i[959];
  assign N3422 = N3419 | N3421;
  assign N3425 = ~sel_i[961];
  assign N3427 = N3424 | N3426;
  assign N3430 = ~sel_i[963];
  assign N3432 = N3429 | N3431;
  assign N3435 = ~sel_i[965];
  assign N3437 = N3434 | N3436;
  assign N3440 = ~sel_i[967];
  assign N3442 = N3439 | N3441;
  assign N3445 = ~sel_i[969];
  assign N3447 = N3444 | N3446;
  assign N3450 = ~sel_i[971];
  assign N3452 = N3449 | N3451;
  assign N3455 = ~sel_i[973];
  assign N3457 = N3454 | N3456;
  assign N3460 = ~sel_i[975];
  assign N3462 = N3459 | N3461;
  assign N3465 = ~sel_i[977];
  assign N3467 = N3464 | N3466;
  assign N3470 = ~sel_i[979];
  assign N3472 = N3469 | N3471;
  assign N3475 = ~sel_i[981];
  assign N3477 = N3474 | N3476;
  assign N3480 = ~sel_i[983];
  assign N3482 = N3479 | N3481;
  assign N3485 = ~sel_i[985];
  assign N3487 = N3484 | N3486;
  assign N3490 = ~sel_i[987];
  assign N3492 = N3489 | N3491;
  assign N3495 = ~sel_i[989];
  assign N3497 = N3494 | N3496;
  assign N3500 = ~sel_i[991];
  assign N3502 = N3499 | N3501;
  assign N3505 = ~sel_i[993];
  assign N3507 = N3504 | N3506;
  assign N3510 = ~sel_i[995];
  assign N3512 = N3509 | N3511;
  assign N3515 = ~sel_i[997];
  assign N3517 = N3514 | N3516;
  assign N3520 = ~sel_i[999];
  assign N3522 = N3519 | N3521;
  assign N3525 = ~sel_i[1001];
  assign N3527 = N3524 | N3526;
  assign N3530 = ~sel_i[1003];
  assign N3532 = N3529 | N3531;
  assign N3535 = ~sel_i[1005];
  assign N3537 = N3534 | N3536;
  assign N3540 = ~sel_i[1007];
  assign N3542 = N3539 | N3541;
  assign N3545 = ~sel_i[1009];
  assign N3547 = N3544 | N3546;
  assign N3550 = ~sel_i[1011];
  assign N3552 = N3549 | N3551;
  assign N3555 = ~sel_i[1013];
  assign N3557 = N3554 | N3556;
  assign N3560 = ~sel_i[1015];
  assign N3562 = N3559 | N3561;
  assign N3565 = ~sel_i[1017];
  assign N3567 = N3564 | N3566;
  assign N3570 = ~sel_i[1019];
  assign N3572 = N3569 | N3571;
  assign N3575 = ~sel_i[1021];
  assign N3577 = N3574 | N3576;
  assign N3580 = ~sel_i[1023];
  assign N3582 = N3579 | N3581;
  assign N3584 = ~N1027;
  assign N3585 = ~N1032;
  assign N3586 = ~N1037;
  assign N3587 = ~N1042;
  assign N3588 = ~N1047;
  assign N3589 = ~N1052;
  assign N3590 = ~N1057;
  assign N3591 = ~N1062;
  assign N3592 = ~N1067;
  assign N3593 = ~N1072;
  assign N3594 = ~N1077;
  assign N3595 = ~N1082;
  assign N3596 = ~N1087;
  assign N3597 = ~N1092;
  assign N3598 = ~N1097;
  assign N3599 = ~N1102;
  assign N3600 = ~N1107;
  assign N3601 = ~N1112;
  assign N3602 = ~N1117;
  assign N3603 = ~N1122;
  assign N3604 = ~N1127;
  assign N3605 = ~N1132;
  assign N3606 = ~N1137;
  assign N3607 = ~N1142;
  assign N3608 = ~N1147;
  assign N3609 = ~N1152;
  assign N3610 = ~N1157;
  assign N3611 = ~N1162;
  assign N3612 = ~N1167;
  assign N3613 = ~N1172;
  assign N3614 = ~N1177;
  assign N3615 = ~N1182;
  assign N3616 = ~N1187;
  assign N3617 = ~N1192;
  assign N3618 = ~N1197;
  assign N3619 = ~N1202;
  assign N3620 = ~N1207;
  assign N3621 = ~N1212;
  assign N3622 = ~N1217;
  assign N3623 = ~N1222;
  assign N3624 = ~N1227;
  assign N3625 = ~N1232;
  assign N3626 = ~N1237;
  assign N3627 = ~N1242;
  assign N3628 = ~N1247;
  assign N3629 = ~N1252;
  assign N3630 = ~N1257;
  assign N3631 = ~N1262;
  assign N3632 = ~N1267;
  assign N3633 = ~N1272;
  assign N3634 = ~N1277;
  assign N3635 = ~N1282;
  assign N3636 = ~N1287;
  assign N3637 = ~N1292;
  assign N3638 = ~N1297;
  assign N3639 = ~N1302;
  assign N3640 = ~N1307;
  assign N3641 = ~N1312;
  assign N3642 = ~N1317;
  assign N3643 = ~N1322;
  assign N3644 = ~N1327;
  assign N3645 = ~N1332;
  assign N3646 = ~N1337;
  assign N3647 = ~N1342;
  assign N3648 = ~N1347;
  assign N3649 = ~N1352;
  assign N3650 = ~N1357;
  assign N3651 = ~N1362;
  assign N3652 = ~N1367;
  assign N3653 = ~N1372;
  assign N3654 = ~N1377;
  assign N3655 = ~N1382;
  assign N3656 = ~N1387;
  assign N3657 = ~N1392;
  assign N3658 = ~N1397;
  assign N3659 = ~N1402;
  assign N3660 = ~N1407;
  assign N3661 = ~N1412;
  assign N3662 = ~N1417;
  assign N3663 = ~N1422;
  assign N3664 = ~N1427;
  assign N3665 = ~N1432;
  assign N3666 = ~N1437;
  assign N3667 = ~N1442;
  assign N3668 = ~N1447;
  assign N3669 = ~N1452;
  assign N3670 = ~N1457;
  assign N3671 = ~N1462;
  assign N3672 = ~N1467;
  assign N3673 = ~N1472;
  assign N3674 = ~N1477;
  assign N3675 = ~N1482;
  assign N3676 = ~N1487;
  assign N3677 = ~N1492;
  assign N3678 = ~N1497;
  assign N3679 = ~N1502;
  assign N3680 = ~N1507;
  assign N3681 = ~N1512;
  assign N3682 = ~N1517;
  assign N3683 = ~N1522;
  assign N3684 = ~N1527;
  assign N3685 = ~N1532;
  assign N3686 = ~N1537;
  assign N3687 = ~N1542;
  assign N3688 = ~N1547;
  assign N3689 = ~N1552;
  assign N3690 = ~N1557;
  assign N3691 = ~N1562;
  assign N3692 = ~N1567;
  assign N3693 = ~N1572;
  assign N3694 = ~N1577;
  assign N3695 = ~N1582;
  assign N3696 = ~N1587;
  assign N3697 = ~N1592;
  assign N3698 = ~N1597;
  assign N3699 = ~N1602;
  assign N3700 = ~N1607;
  assign N3701 = ~N1612;
  assign N3702 = ~N1617;
  assign N3703 = ~N1622;
  assign N3704 = ~N1627;
  assign N3705 = ~N1632;
  assign N3706 = ~N1637;
  assign N3707 = ~N1642;
  assign N3708 = ~N1647;
  assign N3709 = ~N1652;
  assign N3710 = ~N1657;
  assign N3711 = ~N1662;
  assign N3712 = ~N1667;
  assign N3713 = ~N1672;
  assign N3714 = ~N1677;
  assign N3715 = ~N1682;
  assign N3716 = ~N1687;
  assign N3717 = ~N1692;
  assign N3718 = ~N1697;
  assign N3719 = ~N1702;
  assign N3720 = ~N1707;
  assign N3721 = ~N1712;
  assign N3722 = ~N1717;
  assign N3723 = ~N1722;
  assign N3724 = ~N1727;
  assign N3725 = ~N1732;
  assign N3726 = ~N1737;
  assign N3727 = ~N1742;
  assign N3728 = ~N1747;
  assign N3729 = ~N1752;
  assign N3730 = ~N1757;
  assign N3731 = ~N1762;
  assign N3732 = ~N1767;
  assign N3733 = ~N1772;
  assign N3734 = ~N1777;
  assign N3735 = ~N1782;
  assign N3736 = ~N1787;
  assign N3737 = ~N1792;
  assign N3738 = ~N1797;
  assign N3739 = ~N1802;
  assign N3740 = ~N1807;
  assign N3741 = ~N1812;
  assign N3742 = ~N1817;
  assign N3743 = ~N1822;
  assign N3744 = ~N1827;
  assign N3745 = ~N1832;
  assign N3746 = ~N1837;
  assign N3747 = ~N1842;
  assign N3748 = ~N1847;
  assign N3749 = ~N1852;
  assign N3750 = ~N1857;
  assign N3751 = ~N1862;
  assign N3752 = ~N1867;
  assign N3753 = ~N1872;
  assign N3754 = ~N1877;
  assign N3755 = ~N1882;
  assign N3756 = ~N1887;
  assign N3757 = ~N1892;
  assign N3758 = ~N1897;
  assign N3759 = ~N1902;
  assign N3760 = ~N1907;
  assign N3761 = ~N1912;
  assign N3762 = ~N1917;
  assign N3763 = ~N1922;
  assign N3764 = ~N1927;
  assign N3765 = ~N1932;
  assign N3766 = ~N1937;
  assign N3767 = ~N1942;
  assign N3768 = ~N1947;
  assign N3769 = ~N1952;
  assign N3770 = ~N1957;
  assign N3771 = ~N1962;
  assign N3772 = ~N1967;
  assign N3773 = ~N1972;
  assign N3774 = ~N1977;
  assign N3775 = ~N1982;
  assign N3776 = ~N1987;
  assign N3777 = ~N1992;
  assign N3778 = ~N1997;
  assign N3779 = ~N2002;
  assign N3780 = ~N2007;
  assign N3781 = ~N2012;
  assign N3782 = ~N2017;
  assign N3783 = ~N2022;
  assign N3784 = ~N2027;
  assign N3785 = ~N2032;
  assign N3786 = ~N2037;
  assign N3787 = ~N2042;
  assign N3788 = ~N2047;
  assign N3789 = ~N2052;
  assign N3790 = ~N2057;
  assign N3791 = ~N2062;
  assign N3792 = ~N2067;
  assign N3793 = ~N2072;
  assign N3794 = ~N2077;
  assign N3795 = ~N2082;
  assign N3796 = ~N2087;
  assign N3797 = ~N2092;
  assign N3798 = ~N2097;
  assign N3799 = ~N2102;
  assign N3800 = ~N2107;
  assign N3801 = ~N2112;
  assign N3802 = ~N2117;
  assign N3803 = ~N2122;
  assign N3804 = ~N2127;
  assign N3805 = ~N2132;
  assign N3806 = ~N2137;
  assign N3807 = ~N2142;
  assign N3808 = ~N2147;
  assign N3809 = ~N2152;
  assign N3810 = ~N2157;
  assign N3811 = ~N2162;
  assign N3812 = ~N2167;
  assign N3813 = ~N2172;
  assign N3814 = ~N2177;
  assign N3815 = ~N2182;
  assign N3816 = ~N2187;
  assign N3817 = ~N2192;
  assign N3818 = ~N2197;
  assign N3819 = ~N2202;
  assign N3820 = ~N2207;
  assign N3821 = ~N2212;
  assign N3822 = ~N2217;
  assign N3823 = ~N2222;
  assign N3824 = ~N2227;
  assign N3825 = ~N2232;
  assign N3826 = ~N2237;
  assign N3827 = ~N2242;
  assign N3828 = ~N2247;
  assign N3829 = ~N2252;
  assign N3830 = ~N2257;
  assign N3831 = ~N2262;
  assign N3832 = ~N2267;
  assign N3833 = ~N2272;
  assign N3834 = ~N2277;
  assign N3835 = ~N2282;
  assign N3836 = ~N2287;
  assign N3837 = ~N2292;
  assign N3838 = ~N2297;
  assign N3839 = ~N2302;
  assign N3840 = ~N2307;
  assign N3841 = ~N2312;
  assign N3842 = ~N2317;
  assign N3843 = ~N2322;
  assign N3844 = ~N2327;
  assign N3845 = ~N2332;
  assign N3846 = ~N2337;
  assign N3847 = ~N2342;
  assign N3848 = ~N2347;
  assign N3849 = ~N2352;
  assign N3850 = ~N2357;
  assign N3851 = ~N2362;
  assign N3852 = ~N2367;
  assign N3853 = ~N2372;
  assign N3854 = ~N2377;
  assign N3855 = ~N2382;
  assign N3856 = ~N2387;
  assign N3857 = ~N2392;
  assign N3858 = ~N2397;
  assign N3859 = ~N2402;
  assign N3860 = ~N2407;
  assign N3861 = ~N2412;
  assign N3862 = ~N2417;
  assign N3863 = ~N2422;
  assign N3864 = ~N2427;
  assign N3865 = ~N2432;
  assign N3866 = ~N2437;
  assign N3867 = ~N2442;
  assign N3868 = ~N2447;
  assign N3869 = ~N2452;
  assign N3870 = ~N2457;
  assign N3871 = ~N2462;
  assign N3872 = ~N2467;
  assign N3873 = ~N2472;
  assign N3874 = ~N2477;
  assign N3875 = ~N2482;
  assign N3876 = ~N2487;
  assign N3877 = ~N2492;
  assign N3878 = ~N2497;
  assign N3879 = ~N2502;
  assign N3880 = ~N2507;
  assign N3881 = ~N2512;
  assign N3882 = ~N2517;
  assign N3883 = ~N2522;
  assign N3884 = ~N2527;
  assign N3885 = ~N2532;
  assign N3886 = ~N2537;
  assign N3887 = ~N2542;
  assign N3888 = ~N2547;
  assign N3889 = ~N2552;
  assign N3890 = ~N2557;
  assign N3891 = ~N2562;
  assign N3892 = ~N2567;
  assign N3893 = ~N2572;
  assign N3894 = ~N2577;
  assign N3895 = ~N2582;
  assign N3896 = ~N2587;
  assign N3897 = ~N2592;
  assign N3898 = ~N2597;
  assign N3899 = ~N2602;
  assign N3900 = ~N2607;
  assign N3901 = ~N2612;
  assign N3902 = ~N2617;
  assign N3903 = ~N2622;
  assign N3904 = ~N2627;
  assign N3905 = ~N2632;
  assign N3906 = ~N2637;
  assign N3907 = ~N2642;
  assign N3908 = ~N2647;
  assign N3909 = ~N2652;
  assign N3910 = ~N2657;
  assign N3911 = ~N2662;
  assign N3912 = ~N2667;
  assign N3913 = ~N2672;
  assign N3914 = ~N2677;
  assign N3915 = ~N2682;
  assign N3916 = ~N2687;
  assign N3917 = ~N2692;
  assign N3918 = ~N2697;
  assign N3919 = ~N2702;
  assign N3920 = ~N2707;
  assign N3921 = ~N2712;
  assign N3922 = ~N2717;
  assign N3923 = ~N2722;
  assign N3924 = ~N2727;
  assign N3925 = ~N2732;
  assign N3926 = ~N2737;
  assign N3927 = ~N2742;
  assign N3928 = ~N2747;
  assign N3929 = ~N2752;
  assign N3930 = ~N2757;
  assign N3931 = ~N2762;
  assign N3932 = ~N2767;
  assign N3933 = ~N2772;
  assign N3934 = ~N2777;
  assign N3935 = ~N2782;
  assign N3936 = ~N2787;
  assign N3937 = ~N2792;
  assign N3938 = ~N2797;
  assign N3939 = ~N2802;
  assign N3940 = ~N2807;
  assign N3941 = ~N2812;
  assign N3942 = ~N2817;
  assign N3943 = ~N2822;
  assign N3944 = ~N2827;
  assign N3945 = ~N2832;
  assign N3946 = ~N2837;
  assign N3947 = ~N2842;
  assign N3948 = ~N2847;
  assign N3949 = ~N2852;
  assign N3950 = ~N2857;
  assign N3951 = ~N2862;
  assign N3952 = ~N2867;
  assign N3953 = ~N2872;
  assign N3954 = ~N2877;
  assign N3955 = ~N2882;
  assign N3956 = ~N2887;
  assign N3957 = ~N2892;
  assign N3958 = ~N2897;
  assign N3959 = ~N2902;
  assign N3960 = ~N2907;
  assign N3961 = ~N2912;
  assign N3962 = ~N2917;
  assign N3963 = ~N2922;
  assign N3964 = ~N2927;
  assign N3965 = ~N2932;
  assign N3966 = ~N2937;
  assign N3967 = ~N2942;
  assign N3968 = ~N2947;
  assign N3969 = ~N2952;
  assign N3970 = ~N2957;
  assign N3971 = ~N2962;
  assign N3972 = ~N2967;
  assign N3973 = ~N2972;
  assign N3974 = ~N2977;
  assign N3975 = ~N2982;
  assign N3976 = ~N2987;
  assign N3977 = ~N2992;
  assign N3978 = ~N2997;
  assign N3979 = ~N3002;
  assign N3980 = ~N3007;
  assign N3981 = ~N3012;
  assign N3982 = ~N3017;
  assign N3983 = ~N3022;
  assign N3984 = ~N3027;
  assign N3985 = ~N3032;
  assign N3986 = ~N3037;
  assign N3987 = ~N3042;
  assign N3988 = ~N3047;
  assign N3989 = ~N3052;
  assign N3990 = ~N3057;
  assign N3991 = ~N3062;
  assign N3992 = ~N3067;
  assign N3993 = ~N3072;
  assign N3994 = ~N3077;
  assign N3995 = ~N3082;
  assign N3996 = ~N3087;
  assign N3997 = ~N3092;
  assign N3998 = ~N3097;
  assign N3999 = ~N3102;
  assign N4000 = ~N3107;
  assign N4001 = ~N3112;
  assign N4002 = ~N3117;
  assign N4003 = ~N3122;
  assign N4004 = ~N3127;
  assign N4005 = ~N3132;
  assign N4006 = ~N3137;
  assign N4007 = ~N3142;
  assign N4008 = ~N3147;
  assign N4009 = ~N3152;
  assign N4010 = ~N3157;
  assign N4011 = ~N3162;
  assign N4012 = ~N3167;
  assign N4013 = ~N3172;
  assign N4014 = ~N3177;
  assign N4015 = ~N3182;
  assign N4016 = ~N3187;
  assign N4017 = ~N3192;
  assign N4018 = ~N3197;
  assign N4019 = ~N3202;
  assign N4020 = ~N3207;
  assign N4021 = ~N3212;
  assign N4022 = ~N3217;
  assign N4023 = ~N3222;
  assign N4024 = ~N3227;
  assign N4025 = ~N3232;
  assign N4026 = ~N3237;
  assign N4027 = ~N3242;
  assign N4028 = ~N3247;
  assign N4029 = ~N3252;
  assign N4030 = ~N3257;
  assign N4031 = ~N3262;
  assign N4032 = ~N3267;
  assign N4033 = ~N3272;
  assign N4034 = ~N3277;
  assign N4035 = ~N3282;
  assign N4036 = ~N3287;
  assign N4037 = ~N3292;
  assign N4038 = ~N3297;
  assign N4039 = ~N3302;
  assign N4040 = ~N3307;
  assign N4041 = ~N3312;
  assign N4042 = ~N3317;
  assign N4043 = ~N3322;
  assign N4044 = ~N3327;
  assign N4045 = ~N3332;
  assign N4046 = ~N3337;
  assign N4047 = ~N3342;
  assign N4048 = ~N3347;
  assign N4049 = ~N3352;
  assign N4050 = ~N3357;
  assign N4051 = ~N3362;
  assign N4052 = ~N3367;
  assign N4053 = ~N3372;
  assign N4054 = ~N3377;
  assign N4055 = ~N3382;
  assign N4056 = ~N3387;
  assign N4057 = ~N3392;
  assign N4058 = ~N3397;
  assign N4059 = ~N3402;
  assign N4060 = ~N3407;
  assign N4061 = ~N3412;
  assign N4062 = ~N3417;
  assign N4063 = ~N3422;
  assign N4064 = ~N3427;
  assign N4065 = ~N3432;
  assign N4066 = ~N3437;
  assign N4067 = ~N3442;
  assign N4068 = ~N3447;
  assign N4069 = ~N3452;
  assign N4070 = ~N3457;
  assign N4071 = ~N3462;
  assign N4072 = ~N3467;
  assign N4073 = ~N3472;
  assign N4074 = ~N3477;
  assign N4075 = ~N3482;
  assign N4076 = ~N3487;
  assign N4077 = ~N3492;
  assign N4078 = ~N3497;
  assign N4079 = ~N3502;
  assign N4080 = ~N3507;
  assign N4081 = ~N3512;
  assign N4082 = ~N3517;
  assign N4083 = ~N3522;
  assign N4084 = ~N3527;
  assign N4085 = ~N3532;
  assign N4086 = ~N3537;
  assign N4087 = ~N3542;
  assign N4088 = ~N3547;
  assign N4089 = ~N3552;
  assign N4090 = ~N3557;
  assign N4091 = ~N3562;
  assign N4092 = ~N3567;
  assign N4093 = ~N3572;
  assign N4094 = ~N3577;
  assign N4095 = ~N3582;

  always @(posedge clk_i) begin
    if(N3584) begin
      { data_o[63:0] } <= { r_n_0__63_, r_n_0__62_, r_n_0__61_, r_n_0__60_, r_n_0__59_, r_n_0__58_, r_n_0__57_, r_n_0__56_, r_n_0__55_, r_n_0__54_, r_n_0__53_, r_n_0__52_, r_n_0__51_, r_n_0__50_, r_n_0__49_, r_n_0__48_, r_n_0__47_, r_n_0__46_, r_n_0__45_, r_n_0__44_, r_n_0__43_, r_n_0__42_, r_n_0__41_, r_n_0__40_, r_n_0__39_, r_n_0__38_, r_n_0__37_, r_n_0__36_, r_n_0__35_, r_n_0__34_, r_n_0__33_, r_n_0__32_, r_n_0__31_, r_n_0__30_, r_n_0__29_, r_n_0__28_, r_n_0__27_, r_n_0__26_, r_n_0__25_, r_n_0__24_, r_n_0__23_, r_n_0__22_, r_n_0__21_, r_n_0__20_, r_n_0__19_, r_n_0__18_, r_n_0__17_, r_n_0__16_, r_n_0__15_, r_n_0__14_, r_n_0__13_, r_n_0__12_, r_n_0__11_, r_n_0__10_, r_n_0__9_, r_n_0__8_, r_n_0__7_, r_n_0__6_, r_n_0__5_, r_n_0__4_, r_n_0__3_, r_n_0__2_, r_n_0__1_, r_n_0__0_ };
    end 
    if(N3585) begin
      r_1__63_ <= r_n_1__63_;
      r_1__62_ <= r_n_1__62_;
      r_1__61_ <= r_n_1__61_;
      r_1__60_ <= r_n_1__60_;
      r_1__59_ <= r_n_1__59_;
      r_1__58_ <= r_n_1__58_;
      r_1__57_ <= r_n_1__57_;
      r_1__56_ <= r_n_1__56_;
      r_1__55_ <= r_n_1__55_;
      r_1__54_ <= r_n_1__54_;
      r_1__53_ <= r_n_1__53_;
      r_1__52_ <= r_n_1__52_;
      r_1__51_ <= r_n_1__51_;
      r_1__50_ <= r_n_1__50_;
      r_1__49_ <= r_n_1__49_;
      r_1__48_ <= r_n_1__48_;
      r_1__47_ <= r_n_1__47_;
      r_1__46_ <= r_n_1__46_;
      r_1__45_ <= r_n_1__45_;
      r_1__44_ <= r_n_1__44_;
      r_1__43_ <= r_n_1__43_;
      r_1__42_ <= r_n_1__42_;
      r_1__41_ <= r_n_1__41_;
      r_1__40_ <= r_n_1__40_;
      r_1__39_ <= r_n_1__39_;
      r_1__38_ <= r_n_1__38_;
      r_1__37_ <= r_n_1__37_;
      r_1__36_ <= r_n_1__36_;
      r_1__35_ <= r_n_1__35_;
      r_1__34_ <= r_n_1__34_;
      r_1__33_ <= r_n_1__33_;
      r_1__32_ <= r_n_1__32_;
      r_1__31_ <= r_n_1__31_;
      r_1__30_ <= r_n_1__30_;
      r_1__29_ <= r_n_1__29_;
      r_1__28_ <= r_n_1__28_;
      r_1__27_ <= r_n_1__27_;
      r_1__26_ <= r_n_1__26_;
      r_1__25_ <= r_n_1__25_;
      r_1__24_ <= r_n_1__24_;
      r_1__23_ <= r_n_1__23_;
      r_1__22_ <= r_n_1__22_;
      r_1__21_ <= r_n_1__21_;
      r_1__20_ <= r_n_1__20_;
      r_1__19_ <= r_n_1__19_;
      r_1__18_ <= r_n_1__18_;
      r_1__17_ <= r_n_1__17_;
      r_1__16_ <= r_n_1__16_;
      r_1__15_ <= r_n_1__15_;
      r_1__14_ <= r_n_1__14_;
      r_1__13_ <= r_n_1__13_;
      r_1__12_ <= r_n_1__12_;
      r_1__11_ <= r_n_1__11_;
      r_1__10_ <= r_n_1__10_;
      r_1__9_ <= r_n_1__9_;
      r_1__8_ <= r_n_1__8_;
      r_1__7_ <= r_n_1__7_;
      r_1__6_ <= r_n_1__6_;
      r_1__5_ <= r_n_1__5_;
      r_1__4_ <= r_n_1__4_;
      r_1__3_ <= r_n_1__3_;
      r_1__2_ <= r_n_1__2_;
      r_1__1_ <= r_n_1__1_;
      r_1__0_ <= r_n_1__0_;
    end 
    if(N3586) begin
      r_2__63_ <= r_n_2__63_;
      r_2__62_ <= r_n_2__62_;
      r_2__61_ <= r_n_2__61_;
      r_2__60_ <= r_n_2__60_;
      r_2__59_ <= r_n_2__59_;
      r_2__58_ <= r_n_2__58_;
      r_2__57_ <= r_n_2__57_;
      r_2__56_ <= r_n_2__56_;
      r_2__55_ <= r_n_2__55_;
      r_2__54_ <= r_n_2__54_;
      r_2__53_ <= r_n_2__53_;
      r_2__52_ <= r_n_2__52_;
      r_2__51_ <= r_n_2__51_;
      r_2__50_ <= r_n_2__50_;
      r_2__49_ <= r_n_2__49_;
      r_2__48_ <= r_n_2__48_;
      r_2__47_ <= r_n_2__47_;
      r_2__46_ <= r_n_2__46_;
      r_2__45_ <= r_n_2__45_;
      r_2__44_ <= r_n_2__44_;
      r_2__43_ <= r_n_2__43_;
      r_2__42_ <= r_n_2__42_;
      r_2__41_ <= r_n_2__41_;
      r_2__40_ <= r_n_2__40_;
      r_2__39_ <= r_n_2__39_;
      r_2__38_ <= r_n_2__38_;
      r_2__37_ <= r_n_2__37_;
      r_2__36_ <= r_n_2__36_;
      r_2__35_ <= r_n_2__35_;
      r_2__34_ <= r_n_2__34_;
      r_2__33_ <= r_n_2__33_;
      r_2__32_ <= r_n_2__32_;
      r_2__31_ <= r_n_2__31_;
      r_2__30_ <= r_n_2__30_;
      r_2__29_ <= r_n_2__29_;
      r_2__28_ <= r_n_2__28_;
      r_2__27_ <= r_n_2__27_;
      r_2__26_ <= r_n_2__26_;
      r_2__25_ <= r_n_2__25_;
      r_2__24_ <= r_n_2__24_;
      r_2__23_ <= r_n_2__23_;
      r_2__22_ <= r_n_2__22_;
      r_2__21_ <= r_n_2__21_;
      r_2__20_ <= r_n_2__20_;
      r_2__19_ <= r_n_2__19_;
      r_2__18_ <= r_n_2__18_;
      r_2__17_ <= r_n_2__17_;
      r_2__16_ <= r_n_2__16_;
      r_2__15_ <= r_n_2__15_;
      r_2__14_ <= r_n_2__14_;
      r_2__13_ <= r_n_2__13_;
      r_2__12_ <= r_n_2__12_;
      r_2__11_ <= r_n_2__11_;
      r_2__10_ <= r_n_2__10_;
      r_2__9_ <= r_n_2__9_;
      r_2__8_ <= r_n_2__8_;
      r_2__7_ <= r_n_2__7_;
      r_2__6_ <= r_n_2__6_;
      r_2__5_ <= r_n_2__5_;
      r_2__4_ <= r_n_2__4_;
      r_2__3_ <= r_n_2__3_;
      r_2__2_ <= r_n_2__2_;
      r_2__1_ <= r_n_2__1_;
      r_2__0_ <= r_n_2__0_;
    end 
    if(N3587) begin
      r_3__63_ <= r_n_3__63_;
      r_3__62_ <= r_n_3__62_;
      r_3__61_ <= r_n_3__61_;
      r_3__60_ <= r_n_3__60_;
      r_3__59_ <= r_n_3__59_;
      r_3__58_ <= r_n_3__58_;
      r_3__57_ <= r_n_3__57_;
      r_3__56_ <= r_n_3__56_;
      r_3__55_ <= r_n_3__55_;
      r_3__54_ <= r_n_3__54_;
      r_3__53_ <= r_n_3__53_;
      r_3__52_ <= r_n_3__52_;
      r_3__51_ <= r_n_3__51_;
      r_3__50_ <= r_n_3__50_;
      r_3__49_ <= r_n_3__49_;
      r_3__48_ <= r_n_3__48_;
      r_3__47_ <= r_n_3__47_;
      r_3__46_ <= r_n_3__46_;
      r_3__45_ <= r_n_3__45_;
      r_3__44_ <= r_n_3__44_;
      r_3__43_ <= r_n_3__43_;
      r_3__42_ <= r_n_3__42_;
      r_3__41_ <= r_n_3__41_;
      r_3__40_ <= r_n_3__40_;
      r_3__39_ <= r_n_3__39_;
      r_3__38_ <= r_n_3__38_;
      r_3__37_ <= r_n_3__37_;
      r_3__36_ <= r_n_3__36_;
      r_3__35_ <= r_n_3__35_;
      r_3__34_ <= r_n_3__34_;
      r_3__33_ <= r_n_3__33_;
      r_3__32_ <= r_n_3__32_;
      r_3__31_ <= r_n_3__31_;
      r_3__30_ <= r_n_3__30_;
      r_3__29_ <= r_n_3__29_;
      r_3__28_ <= r_n_3__28_;
      r_3__27_ <= r_n_3__27_;
      r_3__26_ <= r_n_3__26_;
      r_3__25_ <= r_n_3__25_;
      r_3__24_ <= r_n_3__24_;
      r_3__23_ <= r_n_3__23_;
      r_3__22_ <= r_n_3__22_;
      r_3__21_ <= r_n_3__21_;
      r_3__20_ <= r_n_3__20_;
      r_3__19_ <= r_n_3__19_;
      r_3__18_ <= r_n_3__18_;
      r_3__17_ <= r_n_3__17_;
      r_3__16_ <= r_n_3__16_;
      r_3__15_ <= r_n_3__15_;
      r_3__14_ <= r_n_3__14_;
      r_3__13_ <= r_n_3__13_;
      r_3__12_ <= r_n_3__12_;
      r_3__11_ <= r_n_3__11_;
      r_3__10_ <= r_n_3__10_;
      r_3__9_ <= r_n_3__9_;
      r_3__8_ <= r_n_3__8_;
      r_3__7_ <= r_n_3__7_;
      r_3__6_ <= r_n_3__6_;
      r_3__5_ <= r_n_3__5_;
      r_3__4_ <= r_n_3__4_;
      r_3__3_ <= r_n_3__3_;
      r_3__2_ <= r_n_3__2_;
      r_3__1_ <= r_n_3__1_;
      r_3__0_ <= r_n_3__0_;
    end 
    if(N3588) begin
      r_4__63_ <= r_n_4__63_;
      r_4__62_ <= r_n_4__62_;
      r_4__61_ <= r_n_4__61_;
      r_4__60_ <= r_n_4__60_;
      r_4__59_ <= r_n_4__59_;
      r_4__58_ <= r_n_4__58_;
      r_4__57_ <= r_n_4__57_;
      r_4__56_ <= r_n_4__56_;
      r_4__55_ <= r_n_4__55_;
      r_4__54_ <= r_n_4__54_;
      r_4__53_ <= r_n_4__53_;
      r_4__52_ <= r_n_4__52_;
      r_4__51_ <= r_n_4__51_;
      r_4__50_ <= r_n_4__50_;
      r_4__49_ <= r_n_4__49_;
      r_4__48_ <= r_n_4__48_;
      r_4__47_ <= r_n_4__47_;
      r_4__46_ <= r_n_4__46_;
      r_4__45_ <= r_n_4__45_;
      r_4__44_ <= r_n_4__44_;
      r_4__43_ <= r_n_4__43_;
      r_4__42_ <= r_n_4__42_;
      r_4__41_ <= r_n_4__41_;
      r_4__40_ <= r_n_4__40_;
      r_4__39_ <= r_n_4__39_;
      r_4__38_ <= r_n_4__38_;
      r_4__37_ <= r_n_4__37_;
      r_4__36_ <= r_n_4__36_;
      r_4__35_ <= r_n_4__35_;
      r_4__34_ <= r_n_4__34_;
      r_4__33_ <= r_n_4__33_;
      r_4__32_ <= r_n_4__32_;
      r_4__31_ <= r_n_4__31_;
      r_4__30_ <= r_n_4__30_;
      r_4__29_ <= r_n_4__29_;
      r_4__28_ <= r_n_4__28_;
      r_4__27_ <= r_n_4__27_;
      r_4__26_ <= r_n_4__26_;
      r_4__25_ <= r_n_4__25_;
      r_4__24_ <= r_n_4__24_;
      r_4__23_ <= r_n_4__23_;
      r_4__22_ <= r_n_4__22_;
      r_4__21_ <= r_n_4__21_;
      r_4__20_ <= r_n_4__20_;
      r_4__19_ <= r_n_4__19_;
      r_4__18_ <= r_n_4__18_;
      r_4__17_ <= r_n_4__17_;
      r_4__16_ <= r_n_4__16_;
      r_4__15_ <= r_n_4__15_;
      r_4__14_ <= r_n_4__14_;
      r_4__13_ <= r_n_4__13_;
      r_4__12_ <= r_n_4__12_;
      r_4__11_ <= r_n_4__11_;
      r_4__10_ <= r_n_4__10_;
      r_4__9_ <= r_n_4__9_;
      r_4__8_ <= r_n_4__8_;
      r_4__7_ <= r_n_4__7_;
      r_4__6_ <= r_n_4__6_;
      r_4__5_ <= r_n_4__5_;
      r_4__4_ <= r_n_4__4_;
      r_4__3_ <= r_n_4__3_;
      r_4__2_ <= r_n_4__2_;
      r_4__1_ <= r_n_4__1_;
      r_4__0_ <= r_n_4__0_;
    end 
    if(N3589) begin
      r_5__63_ <= r_n_5__63_;
      r_5__62_ <= r_n_5__62_;
      r_5__61_ <= r_n_5__61_;
      r_5__60_ <= r_n_5__60_;
      r_5__59_ <= r_n_5__59_;
      r_5__58_ <= r_n_5__58_;
      r_5__57_ <= r_n_5__57_;
      r_5__56_ <= r_n_5__56_;
      r_5__55_ <= r_n_5__55_;
      r_5__54_ <= r_n_5__54_;
      r_5__53_ <= r_n_5__53_;
      r_5__52_ <= r_n_5__52_;
      r_5__51_ <= r_n_5__51_;
      r_5__50_ <= r_n_5__50_;
      r_5__49_ <= r_n_5__49_;
      r_5__48_ <= r_n_5__48_;
      r_5__47_ <= r_n_5__47_;
      r_5__46_ <= r_n_5__46_;
      r_5__45_ <= r_n_5__45_;
      r_5__44_ <= r_n_5__44_;
      r_5__43_ <= r_n_5__43_;
      r_5__42_ <= r_n_5__42_;
      r_5__41_ <= r_n_5__41_;
      r_5__40_ <= r_n_5__40_;
      r_5__39_ <= r_n_5__39_;
      r_5__38_ <= r_n_5__38_;
      r_5__37_ <= r_n_5__37_;
      r_5__36_ <= r_n_5__36_;
      r_5__35_ <= r_n_5__35_;
      r_5__34_ <= r_n_5__34_;
      r_5__33_ <= r_n_5__33_;
      r_5__32_ <= r_n_5__32_;
      r_5__31_ <= r_n_5__31_;
      r_5__30_ <= r_n_5__30_;
      r_5__29_ <= r_n_5__29_;
      r_5__28_ <= r_n_5__28_;
      r_5__27_ <= r_n_5__27_;
      r_5__26_ <= r_n_5__26_;
      r_5__25_ <= r_n_5__25_;
      r_5__24_ <= r_n_5__24_;
      r_5__23_ <= r_n_5__23_;
      r_5__22_ <= r_n_5__22_;
      r_5__21_ <= r_n_5__21_;
      r_5__20_ <= r_n_5__20_;
      r_5__19_ <= r_n_5__19_;
      r_5__18_ <= r_n_5__18_;
      r_5__17_ <= r_n_5__17_;
      r_5__16_ <= r_n_5__16_;
      r_5__15_ <= r_n_5__15_;
      r_5__14_ <= r_n_5__14_;
      r_5__13_ <= r_n_5__13_;
      r_5__12_ <= r_n_5__12_;
      r_5__11_ <= r_n_5__11_;
      r_5__10_ <= r_n_5__10_;
      r_5__9_ <= r_n_5__9_;
      r_5__8_ <= r_n_5__8_;
      r_5__7_ <= r_n_5__7_;
      r_5__6_ <= r_n_5__6_;
      r_5__5_ <= r_n_5__5_;
      r_5__4_ <= r_n_5__4_;
      r_5__3_ <= r_n_5__3_;
      r_5__2_ <= r_n_5__2_;
      r_5__1_ <= r_n_5__1_;
      r_5__0_ <= r_n_5__0_;
    end 
    if(N3590) begin
      r_6__63_ <= r_n_6__63_;
      r_6__62_ <= r_n_6__62_;
      r_6__61_ <= r_n_6__61_;
      r_6__60_ <= r_n_6__60_;
      r_6__59_ <= r_n_6__59_;
      r_6__58_ <= r_n_6__58_;
      r_6__57_ <= r_n_6__57_;
      r_6__56_ <= r_n_6__56_;
      r_6__55_ <= r_n_6__55_;
      r_6__54_ <= r_n_6__54_;
      r_6__53_ <= r_n_6__53_;
      r_6__52_ <= r_n_6__52_;
      r_6__51_ <= r_n_6__51_;
      r_6__50_ <= r_n_6__50_;
      r_6__49_ <= r_n_6__49_;
      r_6__48_ <= r_n_6__48_;
      r_6__47_ <= r_n_6__47_;
      r_6__46_ <= r_n_6__46_;
      r_6__45_ <= r_n_6__45_;
      r_6__44_ <= r_n_6__44_;
      r_6__43_ <= r_n_6__43_;
      r_6__42_ <= r_n_6__42_;
      r_6__41_ <= r_n_6__41_;
      r_6__40_ <= r_n_6__40_;
      r_6__39_ <= r_n_6__39_;
      r_6__38_ <= r_n_6__38_;
      r_6__37_ <= r_n_6__37_;
      r_6__36_ <= r_n_6__36_;
      r_6__35_ <= r_n_6__35_;
      r_6__34_ <= r_n_6__34_;
      r_6__33_ <= r_n_6__33_;
      r_6__32_ <= r_n_6__32_;
      r_6__31_ <= r_n_6__31_;
      r_6__30_ <= r_n_6__30_;
      r_6__29_ <= r_n_6__29_;
      r_6__28_ <= r_n_6__28_;
      r_6__27_ <= r_n_6__27_;
      r_6__26_ <= r_n_6__26_;
      r_6__25_ <= r_n_6__25_;
      r_6__24_ <= r_n_6__24_;
      r_6__23_ <= r_n_6__23_;
      r_6__22_ <= r_n_6__22_;
      r_6__21_ <= r_n_6__21_;
      r_6__20_ <= r_n_6__20_;
      r_6__19_ <= r_n_6__19_;
      r_6__18_ <= r_n_6__18_;
      r_6__17_ <= r_n_6__17_;
      r_6__16_ <= r_n_6__16_;
      r_6__15_ <= r_n_6__15_;
      r_6__14_ <= r_n_6__14_;
      r_6__13_ <= r_n_6__13_;
      r_6__12_ <= r_n_6__12_;
      r_6__11_ <= r_n_6__11_;
      r_6__10_ <= r_n_6__10_;
      r_6__9_ <= r_n_6__9_;
      r_6__8_ <= r_n_6__8_;
      r_6__7_ <= r_n_6__7_;
      r_6__6_ <= r_n_6__6_;
      r_6__5_ <= r_n_6__5_;
      r_6__4_ <= r_n_6__4_;
      r_6__3_ <= r_n_6__3_;
      r_6__2_ <= r_n_6__2_;
      r_6__1_ <= r_n_6__1_;
      r_6__0_ <= r_n_6__0_;
    end 
    if(N3591) begin
      r_7__63_ <= r_n_7__63_;
      r_7__62_ <= r_n_7__62_;
      r_7__61_ <= r_n_7__61_;
      r_7__60_ <= r_n_7__60_;
      r_7__59_ <= r_n_7__59_;
      r_7__58_ <= r_n_7__58_;
      r_7__57_ <= r_n_7__57_;
      r_7__56_ <= r_n_7__56_;
      r_7__55_ <= r_n_7__55_;
      r_7__54_ <= r_n_7__54_;
      r_7__53_ <= r_n_7__53_;
      r_7__52_ <= r_n_7__52_;
      r_7__51_ <= r_n_7__51_;
      r_7__50_ <= r_n_7__50_;
      r_7__49_ <= r_n_7__49_;
      r_7__48_ <= r_n_7__48_;
      r_7__47_ <= r_n_7__47_;
      r_7__46_ <= r_n_7__46_;
      r_7__45_ <= r_n_7__45_;
      r_7__44_ <= r_n_7__44_;
      r_7__43_ <= r_n_7__43_;
      r_7__42_ <= r_n_7__42_;
      r_7__41_ <= r_n_7__41_;
      r_7__40_ <= r_n_7__40_;
      r_7__39_ <= r_n_7__39_;
      r_7__38_ <= r_n_7__38_;
      r_7__37_ <= r_n_7__37_;
      r_7__36_ <= r_n_7__36_;
      r_7__35_ <= r_n_7__35_;
      r_7__34_ <= r_n_7__34_;
      r_7__33_ <= r_n_7__33_;
      r_7__32_ <= r_n_7__32_;
      r_7__31_ <= r_n_7__31_;
      r_7__30_ <= r_n_7__30_;
      r_7__29_ <= r_n_7__29_;
      r_7__28_ <= r_n_7__28_;
      r_7__27_ <= r_n_7__27_;
      r_7__26_ <= r_n_7__26_;
      r_7__25_ <= r_n_7__25_;
      r_7__24_ <= r_n_7__24_;
      r_7__23_ <= r_n_7__23_;
      r_7__22_ <= r_n_7__22_;
      r_7__21_ <= r_n_7__21_;
      r_7__20_ <= r_n_7__20_;
      r_7__19_ <= r_n_7__19_;
      r_7__18_ <= r_n_7__18_;
      r_7__17_ <= r_n_7__17_;
      r_7__16_ <= r_n_7__16_;
      r_7__15_ <= r_n_7__15_;
      r_7__14_ <= r_n_7__14_;
      r_7__13_ <= r_n_7__13_;
      r_7__12_ <= r_n_7__12_;
      r_7__11_ <= r_n_7__11_;
      r_7__10_ <= r_n_7__10_;
      r_7__9_ <= r_n_7__9_;
      r_7__8_ <= r_n_7__8_;
      r_7__7_ <= r_n_7__7_;
      r_7__6_ <= r_n_7__6_;
      r_7__5_ <= r_n_7__5_;
      r_7__4_ <= r_n_7__4_;
      r_7__3_ <= r_n_7__3_;
      r_7__2_ <= r_n_7__2_;
      r_7__1_ <= r_n_7__1_;
      r_7__0_ <= r_n_7__0_;
    end 
    if(N3592) begin
      r_8__63_ <= r_n_8__63_;
      r_8__62_ <= r_n_8__62_;
      r_8__61_ <= r_n_8__61_;
      r_8__60_ <= r_n_8__60_;
      r_8__59_ <= r_n_8__59_;
      r_8__58_ <= r_n_8__58_;
      r_8__57_ <= r_n_8__57_;
      r_8__56_ <= r_n_8__56_;
      r_8__55_ <= r_n_8__55_;
      r_8__54_ <= r_n_8__54_;
      r_8__53_ <= r_n_8__53_;
      r_8__52_ <= r_n_8__52_;
      r_8__51_ <= r_n_8__51_;
      r_8__50_ <= r_n_8__50_;
      r_8__49_ <= r_n_8__49_;
      r_8__48_ <= r_n_8__48_;
      r_8__47_ <= r_n_8__47_;
      r_8__46_ <= r_n_8__46_;
      r_8__45_ <= r_n_8__45_;
      r_8__44_ <= r_n_8__44_;
      r_8__43_ <= r_n_8__43_;
      r_8__42_ <= r_n_8__42_;
      r_8__41_ <= r_n_8__41_;
      r_8__40_ <= r_n_8__40_;
      r_8__39_ <= r_n_8__39_;
      r_8__38_ <= r_n_8__38_;
      r_8__37_ <= r_n_8__37_;
      r_8__36_ <= r_n_8__36_;
      r_8__35_ <= r_n_8__35_;
      r_8__34_ <= r_n_8__34_;
      r_8__33_ <= r_n_8__33_;
      r_8__32_ <= r_n_8__32_;
      r_8__31_ <= r_n_8__31_;
      r_8__30_ <= r_n_8__30_;
      r_8__29_ <= r_n_8__29_;
      r_8__28_ <= r_n_8__28_;
      r_8__27_ <= r_n_8__27_;
      r_8__26_ <= r_n_8__26_;
      r_8__25_ <= r_n_8__25_;
      r_8__24_ <= r_n_8__24_;
      r_8__23_ <= r_n_8__23_;
      r_8__22_ <= r_n_8__22_;
      r_8__21_ <= r_n_8__21_;
      r_8__20_ <= r_n_8__20_;
      r_8__19_ <= r_n_8__19_;
      r_8__18_ <= r_n_8__18_;
      r_8__17_ <= r_n_8__17_;
      r_8__16_ <= r_n_8__16_;
      r_8__15_ <= r_n_8__15_;
      r_8__14_ <= r_n_8__14_;
      r_8__13_ <= r_n_8__13_;
      r_8__12_ <= r_n_8__12_;
      r_8__11_ <= r_n_8__11_;
      r_8__10_ <= r_n_8__10_;
      r_8__9_ <= r_n_8__9_;
      r_8__8_ <= r_n_8__8_;
      r_8__7_ <= r_n_8__7_;
      r_8__6_ <= r_n_8__6_;
      r_8__5_ <= r_n_8__5_;
      r_8__4_ <= r_n_8__4_;
      r_8__3_ <= r_n_8__3_;
      r_8__2_ <= r_n_8__2_;
      r_8__1_ <= r_n_8__1_;
      r_8__0_ <= r_n_8__0_;
    end 
    if(N3593) begin
      r_9__63_ <= r_n_9__63_;
      r_9__62_ <= r_n_9__62_;
      r_9__61_ <= r_n_9__61_;
      r_9__60_ <= r_n_9__60_;
      r_9__59_ <= r_n_9__59_;
      r_9__58_ <= r_n_9__58_;
      r_9__57_ <= r_n_9__57_;
      r_9__56_ <= r_n_9__56_;
      r_9__55_ <= r_n_9__55_;
      r_9__54_ <= r_n_9__54_;
      r_9__53_ <= r_n_9__53_;
      r_9__52_ <= r_n_9__52_;
      r_9__51_ <= r_n_9__51_;
      r_9__50_ <= r_n_9__50_;
      r_9__49_ <= r_n_9__49_;
      r_9__48_ <= r_n_9__48_;
      r_9__47_ <= r_n_9__47_;
      r_9__46_ <= r_n_9__46_;
      r_9__45_ <= r_n_9__45_;
      r_9__44_ <= r_n_9__44_;
      r_9__43_ <= r_n_9__43_;
      r_9__42_ <= r_n_9__42_;
      r_9__41_ <= r_n_9__41_;
      r_9__40_ <= r_n_9__40_;
      r_9__39_ <= r_n_9__39_;
      r_9__38_ <= r_n_9__38_;
      r_9__37_ <= r_n_9__37_;
      r_9__36_ <= r_n_9__36_;
      r_9__35_ <= r_n_9__35_;
      r_9__34_ <= r_n_9__34_;
      r_9__33_ <= r_n_9__33_;
      r_9__32_ <= r_n_9__32_;
      r_9__31_ <= r_n_9__31_;
      r_9__30_ <= r_n_9__30_;
      r_9__29_ <= r_n_9__29_;
      r_9__28_ <= r_n_9__28_;
      r_9__27_ <= r_n_9__27_;
      r_9__26_ <= r_n_9__26_;
      r_9__25_ <= r_n_9__25_;
      r_9__24_ <= r_n_9__24_;
      r_9__23_ <= r_n_9__23_;
      r_9__22_ <= r_n_9__22_;
      r_9__21_ <= r_n_9__21_;
      r_9__20_ <= r_n_9__20_;
      r_9__19_ <= r_n_9__19_;
      r_9__18_ <= r_n_9__18_;
      r_9__17_ <= r_n_9__17_;
      r_9__16_ <= r_n_9__16_;
      r_9__15_ <= r_n_9__15_;
      r_9__14_ <= r_n_9__14_;
      r_9__13_ <= r_n_9__13_;
      r_9__12_ <= r_n_9__12_;
      r_9__11_ <= r_n_9__11_;
      r_9__10_ <= r_n_9__10_;
      r_9__9_ <= r_n_9__9_;
      r_9__8_ <= r_n_9__8_;
      r_9__7_ <= r_n_9__7_;
      r_9__6_ <= r_n_9__6_;
      r_9__5_ <= r_n_9__5_;
      r_9__4_ <= r_n_9__4_;
      r_9__3_ <= r_n_9__3_;
      r_9__2_ <= r_n_9__2_;
      r_9__1_ <= r_n_9__1_;
      r_9__0_ <= r_n_9__0_;
    end 
    if(N3594) begin
      r_10__63_ <= r_n_10__63_;
      r_10__62_ <= r_n_10__62_;
      r_10__61_ <= r_n_10__61_;
      r_10__60_ <= r_n_10__60_;
      r_10__59_ <= r_n_10__59_;
      r_10__58_ <= r_n_10__58_;
      r_10__57_ <= r_n_10__57_;
      r_10__56_ <= r_n_10__56_;
      r_10__55_ <= r_n_10__55_;
      r_10__54_ <= r_n_10__54_;
      r_10__53_ <= r_n_10__53_;
      r_10__52_ <= r_n_10__52_;
      r_10__51_ <= r_n_10__51_;
      r_10__50_ <= r_n_10__50_;
      r_10__49_ <= r_n_10__49_;
      r_10__48_ <= r_n_10__48_;
      r_10__47_ <= r_n_10__47_;
      r_10__46_ <= r_n_10__46_;
      r_10__45_ <= r_n_10__45_;
      r_10__44_ <= r_n_10__44_;
      r_10__43_ <= r_n_10__43_;
      r_10__42_ <= r_n_10__42_;
      r_10__41_ <= r_n_10__41_;
      r_10__40_ <= r_n_10__40_;
      r_10__39_ <= r_n_10__39_;
      r_10__38_ <= r_n_10__38_;
      r_10__37_ <= r_n_10__37_;
      r_10__36_ <= r_n_10__36_;
      r_10__35_ <= r_n_10__35_;
      r_10__34_ <= r_n_10__34_;
      r_10__33_ <= r_n_10__33_;
      r_10__32_ <= r_n_10__32_;
      r_10__31_ <= r_n_10__31_;
      r_10__30_ <= r_n_10__30_;
      r_10__29_ <= r_n_10__29_;
      r_10__28_ <= r_n_10__28_;
      r_10__27_ <= r_n_10__27_;
      r_10__26_ <= r_n_10__26_;
      r_10__25_ <= r_n_10__25_;
      r_10__24_ <= r_n_10__24_;
      r_10__23_ <= r_n_10__23_;
      r_10__22_ <= r_n_10__22_;
      r_10__21_ <= r_n_10__21_;
      r_10__20_ <= r_n_10__20_;
      r_10__19_ <= r_n_10__19_;
      r_10__18_ <= r_n_10__18_;
      r_10__17_ <= r_n_10__17_;
      r_10__16_ <= r_n_10__16_;
      r_10__15_ <= r_n_10__15_;
      r_10__14_ <= r_n_10__14_;
      r_10__13_ <= r_n_10__13_;
      r_10__12_ <= r_n_10__12_;
      r_10__11_ <= r_n_10__11_;
      r_10__10_ <= r_n_10__10_;
      r_10__9_ <= r_n_10__9_;
      r_10__8_ <= r_n_10__8_;
      r_10__7_ <= r_n_10__7_;
      r_10__6_ <= r_n_10__6_;
      r_10__5_ <= r_n_10__5_;
      r_10__4_ <= r_n_10__4_;
      r_10__3_ <= r_n_10__3_;
      r_10__2_ <= r_n_10__2_;
      r_10__1_ <= r_n_10__1_;
      r_10__0_ <= r_n_10__0_;
    end 
    if(N3595) begin
      r_11__63_ <= r_n_11__63_;
      r_11__62_ <= r_n_11__62_;
      r_11__61_ <= r_n_11__61_;
      r_11__60_ <= r_n_11__60_;
      r_11__59_ <= r_n_11__59_;
      r_11__58_ <= r_n_11__58_;
      r_11__57_ <= r_n_11__57_;
      r_11__56_ <= r_n_11__56_;
      r_11__55_ <= r_n_11__55_;
      r_11__54_ <= r_n_11__54_;
      r_11__53_ <= r_n_11__53_;
      r_11__52_ <= r_n_11__52_;
      r_11__51_ <= r_n_11__51_;
      r_11__50_ <= r_n_11__50_;
      r_11__49_ <= r_n_11__49_;
      r_11__48_ <= r_n_11__48_;
      r_11__47_ <= r_n_11__47_;
      r_11__46_ <= r_n_11__46_;
      r_11__45_ <= r_n_11__45_;
      r_11__44_ <= r_n_11__44_;
      r_11__43_ <= r_n_11__43_;
      r_11__42_ <= r_n_11__42_;
      r_11__41_ <= r_n_11__41_;
      r_11__40_ <= r_n_11__40_;
      r_11__39_ <= r_n_11__39_;
      r_11__38_ <= r_n_11__38_;
      r_11__37_ <= r_n_11__37_;
      r_11__36_ <= r_n_11__36_;
      r_11__35_ <= r_n_11__35_;
      r_11__34_ <= r_n_11__34_;
      r_11__33_ <= r_n_11__33_;
      r_11__32_ <= r_n_11__32_;
      r_11__31_ <= r_n_11__31_;
      r_11__30_ <= r_n_11__30_;
      r_11__29_ <= r_n_11__29_;
      r_11__28_ <= r_n_11__28_;
      r_11__27_ <= r_n_11__27_;
      r_11__26_ <= r_n_11__26_;
      r_11__25_ <= r_n_11__25_;
      r_11__24_ <= r_n_11__24_;
      r_11__23_ <= r_n_11__23_;
      r_11__22_ <= r_n_11__22_;
      r_11__21_ <= r_n_11__21_;
      r_11__20_ <= r_n_11__20_;
      r_11__19_ <= r_n_11__19_;
      r_11__18_ <= r_n_11__18_;
      r_11__17_ <= r_n_11__17_;
      r_11__16_ <= r_n_11__16_;
      r_11__15_ <= r_n_11__15_;
      r_11__14_ <= r_n_11__14_;
      r_11__13_ <= r_n_11__13_;
      r_11__12_ <= r_n_11__12_;
      r_11__11_ <= r_n_11__11_;
      r_11__10_ <= r_n_11__10_;
      r_11__9_ <= r_n_11__9_;
      r_11__8_ <= r_n_11__8_;
      r_11__7_ <= r_n_11__7_;
      r_11__6_ <= r_n_11__6_;
      r_11__5_ <= r_n_11__5_;
      r_11__4_ <= r_n_11__4_;
      r_11__3_ <= r_n_11__3_;
      r_11__2_ <= r_n_11__2_;
      r_11__1_ <= r_n_11__1_;
      r_11__0_ <= r_n_11__0_;
    end 
    if(N3596) begin
      r_12__63_ <= r_n_12__63_;
      r_12__62_ <= r_n_12__62_;
      r_12__61_ <= r_n_12__61_;
      r_12__60_ <= r_n_12__60_;
      r_12__59_ <= r_n_12__59_;
      r_12__58_ <= r_n_12__58_;
      r_12__57_ <= r_n_12__57_;
      r_12__56_ <= r_n_12__56_;
      r_12__55_ <= r_n_12__55_;
      r_12__54_ <= r_n_12__54_;
      r_12__53_ <= r_n_12__53_;
      r_12__52_ <= r_n_12__52_;
      r_12__51_ <= r_n_12__51_;
      r_12__50_ <= r_n_12__50_;
      r_12__49_ <= r_n_12__49_;
      r_12__48_ <= r_n_12__48_;
      r_12__47_ <= r_n_12__47_;
      r_12__46_ <= r_n_12__46_;
      r_12__45_ <= r_n_12__45_;
      r_12__44_ <= r_n_12__44_;
      r_12__43_ <= r_n_12__43_;
      r_12__42_ <= r_n_12__42_;
      r_12__41_ <= r_n_12__41_;
      r_12__40_ <= r_n_12__40_;
      r_12__39_ <= r_n_12__39_;
      r_12__38_ <= r_n_12__38_;
      r_12__37_ <= r_n_12__37_;
      r_12__36_ <= r_n_12__36_;
      r_12__35_ <= r_n_12__35_;
      r_12__34_ <= r_n_12__34_;
      r_12__33_ <= r_n_12__33_;
      r_12__32_ <= r_n_12__32_;
      r_12__31_ <= r_n_12__31_;
      r_12__30_ <= r_n_12__30_;
      r_12__29_ <= r_n_12__29_;
      r_12__28_ <= r_n_12__28_;
      r_12__27_ <= r_n_12__27_;
      r_12__26_ <= r_n_12__26_;
      r_12__25_ <= r_n_12__25_;
      r_12__24_ <= r_n_12__24_;
      r_12__23_ <= r_n_12__23_;
      r_12__22_ <= r_n_12__22_;
      r_12__21_ <= r_n_12__21_;
      r_12__20_ <= r_n_12__20_;
      r_12__19_ <= r_n_12__19_;
      r_12__18_ <= r_n_12__18_;
      r_12__17_ <= r_n_12__17_;
      r_12__16_ <= r_n_12__16_;
      r_12__15_ <= r_n_12__15_;
      r_12__14_ <= r_n_12__14_;
      r_12__13_ <= r_n_12__13_;
      r_12__12_ <= r_n_12__12_;
      r_12__11_ <= r_n_12__11_;
      r_12__10_ <= r_n_12__10_;
      r_12__9_ <= r_n_12__9_;
      r_12__8_ <= r_n_12__8_;
      r_12__7_ <= r_n_12__7_;
      r_12__6_ <= r_n_12__6_;
      r_12__5_ <= r_n_12__5_;
      r_12__4_ <= r_n_12__4_;
      r_12__3_ <= r_n_12__3_;
      r_12__2_ <= r_n_12__2_;
      r_12__1_ <= r_n_12__1_;
      r_12__0_ <= r_n_12__0_;
    end 
    if(N3597) begin
      r_13__63_ <= r_n_13__63_;
      r_13__62_ <= r_n_13__62_;
      r_13__61_ <= r_n_13__61_;
      r_13__60_ <= r_n_13__60_;
      r_13__59_ <= r_n_13__59_;
      r_13__58_ <= r_n_13__58_;
      r_13__57_ <= r_n_13__57_;
      r_13__56_ <= r_n_13__56_;
      r_13__55_ <= r_n_13__55_;
      r_13__54_ <= r_n_13__54_;
      r_13__53_ <= r_n_13__53_;
      r_13__52_ <= r_n_13__52_;
      r_13__51_ <= r_n_13__51_;
      r_13__50_ <= r_n_13__50_;
      r_13__49_ <= r_n_13__49_;
      r_13__48_ <= r_n_13__48_;
      r_13__47_ <= r_n_13__47_;
      r_13__46_ <= r_n_13__46_;
      r_13__45_ <= r_n_13__45_;
      r_13__44_ <= r_n_13__44_;
      r_13__43_ <= r_n_13__43_;
      r_13__42_ <= r_n_13__42_;
      r_13__41_ <= r_n_13__41_;
      r_13__40_ <= r_n_13__40_;
      r_13__39_ <= r_n_13__39_;
      r_13__38_ <= r_n_13__38_;
      r_13__37_ <= r_n_13__37_;
      r_13__36_ <= r_n_13__36_;
      r_13__35_ <= r_n_13__35_;
      r_13__34_ <= r_n_13__34_;
      r_13__33_ <= r_n_13__33_;
      r_13__32_ <= r_n_13__32_;
      r_13__31_ <= r_n_13__31_;
      r_13__30_ <= r_n_13__30_;
      r_13__29_ <= r_n_13__29_;
      r_13__28_ <= r_n_13__28_;
      r_13__27_ <= r_n_13__27_;
      r_13__26_ <= r_n_13__26_;
      r_13__25_ <= r_n_13__25_;
      r_13__24_ <= r_n_13__24_;
      r_13__23_ <= r_n_13__23_;
      r_13__22_ <= r_n_13__22_;
      r_13__21_ <= r_n_13__21_;
      r_13__20_ <= r_n_13__20_;
      r_13__19_ <= r_n_13__19_;
      r_13__18_ <= r_n_13__18_;
      r_13__17_ <= r_n_13__17_;
      r_13__16_ <= r_n_13__16_;
      r_13__15_ <= r_n_13__15_;
      r_13__14_ <= r_n_13__14_;
      r_13__13_ <= r_n_13__13_;
      r_13__12_ <= r_n_13__12_;
      r_13__11_ <= r_n_13__11_;
      r_13__10_ <= r_n_13__10_;
      r_13__9_ <= r_n_13__9_;
      r_13__8_ <= r_n_13__8_;
      r_13__7_ <= r_n_13__7_;
      r_13__6_ <= r_n_13__6_;
      r_13__5_ <= r_n_13__5_;
      r_13__4_ <= r_n_13__4_;
      r_13__3_ <= r_n_13__3_;
      r_13__2_ <= r_n_13__2_;
      r_13__1_ <= r_n_13__1_;
      r_13__0_ <= r_n_13__0_;
    end 
    if(N3598) begin
      r_14__63_ <= r_n_14__63_;
      r_14__62_ <= r_n_14__62_;
      r_14__61_ <= r_n_14__61_;
      r_14__60_ <= r_n_14__60_;
      r_14__59_ <= r_n_14__59_;
      r_14__58_ <= r_n_14__58_;
      r_14__57_ <= r_n_14__57_;
      r_14__56_ <= r_n_14__56_;
      r_14__55_ <= r_n_14__55_;
      r_14__54_ <= r_n_14__54_;
      r_14__53_ <= r_n_14__53_;
      r_14__52_ <= r_n_14__52_;
      r_14__51_ <= r_n_14__51_;
      r_14__50_ <= r_n_14__50_;
      r_14__49_ <= r_n_14__49_;
      r_14__48_ <= r_n_14__48_;
      r_14__47_ <= r_n_14__47_;
      r_14__46_ <= r_n_14__46_;
      r_14__45_ <= r_n_14__45_;
      r_14__44_ <= r_n_14__44_;
      r_14__43_ <= r_n_14__43_;
      r_14__42_ <= r_n_14__42_;
      r_14__41_ <= r_n_14__41_;
      r_14__40_ <= r_n_14__40_;
      r_14__39_ <= r_n_14__39_;
      r_14__38_ <= r_n_14__38_;
      r_14__37_ <= r_n_14__37_;
      r_14__36_ <= r_n_14__36_;
      r_14__35_ <= r_n_14__35_;
      r_14__34_ <= r_n_14__34_;
      r_14__33_ <= r_n_14__33_;
      r_14__32_ <= r_n_14__32_;
      r_14__31_ <= r_n_14__31_;
      r_14__30_ <= r_n_14__30_;
      r_14__29_ <= r_n_14__29_;
      r_14__28_ <= r_n_14__28_;
      r_14__27_ <= r_n_14__27_;
      r_14__26_ <= r_n_14__26_;
      r_14__25_ <= r_n_14__25_;
      r_14__24_ <= r_n_14__24_;
      r_14__23_ <= r_n_14__23_;
      r_14__22_ <= r_n_14__22_;
      r_14__21_ <= r_n_14__21_;
      r_14__20_ <= r_n_14__20_;
      r_14__19_ <= r_n_14__19_;
      r_14__18_ <= r_n_14__18_;
      r_14__17_ <= r_n_14__17_;
      r_14__16_ <= r_n_14__16_;
      r_14__15_ <= r_n_14__15_;
      r_14__14_ <= r_n_14__14_;
      r_14__13_ <= r_n_14__13_;
      r_14__12_ <= r_n_14__12_;
      r_14__11_ <= r_n_14__11_;
      r_14__10_ <= r_n_14__10_;
      r_14__9_ <= r_n_14__9_;
      r_14__8_ <= r_n_14__8_;
      r_14__7_ <= r_n_14__7_;
      r_14__6_ <= r_n_14__6_;
      r_14__5_ <= r_n_14__5_;
      r_14__4_ <= r_n_14__4_;
      r_14__3_ <= r_n_14__3_;
      r_14__2_ <= r_n_14__2_;
      r_14__1_ <= r_n_14__1_;
      r_14__0_ <= r_n_14__0_;
    end 
    if(N3599) begin
      r_15__63_ <= r_n_15__63_;
      r_15__62_ <= r_n_15__62_;
      r_15__61_ <= r_n_15__61_;
      r_15__60_ <= r_n_15__60_;
      r_15__59_ <= r_n_15__59_;
      r_15__58_ <= r_n_15__58_;
      r_15__57_ <= r_n_15__57_;
      r_15__56_ <= r_n_15__56_;
      r_15__55_ <= r_n_15__55_;
      r_15__54_ <= r_n_15__54_;
      r_15__53_ <= r_n_15__53_;
      r_15__52_ <= r_n_15__52_;
      r_15__51_ <= r_n_15__51_;
      r_15__50_ <= r_n_15__50_;
      r_15__49_ <= r_n_15__49_;
      r_15__48_ <= r_n_15__48_;
      r_15__47_ <= r_n_15__47_;
      r_15__46_ <= r_n_15__46_;
      r_15__45_ <= r_n_15__45_;
      r_15__44_ <= r_n_15__44_;
      r_15__43_ <= r_n_15__43_;
      r_15__42_ <= r_n_15__42_;
      r_15__41_ <= r_n_15__41_;
      r_15__40_ <= r_n_15__40_;
      r_15__39_ <= r_n_15__39_;
      r_15__38_ <= r_n_15__38_;
      r_15__37_ <= r_n_15__37_;
      r_15__36_ <= r_n_15__36_;
      r_15__35_ <= r_n_15__35_;
      r_15__34_ <= r_n_15__34_;
      r_15__33_ <= r_n_15__33_;
      r_15__32_ <= r_n_15__32_;
      r_15__31_ <= r_n_15__31_;
      r_15__30_ <= r_n_15__30_;
      r_15__29_ <= r_n_15__29_;
      r_15__28_ <= r_n_15__28_;
      r_15__27_ <= r_n_15__27_;
      r_15__26_ <= r_n_15__26_;
      r_15__25_ <= r_n_15__25_;
      r_15__24_ <= r_n_15__24_;
      r_15__23_ <= r_n_15__23_;
      r_15__22_ <= r_n_15__22_;
      r_15__21_ <= r_n_15__21_;
      r_15__20_ <= r_n_15__20_;
      r_15__19_ <= r_n_15__19_;
      r_15__18_ <= r_n_15__18_;
      r_15__17_ <= r_n_15__17_;
      r_15__16_ <= r_n_15__16_;
      r_15__15_ <= r_n_15__15_;
      r_15__14_ <= r_n_15__14_;
      r_15__13_ <= r_n_15__13_;
      r_15__12_ <= r_n_15__12_;
      r_15__11_ <= r_n_15__11_;
      r_15__10_ <= r_n_15__10_;
      r_15__9_ <= r_n_15__9_;
      r_15__8_ <= r_n_15__8_;
      r_15__7_ <= r_n_15__7_;
      r_15__6_ <= r_n_15__6_;
      r_15__5_ <= r_n_15__5_;
      r_15__4_ <= r_n_15__4_;
      r_15__3_ <= r_n_15__3_;
      r_15__2_ <= r_n_15__2_;
      r_15__1_ <= r_n_15__1_;
      r_15__0_ <= r_n_15__0_;
    end 
    if(N3600) begin
      r_16__63_ <= r_n_16__63_;
      r_16__62_ <= r_n_16__62_;
      r_16__61_ <= r_n_16__61_;
      r_16__60_ <= r_n_16__60_;
      r_16__59_ <= r_n_16__59_;
      r_16__58_ <= r_n_16__58_;
      r_16__57_ <= r_n_16__57_;
      r_16__56_ <= r_n_16__56_;
      r_16__55_ <= r_n_16__55_;
      r_16__54_ <= r_n_16__54_;
      r_16__53_ <= r_n_16__53_;
      r_16__52_ <= r_n_16__52_;
      r_16__51_ <= r_n_16__51_;
      r_16__50_ <= r_n_16__50_;
      r_16__49_ <= r_n_16__49_;
      r_16__48_ <= r_n_16__48_;
      r_16__47_ <= r_n_16__47_;
      r_16__46_ <= r_n_16__46_;
      r_16__45_ <= r_n_16__45_;
      r_16__44_ <= r_n_16__44_;
      r_16__43_ <= r_n_16__43_;
      r_16__42_ <= r_n_16__42_;
      r_16__41_ <= r_n_16__41_;
      r_16__40_ <= r_n_16__40_;
      r_16__39_ <= r_n_16__39_;
      r_16__38_ <= r_n_16__38_;
      r_16__37_ <= r_n_16__37_;
      r_16__36_ <= r_n_16__36_;
      r_16__35_ <= r_n_16__35_;
      r_16__34_ <= r_n_16__34_;
      r_16__33_ <= r_n_16__33_;
      r_16__32_ <= r_n_16__32_;
      r_16__31_ <= r_n_16__31_;
      r_16__30_ <= r_n_16__30_;
      r_16__29_ <= r_n_16__29_;
      r_16__28_ <= r_n_16__28_;
      r_16__27_ <= r_n_16__27_;
      r_16__26_ <= r_n_16__26_;
      r_16__25_ <= r_n_16__25_;
      r_16__24_ <= r_n_16__24_;
      r_16__23_ <= r_n_16__23_;
      r_16__22_ <= r_n_16__22_;
      r_16__21_ <= r_n_16__21_;
      r_16__20_ <= r_n_16__20_;
      r_16__19_ <= r_n_16__19_;
      r_16__18_ <= r_n_16__18_;
      r_16__17_ <= r_n_16__17_;
      r_16__16_ <= r_n_16__16_;
      r_16__15_ <= r_n_16__15_;
      r_16__14_ <= r_n_16__14_;
      r_16__13_ <= r_n_16__13_;
      r_16__12_ <= r_n_16__12_;
      r_16__11_ <= r_n_16__11_;
      r_16__10_ <= r_n_16__10_;
      r_16__9_ <= r_n_16__9_;
      r_16__8_ <= r_n_16__8_;
      r_16__7_ <= r_n_16__7_;
      r_16__6_ <= r_n_16__6_;
      r_16__5_ <= r_n_16__5_;
      r_16__4_ <= r_n_16__4_;
      r_16__3_ <= r_n_16__3_;
      r_16__2_ <= r_n_16__2_;
      r_16__1_ <= r_n_16__1_;
      r_16__0_ <= r_n_16__0_;
    end 
    if(N3601) begin
      r_17__63_ <= r_n_17__63_;
      r_17__62_ <= r_n_17__62_;
      r_17__61_ <= r_n_17__61_;
      r_17__60_ <= r_n_17__60_;
      r_17__59_ <= r_n_17__59_;
      r_17__58_ <= r_n_17__58_;
      r_17__57_ <= r_n_17__57_;
      r_17__56_ <= r_n_17__56_;
      r_17__55_ <= r_n_17__55_;
      r_17__54_ <= r_n_17__54_;
      r_17__53_ <= r_n_17__53_;
      r_17__52_ <= r_n_17__52_;
      r_17__51_ <= r_n_17__51_;
      r_17__50_ <= r_n_17__50_;
      r_17__49_ <= r_n_17__49_;
      r_17__48_ <= r_n_17__48_;
      r_17__47_ <= r_n_17__47_;
      r_17__46_ <= r_n_17__46_;
      r_17__45_ <= r_n_17__45_;
      r_17__44_ <= r_n_17__44_;
      r_17__43_ <= r_n_17__43_;
      r_17__42_ <= r_n_17__42_;
      r_17__41_ <= r_n_17__41_;
      r_17__40_ <= r_n_17__40_;
      r_17__39_ <= r_n_17__39_;
      r_17__38_ <= r_n_17__38_;
      r_17__37_ <= r_n_17__37_;
      r_17__36_ <= r_n_17__36_;
      r_17__35_ <= r_n_17__35_;
      r_17__34_ <= r_n_17__34_;
      r_17__33_ <= r_n_17__33_;
      r_17__32_ <= r_n_17__32_;
      r_17__31_ <= r_n_17__31_;
      r_17__30_ <= r_n_17__30_;
      r_17__29_ <= r_n_17__29_;
      r_17__28_ <= r_n_17__28_;
      r_17__27_ <= r_n_17__27_;
      r_17__26_ <= r_n_17__26_;
      r_17__25_ <= r_n_17__25_;
      r_17__24_ <= r_n_17__24_;
      r_17__23_ <= r_n_17__23_;
      r_17__22_ <= r_n_17__22_;
      r_17__21_ <= r_n_17__21_;
      r_17__20_ <= r_n_17__20_;
      r_17__19_ <= r_n_17__19_;
      r_17__18_ <= r_n_17__18_;
      r_17__17_ <= r_n_17__17_;
      r_17__16_ <= r_n_17__16_;
      r_17__15_ <= r_n_17__15_;
      r_17__14_ <= r_n_17__14_;
      r_17__13_ <= r_n_17__13_;
      r_17__12_ <= r_n_17__12_;
      r_17__11_ <= r_n_17__11_;
      r_17__10_ <= r_n_17__10_;
      r_17__9_ <= r_n_17__9_;
      r_17__8_ <= r_n_17__8_;
      r_17__7_ <= r_n_17__7_;
      r_17__6_ <= r_n_17__6_;
      r_17__5_ <= r_n_17__5_;
      r_17__4_ <= r_n_17__4_;
      r_17__3_ <= r_n_17__3_;
      r_17__2_ <= r_n_17__2_;
      r_17__1_ <= r_n_17__1_;
      r_17__0_ <= r_n_17__0_;
    end 
    if(N3602) begin
      r_18__63_ <= r_n_18__63_;
      r_18__62_ <= r_n_18__62_;
      r_18__61_ <= r_n_18__61_;
      r_18__60_ <= r_n_18__60_;
      r_18__59_ <= r_n_18__59_;
      r_18__58_ <= r_n_18__58_;
      r_18__57_ <= r_n_18__57_;
      r_18__56_ <= r_n_18__56_;
      r_18__55_ <= r_n_18__55_;
      r_18__54_ <= r_n_18__54_;
      r_18__53_ <= r_n_18__53_;
      r_18__52_ <= r_n_18__52_;
      r_18__51_ <= r_n_18__51_;
      r_18__50_ <= r_n_18__50_;
      r_18__49_ <= r_n_18__49_;
      r_18__48_ <= r_n_18__48_;
      r_18__47_ <= r_n_18__47_;
      r_18__46_ <= r_n_18__46_;
      r_18__45_ <= r_n_18__45_;
      r_18__44_ <= r_n_18__44_;
      r_18__43_ <= r_n_18__43_;
      r_18__42_ <= r_n_18__42_;
      r_18__41_ <= r_n_18__41_;
      r_18__40_ <= r_n_18__40_;
      r_18__39_ <= r_n_18__39_;
      r_18__38_ <= r_n_18__38_;
      r_18__37_ <= r_n_18__37_;
      r_18__36_ <= r_n_18__36_;
      r_18__35_ <= r_n_18__35_;
      r_18__34_ <= r_n_18__34_;
      r_18__33_ <= r_n_18__33_;
      r_18__32_ <= r_n_18__32_;
      r_18__31_ <= r_n_18__31_;
      r_18__30_ <= r_n_18__30_;
      r_18__29_ <= r_n_18__29_;
      r_18__28_ <= r_n_18__28_;
      r_18__27_ <= r_n_18__27_;
      r_18__26_ <= r_n_18__26_;
      r_18__25_ <= r_n_18__25_;
      r_18__24_ <= r_n_18__24_;
      r_18__23_ <= r_n_18__23_;
      r_18__22_ <= r_n_18__22_;
      r_18__21_ <= r_n_18__21_;
      r_18__20_ <= r_n_18__20_;
      r_18__19_ <= r_n_18__19_;
      r_18__18_ <= r_n_18__18_;
      r_18__17_ <= r_n_18__17_;
      r_18__16_ <= r_n_18__16_;
      r_18__15_ <= r_n_18__15_;
      r_18__14_ <= r_n_18__14_;
      r_18__13_ <= r_n_18__13_;
      r_18__12_ <= r_n_18__12_;
      r_18__11_ <= r_n_18__11_;
      r_18__10_ <= r_n_18__10_;
      r_18__9_ <= r_n_18__9_;
      r_18__8_ <= r_n_18__8_;
      r_18__7_ <= r_n_18__7_;
      r_18__6_ <= r_n_18__6_;
      r_18__5_ <= r_n_18__5_;
      r_18__4_ <= r_n_18__4_;
      r_18__3_ <= r_n_18__3_;
      r_18__2_ <= r_n_18__2_;
      r_18__1_ <= r_n_18__1_;
      r_18__0_ <= r_n_18__0_;
    end 
    if(N3603) begin
      r_19__63_ <= r_n_19__63_;
      r_19__62_ <= r_n_19__62_;
      r_19__61_ <= r_n_19__61_;
      r_19__60_ <= r_n_19__60_;
      r_19__59_ <= r_n_19__59_;
      r_19__58_ <= r_n_19__58_;
      r_19__57_ <= r_n_19__57_;
      r_19__56_ <= r_n_19__56_;
      r_19__55_ <= r_n_19__55_;
      r_19__54_ <= r_n_19__54_;
      r_19__53_ <= r_n_19__53_;
      r_19__52_ <= r_n_19__52_;
      r_19__51_ <= r_n_19__51_;
      r_19__50_ <= r_n_19__50_;
      r_19__49_ <= r_n_19__49_;
      r_19__48_ <= r_n_19__48_;
      r_19__47_ <= r_n_19__47_;
      r_19__46_ <= r_n_19__46_;
      r_19__45_ <= r_n_19__45_;
      r_19__44_ <= r_n_19__44_;
      r_19__43_ <= r_n_19__43_;
      r_19__42_ <= r_n_19__42_;
      r_19__41_ <= r_n_19__41_;
      r_19__40_ <= r_n_19__40_;
      r_19__39_ <= r_n_19__39_;
      r_19__38_ <= r_n_19__38_;
      r_19__37_ <= r_n_19__37_;
      r_19__36_ <= r_n_19__36_;
      r_19__35_ <= r_n_19__35_;
      r_19__34_ <= r_n_19__34_;
      r_19__33_ <= r_n_19__33_;
      r_19__32_ <= r_n_19__32_;
      r_19__31_ <= r_n_19__31_;
      r_19__30_ <= r_n_19__30_;
      r_19__29_ <= r_n_19__29_;
      r_19__28_ <= r_n_19__28_;
      r_19__27_ <= r_n_19__27_;
      r_19__26_ <= r_n_19__26_;
      r_19__25_ <= r_n_19__25_;
      r_19__24_ <= r_n_19__24_;
      r_19__23_ <= r_n_19__23_;
      r_19__22_ <= r_n_19__22_;
      r_19__21_ <= r_n_19__21_;
      r_19__20_ <= r_n_19__20_;
      r_19__19_ <= r_n_19__19_;
      r_19__18_ <= r_n_19__18_;
      r_19__17_ <= r_n_19__17_;
      r_19__16_ <= r_n_19__16_;
      r_19__15_ <= r_n_19__15_;
      r_19__14_ <= r_n_19__14_;
      r_19__13_ <= r_n_19__13_;
      r_19__12_ <= r_n_19__12_;
      r_19__11_ <= r_n_19__11_;
      r_19__10_ <= r_n_19__10_;
      r_19__9_ <= r_n_19__9_;
      r_19__8_ <= r_n_19__8_;
      r_19__7_ <= r_n_19__7_;
      r_19__6_ <= r_n_19__6_;
      r_19__5_ <= r_n_19__5_;
      r_19__4_ <= r_n_19__4_;
      r_19__3_ <= r_n_19__3_;
      r_19__2_ <= r_n_19__2_;
      r_19__1_ <= r_n_19__1_;
      r_19__0_ <= r_n_19__0_;
    end 
    if(N3604) begin
      r_20__63_ <= r_n_20__63_;
      r_20__62_ <= r_n_20__62_;
      r_20__61_ <= r_n_20__61_;
      r_20__60_ <= r_n_20__60_;
      r_20__59_ <= r_n_20__59_;
      r_20__58_ <= r_n_20__58_;
      r_20__57_ <= r_n_20__57_;
      r_20__56_ <= r_n_20__56_;
      r_20__55_ <= r_n_20__55_;
      r_20__54_ <= r_n_20__54_;
      r_20__53_ <= r_n_20__53_;
      r_20__52_ <= r_n_20__52_;
      r_20__51_ <= r_n_20__51_;
      r_20__50_ <= r_n_20__50_;
      r_20__49_ <= r_n_20__49_;
      r_20__48_ <= r_n_20__48_;
      r_20__47_ <= r_n_20__47_;
      r_20__46_ <= r_n_20__46_;
      r_20__45_ <= r_n_20__45_;
      r_20__44_ <= r_n_20__44_;
      r_20__43_ <= r_n_20__43_;
      r_20__42_ <= r_n_20__42_;
      r_20__41_ <= r_n_20__41_;
      r_20__40_ <= r_n_20__40_;
      r_20__39_ <= r_n_20__39_;
      r_20__38_ <= r_n_20__38_;
      r_20__37_ <= r_n_20__37_;
      r_20__36_ <= r_n_20__36_;
      r_20__35_ <= r_n_20__35_;
      r_20__34_ <= r_n_20__34_;
      r_20__33_ <= r_n_20__33_;
      r_20__32_ <= r_n_20__32_;
      r_20__31_ <= r_n_20__31_;
      r_20__30_ <= r_n_20__30_;
      r_20__29_ <= r_n_20__29_;
      r_20__28_ <= r_n_20__28_;
      r_20__27_ <= r_n_20__27_;
      r_20__26_ <= r_n_20__26_;
      r_20__25_ <= r_n_20__25_;
      r_20__24_ <= r_n_20__24_;
      r_20__23_ <= r_n_20__23_;
      r_20__22_ <= r_n_20__22_;
      r_20__21_ <= r_n_20__21_;
      r_20__20_ <= r_n_20__20_;
      r_20__19_ <= r_n_20__19_;
      r_20__18_ <= r_n_20__18_;
      r_20__17_ <= r_n_20__17_;
      r_20__16_ <= r_n_20__16_;
      r_20__15_ <= r_n_20__15_;
      r_20__14_ <= r_n_20__14_;
      r_20__13_ <= r_n_20__13_;
      r_20__12_ <= r_n_20__12_;
      r_20__11_ <= r_n_20__11_;
      r_20__10_ <= r_n_20__10_;
      r_20__9_ <= r_n_20__9_;
      r_20__8_ <= r_n_20__8_;
      r_20__7_ <= r_n_20__7_;
      r_20__6_ <= r_n_20__6_;
      r_20__5_ <= r_n_20__5_;
      r_20__4_ <= r_n_20__4_;
      r_20__3_ <= r_n_20__3_;
      r_20__2_ <= r_n_20__2_;
      r_20__1_ <= r_n_20__1_;
      r_20__0_ <= r_n_20__0_;
    end 
    if(N3605) begin
      r_21__63_ <= r_n_21__63_;
      r_21__62_ <= r_n_21__62_;
      r_21__61_ <= r_n_21__61_;
      r_21__60_ <= r_n_21__60_;
      r_21__59_ <= r_n_21__59_;
      r_21__58_ <= r_n_21__58_;
      r_21__57_ <= r_n_21__57_;
      r_21__56_ <= r_n_21__56_;
      r_21__55_ <= r_n_21__55_;
      r_21__54_ <= r_n_21__54_;
      r_21__53_ <= r_n_21__53_;
      r_21__52_ <= r_n_21__52_;
      r_21__51_ <= r_n_21__51_;
      r_21__50_ <= r_n_21__50_;
      r_21__49_ <= r_n_21__49_;
      r_21__48_ <= r_n_21__48_;
      r_21__47_ <= r_n_21__47_;
      r_21__46_ <= r_n_21__46_;
      r_21__45_ <= r_n_21__45_;
      r_21__44_ <= r_n_21__44_;
      r_21__43_ <= r_n_21__43_;
      r_21__42_ <= r_n_21__42_;
      r_21__41_ <= r_n_21__41_;
      r_21__40_ <= r_n_21__40_;
      r_21__39_ <= r_n_21__39_;
      r_21__38_ <= r_n_21__38_;
      r_21__37_ <= r_n_21__37_;
      r_21__36_ <= r_n_21__36_;
      r_21__35_ <= r_n_21__35_;
      r_21__34_ <= r_n_21__34_;
      r_21__33_ <= r_n_21__33_;
      r_21__32_ <= r_n_21__32_;
      r_21__31_ <= r_n_21__31_;
      r_21__30_ <= r_n_21__30_;
      r_21__29_ <= r_n_21__29_;
      r_21__28_ <= r_n_21__28_;
      r_21__27_ <= r_n_21__27_;
      r_21__26_ <= r_n_21__26_;
      r_21__25_ <= r_n_21__25_;
      r_21__24_ <= r_n_21__24_;
      r_21__23_ <= r_n_21__23_;
      r_21__22_ <= r_n_21__22_;
      r_21__21_ <= r_n_21__21_;
      r_21__20_ <= r_n_21__20_;
      r_21__19_ <= r_n_21__19_;
      r_21__18_ <= r_n_21__18_;
      r_21__17_ <= r_n_21__17_;
      r_21__16_ <= r_n_21__16_;
      r_21__15_ <= r_n_21__15_;
      r_21__14_ <= r_n_21__14_;
      r_21__13_ <= r_n_21__13_;
      r_21__12_ <= r_n_21__12_;
      r_21__11_ <= r_n_21__11_;
      r_21__10_ <= r_n_21__10_;
      r_21__9_ <= r_n_21__9_;
      r_21__8_ <= r_n_21__8_;
      r_21__7_ <= r_n_21__7_;
      r_21__6_ <= r_n_21__6_;
      r_21__5_ <= r_n_21__5_;
      r_21__4_ <= r_n_21__4_;
      r_21__3_ <= r_n_21__3_;
      r_21__2_ <= r_n_21__2_;
      r_21__1_ <= r_n_21__1_;
      r_21__0_ <= r_n_21__0_;
    end 
    if(N3606) begin
      r_22__63_ <= r_n_22__63_;
      r_22__62_ <= r_n_22__62_;
      r_22__61_ <= r_n_22__61_;
      r_22__60_ <= r_n_22__60_;
      r_22__59_ <= r_n_22__59_;
      r_22__58_ <= r_n_22__58_;
      r_22__57_ <= r_n_22__57_;
      r_22__56_ <= r_n_22__56_;
      r_22__55_ <= r_n_22__55_;
      r_22__54_ <= r_n_22__54_;
      r_22__53_ <= r_n_22__53_;
      r_22__52_ <= r_n_22__52_;
      r_22__51_ <= r_n_22__51_;
      r_22__50_ <= r_n_22__50_;
      r_22__49_ <= r_n_22__49_;
      r_22__48_ <= r_n_22__48_;
      r_22__47_ <= r_n_22__47_;
      r_22__46_ <= r_n_22__46_;
      r_22__45_ <= r_n_22__45_;
      r_22__44_ <= r_n_22__44_;
      r_22__43_ <= r_n_22__43_;
      r_22__42_ <= r_n_22__42_;
      r_22__41_ <= r_n_22__41_;
      r_22__40_ <= r_n_22__40_;
      r_22__39_ <= r_n_22__39_;
      r_22__38_ <= r_n_22__38_;
      r_22__37_ <= r_n_22__37_;
      r_22__36_ <= r_n_22__36_;
      r_22__35_ <= r_n_22__35_;
      r_22__34_ <= r_n_22__34_;
      r_22__33_ <= r_n_22__33_;
      r_22__32_ <= r_n_22__32_;
      r_22__31_ <= r_n_22__31_;
      r_22__30_ <= r_n_22__30_;
      r_22__29_ <= r_n_22__29_;
      r_22__28_ <= r_n_22__28_;
      r_22__27_ <= r_n_22__27_;
      r_22__26_ <= r_n_22__26_;
      r_22__25_ <= r_n_22__25_;
      r_22__24_ <= r_n_22__24_;
      r_22__23_ <= r_n_22__23_;
      r_22__22_ <= r_n_22__22_;
      r_22__21_ <= r_n_22__21_;
      r_22__20_ <= r_n_22__20_;
      r_22__19_ <= r_n_22__19_;
      r_22__18_ <= r_n_22__18_;
      r_22__17_ <= r_n_22__17_;
      r_22__16_ <= r_n_22__16_;
      r_22__15_ <= r_n_22__15_;
      r_22__14_ <= r_n_22__14_;
      r_22__13_ <= r_n_22__13_;
      r_22__12_ <= r_n_22__12_;
      r_22__11_ <= r_n_22__11_;
      r_22__10_ <= r_n_22__10_;
      r_22__9_ <= r_n_22__9_;
      r_22__8_ <= r_n_22__8_;
      r_22__7_ <= r_n_22__7_;
      r_22__6_ <= r_n_22__6_;
      r_22__5_ <= r_n_22__5_;
      r_22__4_ <= r_n_22__4_;
      r_22__3_ <= r_n_22__3_;
      r_22__2_ <= r_n_22__2_;
      r_22__1_ <= r_n_22__1_;
      r_22__0_ <= r_n_22__0_;
    end 
    if(N3607) begin
      r_23__63_ <= r_n_23__63_;
      r_23__62_ <= r_n_23__62_;
      r_23__61_ <= r_n_23__61_;
      r_23__60_ <= r_n_23__60_;
      r_23__59_ <= r_n_23__59_;
      r_23__58_ <= r_n_23__58_;
      r_23__57_ <= r_n_23__57_;
      r_23__56_ <= r_n_23__56_;
      r_23__55_ <= r_n_23__55_;
      r_23__54_ <= r_n_23__54_;
      r_23__53_ <= r_n_23__53_;
      r_23__52_ <= r_n_23__52_;
      r_23__51_ <= r_n_23__51_;
      r_23__50_ <= r_n_23__50_;
      r_23__49_ <= r_n_23__49_;
      r_23__48_ <= r_n_23__48_;
      r_23__47_ <= r_n_23__47_;
      r_23__46_ <= r_n_23__46_;
      r_23__45_ <= r_n_23__45_;
      r_23__44_ <= r_n_23__44_;
      r_23__43_ <= r_n_23__43_;
      r_23__42_ <= r_n_23__42_;
      r_23__41_ <= r_n_23__41_;
      r_23__40_ <= r_n_23__40_;
      r_23__39_ <= r_n_23__39_;
      r_23__38_ <= r_n_23__38_;
      r_23__37_ <= r_n_23__37_;
      r_23__36_ <= r_n_23__36_;
      r_23__35_ <= r_n_23__35_;
      r_23__34_ <= r_n_23__34_;
      r_23__33_ <= r_n_23__33_;
      r_23__32_ <= r_n_23__32_;
      r_23__31_ <= r_n_23__31_;
      r_23__30_ <= r_n_23__30_;
      r_23__29_ <= r_n_23__29_;
      r_23__28_ <= r_n_23__28_;
      r_23__27_ <= r_n_23__27_;
      r_23__26_ <= r_n_23__26_;
      r_23__25_ <= r_n_23__25_;
      r_23__24_ <= r_n_23__24_;
      r_23__23_ <= r_n_23__23_;
      r_23__22_ <= r_n_23__22_;
      r_23__21_ <= r_n_23__21_;
      r_23__20_ <= r_n_23__20_;
      r_23__19_ <= r_n_23__19_;
      r_23__18_ <= r_n_23__18_;
      r_23__17_ <= r_n_23__17_;
      r_23__16_ <= r_n_23__16_;
      r_23__15_ <= r_n_23__15_;
      r_23__14_ <= r_n_23__14_;
      r_23__13_ <= r_n_23__13_;
      r_23__12_ <= r_n_23__12_;
      r_23__11_ <= r_n_23__11_;
      r_23__10_ <= r_n_23__10_;
      r_23__9_ <= r_n_23__9_;
      r_23__8_ <= r_n_23__8_;
      r_23__7_ <= r_n_23__7_;
      r_23__6_ <= r_n_23__6_;
      r_23__5_ <= r_n_23__5_;
      r_23__4_ <= r_n_23__4_;
      r_23__3_ <= r_n_23__3_;
      r_23__2_ <= r_n_23__2_;
      r_23__1_ <= r_n_23__1_;
      r_23__0_ <= r_n_23__0_;
    end 
    if(N3608) begin
      r_24__63_ <= r_n_24__63_;
      r_24__62_ <= r_n_24__62_;
      r_24__61_ <= r_n_24__61_;
      r_24__60_ <= r_n_24__60_;
      r_24__59_ <= r_n_24__59_;
      r_24__58_ <= r_n_24__58_;
      r_24__57_ <= r_n_24__57_;
      r_24__56_ <= r_n_24__56_;
      r_24__55_ <= r_n_24__55_;
      r_24__54_ <= r_n_24__54_;
      r_24__53_ <= r_n_24__53_;
      r_24__52_ <= r_n_24__52_;
      r_24__51_ <= r_n_24__51_;
      r_24__50_ <= r_n_24__50_;
      r_24__49_ <= r_n_24__49_;
      r_24__48_ <= r_n_24__48_;
      r_24__47_ <= r_n_24__47_;
      r_24__46_ <= r_n_24__46_;
      r_24__45_ <= r_n_24__45_;
      r_24__44_ <= r_n_24__44_;
      r_24__43_ <= r_n_24__43_;
      r_24__42_ <= r_n_24__42_;
      r_24__41_ <= r_n_24__41_;
      r_24__40_ <= r_n_24__40_;
      r_24__39_ <= r_n_24__39_;
      r_24__38_ <= r_n_24__38_;
      r_24__37_ <= r_n_24__37_;
      r_24__36_ <= r_n_24__36_;
      r_24__35_ <= r_n_24__35_;
      r_24__34_ <= r_n_24__34_;
      r_24__33_ <= r_n_24__33_;
      r_24__32_ <= r_n_24__32_;
      r_24__31_ <= r_n_24__31_;
      r_24__30_ <= r_n_24__30_;
      r_24__29_ <= r_n_24__29_;
      r_24__28_ <= r_n_24__28_;
      r_24__27_ <= r_n_24__27_;
      r_24__26_ <= r_n_24__26_;
      r_24__25_ <= r_n_24__25_;
      r_24__24_ <= r_n_24__24_;
      r_24__23_ <= r_n_24__23_;
      r_24__22_ <= r_n_24__22_;
      r_24__21_ <= r_n_24__21_;
      r_24__20_ <= r_n_24__20_;
      r_24__19_ <= r_n_24__19_;
      r_24__18_ <= r_n_24__18_;
      r_24__17_ <= r_n_24__17_;
      r_24__16_ <= r_n_24__16_;
      r_24__15_ <= r_n_24__15_;
      r_24__14_ <= r_n_24__14_;
      r_24__13_ <= r_n_24__13_;
      r_24__12_ <= r_n_24__12_;
      r_24__11_ <= r_n_24__11_;
      r_24__10_ <= r_n_24__10_;
      r_24__9_ <= r_n_24__9_;
      r_24__8_ <= r_n_24__8_;
      r_24__7_ <= r_n_24__7_;
      r_24__6_ <= r_n_24__6_;
      r_24__5_ <= r_n_24__5_;
      r_24__4_ <= r_n_24__4_;
      r_24__3_ <= r_n_24__3_;
      r_24__2_ <= r_n_24__2_;
      r_24__1_ <= r_n_24__1_;
      r_24__0_ <= r_n_24__0_;
    end 
    if(N3609) begin
      r_25__63_ <= r_n_25__63_;
      r_25__62_ <= r_n_25__62_;
      r_25__61_ <= r_n_25__61_;
      r_25__60_ <= r_n_25__60_;
      r_25__59_ <= r_n_25__59_;
      r_25__58_ <= r_n_25__58_;
      r_25__57_ <= r_n_25__57_;
      r_25__56_ <= r_n_25__56_;
      r_25__55_ <= r_n_25__55_;
      r_25__54_ <= r_n_25__54_;
      r_25__53_ <= r_n_25__53_;
      r_25__52_ <= r_n_25__52_;
      r_25__51_ <= r_n_25__51_;
      r_25__50_ <= r_n_25__50_;
      r_25__49_ <= r_n_25__49_;
      r_25__48_ <= r_n_25__48_;
      r_25__47_ <= r_n_25__47_;
      r_25__46_ <= r_n_25__46_;
      r_25__45_ <= r_n_25__45_;
      r_25__44_ <= r_n_25__44_;
      r_25__43_ <= r_n_25__43_;
      r_25__42_ <= r_n_25__42_;
      r_25__41_ <= r_n_25__41_;
      r_25__40_ <= r_n_25__40_;
      r_25__39_ <= r_n_25__39_;
      r_25__38_ <= r_n_25__38_;
      r_25__37_ <= r_n_25__37_;
      r_25__36_ <= r_n_25__36_;
      r_25__35_ <= r_n_25__35_;
      r_25__34_ <= r_n_25__34_;
      r_25__33_ <= r_n_25__33_;
      r_25__32_ <= r_n_25__32_;
      r_25__31_ <= r_n_25__31_;
      r_25__30_ <= r_n_25__30_;
      r_25__29_ <= r_n_25__29_;
      r_25__28_ <= r_n_25__28_;
      r_25__27_ <= r_n_25__27_;
      r_25__26_ <= r_n_25__26_;
      r_25__25_ <= r_n_25__25_;
      r_25__24_ <= r_n_25__24_;
      r_25__23_ <= r_n_25__23_;
      r_25__22_ <= r_n_25__22_;
      r_25__21_ <= r_n_25__21_;
      r_25__20_ <= r_n_25__20_;
      r_25__19_ <= r_n_25__19_;
      r_25__18_ <= r_n_25__18_;
      r_25__17_ <= r_n_25__17_;
      r_25__16_ <= r_n_25__16_;
      r_25__15_ <= r_n_25__15_;
      r_25__14_ <= r_n_25__14_;
      r_25__13_ <= r_n_25__13_;
      r_25__12_ <= r_n_25__12_;
      r_25__11_ <= r_n_25__11_;
      r_25__10_ <= r_n_25__10_;
      r_25__9_ <= r_n_25__9_;
      r_25__8_ <= r_n_25__8_;
      r_25__7_ <= r_n_25__7_;
      r_25__6_ <= r_n_25__6_;
      r_25__5_ <= r_n_25__5_;
      r_25__4_ <= r_n_25__4_;
      r_25__3_ <= r_n_25__3_;
      r_25__2_ <= r_n_25__2_;
      r_25__1_ <= r_n_25__1_;
      r_25__0_ <= r_n_25__0_;
    end 
    if(N3610) begin
      r_26__63_ <= r_n_26__63_;
      r_26__62_ <= r_n_26__62_;
      r_26__61_ <= r_n_26__61_;
      r_26__60_ <= r_n_26__60_;
      r_26__59_ <= r_n_26__59_;
      r_26__58_ <= r_n_26__58_;
      r_26__57_ <= r_n_26__57_;
      r_26__56_ <= r_n_26__56_;
      r_26__55_ <= r_n_26__55_;
      r_26__54_ <= r_n_26__54_;
      r_26__53_ <= r_n_26__53_;
      r_26__52_ <= r_n_26__52_;
      r_26__51_ <= r_n_26__51_;
      r_26__50_ <= r_n_26__50_;
      r_26__49_ <= r_n_26__49_;
      r_26__48_ <= r_n_26__48_;
      r_26__47_ <= r_n_26__47_;
      r_26__46_ <= r_n_26__46_;
      r_26__45_ <= r_n_26__45_;
      r_26__44_ <= r_n_26__44_;
      r_26__43_ <= r_n_26__43_;
      r_26__42_ <= r_n_26__42_;
      r_26__41_ <= r_n_26__41_;
      r_26__40_ <= r_n_26__40_;
      r_26__39_ <= r_n_26__39_;
      r_26__38_ <= r_n_26__38_;
      r_26__37_ <= r_n_26__37_;
      r_26__36_ <= r_n_26__36_;
      r_26__35_ <= r_n_26__35_;
      r_26__34_ <= r_n_26__34_;
      r_26__33_ <= r_n_26__33_;
      r_26__32_ <= r_n_26__32_;
      r_26__31_ <= r_n_26__31_;
      r_26__30_ <= r_n_26__30_;
      r_26__29_ <= r_n_26__29_;
      r_26__28_ <= r_n_26__28_;
      r_26__27_ <= r_n_26__27_;
      r_26__26_ <= r_n_26__26_;
      r_26__25_ <= r_n_26__25_;
      r_26__24_ <= r_n_26__24_;
      r_26__23_ <= r_n_26__23_;
      r_26__22_ <= r_n_26__22_;
      r_26__21_ <= r_n_26__21_;
      r_26__20_ <= r_n_26__20_;
      r_26__19_ <= r_n_26__19_;
      r_26__18_ <= r_n_26__18_;
      r_26__17_ <= r_n_26__17_;
      r_26__16_ <= r_n_26__16_;
      r_26__15_ <= r_n_26__15_;
      r_26__14_ <= r_n_26__14_;
      r_26__13_ <= r_n_26__13_;
      r_26__12_ <= r_n_26__12_;
      r_26__11_ <= r_n_26__11_;
      r_26__10_ <= r_n_26__10_;
      r_26__9_ <= r_n_26__9_;
      r_26__8_ <= r_n_26__8_;
      r_26__7_ <= r_n_26__7_;
      r_26__6_ <= r_n_26__6_;
      r_26__5_ <= r_n_26__5_;
      r_26__4_ <= r_n_26__4_;
      r_26__3_ <= r_n_26__3_;
      r_26__2_ <= r_n_26__2_;
      r_26__1_ <= r_n_26__1_;
      r_26__0_ <= r_n_26__0_;
    end 
    if(N3611) begin
      r_27__63_ <= r_n_27__63_;
      r_27__62_ <= r_n_27__62_;
      r_27__61_ <= r_n_27__61_;
      r_27__60_ <= r_n_27__60_;
      r_27__59_ <= r_n_27__59_;
      r_27__58_ <= r_n_27__58_;
      r_27__57_ <= r_n_27__57_;
      r_27__56_ <= r_n_27__56_;
      r_27__55_ <= r_n_27__55_;
      r_27__54_ <= r_n_27__54_;
      r_27__53_ <= r_n_27__53_;
      r_27__52_ <= r_n_27__52_;
      r_27__51_ <= r_n_27__51_;
      r_27__50_ <= r_n_27__50_;
      r_27__49_ <= r_n_27__49_;
      r_27__48_ <= r_n_27__48_;
      r_27__47_ <= r_n_27__47_;
      r_27__46_ <= r_n_27__46_;
      r_27__45_ <= r_n_27__45_;
      r_27__44_ <= r_n_27__44_;
      r_27__43_ <= r_n_27__43_;
      r_27__42_ <= r_n_27__42_;
      r_27__41_ <= r_n_27__41_;
      r_27__40_ <= r_n_27__40_;
      r_27__39_ <= r_n_27__39_;
      r_27__38_ <= r_n_27__38_;
      r_27__37_ <= r_n_27__37_;
      r_27__36_ <= r_n_27__36_;
      r_27__35_ <= r_n_27__35_;
      r_27__34_ <= r_n_27__34_;
      r_27__33_ <= r_n_27__33_;
      r_27__32_ <= r_n_27__32_;
      r_27__31_ <= r_n_27__31_;
      r_27__30_ <= r_n_27__30_;
      r_27__29_ <= r_n_27__29_;
      r_27__28_ <= r_n_27__28_;
      r_27__27_ <= r_n_27__27_;
      r_27__26_ <= r_n_27__26_;
      r_27__25_ <= r_n_27__25_;
      r_27__24_ <= r_n_27__24_;
      r_27__23_ <= r_n_27__23_;
      r_27__22_ <= r_n_27__22_;
      r_27__21_ <= r_n_27__21_;
      r_27__20_ <= r_n_27__20_;
      r_27__19_ <= r_n_27__19_;
      r_27__18_ <= r_n_27__18_;
      r_27__17_ <= r_n_27__17_;
      r_27__16_ <= r_n_27__16_;
      r_27__15_ <= r_n_27__15_;
      r_27__14_ <= r_n_27__14_;
      r_27__13_ <= r_n_27__13_;
      r_27__12_ <= r_n_27__12_;
      r_27__11_ <= r_n_27__11_;
      r_27__10_ <= r_n_27__10_;
      r_27__9_ <= r_n_27__9_;
      r_27__8_ <= r_n_27__8_;
      r_27__7_ <= r_n_27__7_;
      r_27__6_ <= r_n_27__6_;
      r_27__5_ <= r_n_27__5_;
      r_27__4_ <= r_n_27__4_;
      r_27__3_ <= r_n_27__3_;
      r_27__2_ <= r_n_27__2_;
      r_27__1_ <= r_n_27__1_;
      r_27__0_ <= r_n_27__0_;
    end 
    if(N3612) begin
      r_28__63_ <= r_n_28__63_;
      r_28__62_ <= r_n_28__62_;
      r_28__61_ <= r_n_28__61_;
      r_28__60_ <= r_n_28__60_;
      r_28__59_ <= r_n_28__59_;
      r_28__58_ <= r_n_28__58_;
      r_28__57_ <= r_n_28__57_;
      r_28__56_ <= r_n_28__56_;
      r_28__55_ <= r_n_28__55_;
      r_28__54_ <= r_n_28__54_;
      r_28__53_ <= r_n_28__53_;
      r_28__52_ <= r_n_28__52_;
      r_28__51_ <= r_n_28__51_;
      r_28__50_ <= r_n_28__50_;
      r_28__49_ <= r_n_28__49_;
      r_28__48_ <= r_n_28__48_;
      r_28__47_ <= r_n_28__47_;
      r_28__46_ <= r_n_28__46_;
      r_28__45_ <= r_n_28__45_;
      r_28__44_ <= r_n_28__44_;
      r_28__43_ <= r_n_28__43_;
      r_28__42_ <= r_n_28__42_;
      r_28__41_ <= r_n_28__41_;
      r_28__40_ <= r_n_28__40_;
      r_28__39_ <= r_n_28__39_;
      r_28__38_ <= r_n_28__38_;
      r_28__37_ <= r_n_28__37_;
      r_28__36_ <= r_n_28__36_;
      r_28__35_ <= r_n_28__35_;
      r_28__34_ <= r_n_28__34_;
      r_28__33_ <= r_n_28__33_;
      r_28__32_ <= r_n_28__32_;
      r_28__31_ <= r_n_28__31_;
      r_28__30_ <= r_n_28__30_;
      r_28__29_ <= r_n_28__29_;
      r_28__28_ <= r_n_28__28_;
      r_28__27_ <= r_n_28__27_;
      r_28__26_ <= r_n_28__26_;
      r_28__25_ <= r_n_28__25_;
      r_28__24_ <= r_n_28__24_;
      r_28__23_ <= r_n_28__23_;
      r_28__22_ <= r_n_28__22_;
      r_28__21_ <= r_n_28__21_;
      r_28__20_ <= r_n_28__20_;
      r_28__19_ <= r_n_28__19_;
      r_28__18_ <= r_n_28__18_;
      r_28__17_ <= r_n_28__17_;
      r_28__16_ <= r_n_28__16_;
      r_28__15_ <= r_n_28__15_;
      r_28__14_ <= r_n_28__14_;
      r_28__13_ <= r_n_28__13_;
      r_28__12_ <= r_n_28__12_;
      r_28__11_ <= r_n_28__11_;
      r_28__10_ <= r_n_28__10_;
      r_28__9_ <= r_n_28__9_;
      r_28__8_ <= r_n_28__8_;
      r_28__7_ <= r_n_28__7_;
      r_28__6_ <= r_n_28__6_;
      r_28__5_ <= r_n_28__5_;
      r_28__4_ <= r_n_28__4_;
      r_28__3_ <= r_n_28__3_;
      r_28__2_ <= r_n_28__2_;
      r_28__1_ <= r_n_28__1_;
      r_28__0_ <= r_n_28__0_;
    end 
    if(N3613) begin
      r_29__63_ <= r_n_29__63_;
      r_29__62_ <= r_n_29__62_;
      r_29__61_ <= r_n_29__61_;
      r_29__60_ <= r_n_29__60_;
      r_29__59_ <= r_n_29__59_;
      r_29__58_ <= r_n_29__58_;
      r_29__57_ <= r_n_29__57_;
      r_29__56_ <= r_n_29__56_;
      r_29__55_ <= r_n_29__55_;
      r_29__54_ <= r_n_29__54_;
      r_29__53_ <= r_n_29__53_;
      r_29__52_ <= r_n_29__52_;
      r_29__51_ <= r_n_29__51_;
      r_29__50_ <= r_n_29__50_;
      r_29__49_ <= r_n_29__49_;
      r_29__48_ <= r_n_29__48_;
      r_29__47_ <= r_n_29__47_;
      r_29__46_ <= r_n_29__46_;
      r_29__45_ <= r_n_29__45_;
      r_29__44_ <= r_n_29__44_;
      r_29__43_ <= r_n_29__43_;
      r_29__42_ <= r_n_29__42_;
      r_29__41_ <= r_n_29__41_;
      r_29__40_ <= r_n_29__40_;
      r_29__39_ <= r_n_29__39_;
      r_29__38_ <= r_n_29__38_;
      r_29__37_ <= r_n_29__37_;
      r_29__36_ <= r_n_29__36_;
      r_29__35_ <= r_n_29__35_;
      r_29__34_ <= r_n_29__34_;
      r_29__33_ <= r_n_29__33_;
      r_29__32_ <= r_n_29__32_;
      r_29__31_ <= r_n_29__31_;
      r_29__30_ <= r_n_29__30_;
      r_29__29_ <= r_n_29__29_;
      r_29__28_ <= r_n_29__28_;
      r_29__27_ <= r_n_29__27_;
      r_29__26_ <= r_n_29__26_;
      r_29__25_ <= r_n_29__25_;
      r_29__24_ <= r_n_29__24_;
      r_29__23_ <= r_n_29__23_;
      r_29__22_ <= r_n_29__22_;
      r_29__21_ <= r_n_29__21_;
      r_29__20_ <= r_n_29__20_;
      r_29__19_ <= r_n_29__19_;
      r_29__18_ <= r_n_29__18_;
      r_29__17_ <= r_n_29__17_;
      r_29__16_ <= r_n_29__16_;
      r_29__15_ <= r_n_29__15_;
      r_29__14_ <= r_n_29__14_;
      r_29__13_ <= r_n_29__13_;
      r_29__12_ <= r_n_29__12_;
      r_29__11_ <= r_n_29__11_;
      r_29__10_ <= r_n_29__10_;
      r_29__9_ <= r_n_29__9_;
      r_29__8_ <= r_n_29__8_;
      r_29__7_ <= r_n_29__7_;
      r_29__6_ <= r_n_29__6_;
      r_29__5_ <= r_n_29__5_;
      r_29__4_ <= r_n_29__4_;
      r_29__3_ <= r_n_29__3_;
      r_29__2_ <= r_n_29__2_;
      r_29__1_ <= r_n_29__1_;
      r_29__0_ <= r_n_29__0_;
    end 
    if(N3614) begin
      r_30__63_ <= r_n_30__63_;
      r_30__62_ <= r_n_30__62_;
      r_30__61_ <= r_n_30__61_;
      r_30__60_ <= r_n_30__60_;
      r_30__59_ <= r_n_30__59_;
      r_30__58_ <= r_n_30__58_;
      r_30__57_ <= r_n_30__57_;
      r_30__56_ <= r_n_30__56_;
      r_30__55_ <= r_n_30__55_;
      r_30__54_ <= r_n_30__54_;
      r_30__53_ <= r_n_30__53_;
      r_30__52_ <= r_n_30__52_;
      r_30__51_ <= r_n_30__51_;
      r_30__50_ <= r_n_30__50_;
      r_30__49_ <= r_n_30__49_;
      r_30__48_ <= r_n_30__48_;
      r_30__47_ <= r_n_30__47_;
      r_30__46_ <= r_n_30__46_;
      r_30__45_ <= r_n_30__45_;
      r_30__44_ <= r_n_30__44_;
      r_30__43_ <= r_n_30__43_;
      r_30__42_ <= r_n_30__42_;
      r_30__41_ <= r_n_30__41_;
      r_30__40_ <= r_n_30__40_;
      r_30__39_ <= r_n_30__39_;
      r_30__38_ <= r_n_30__38_;
      r_30__37_ <= r_n_30__37_;
      r_30__36_ <= r_n_30__36_;
      r_30__35_ <= r_n_30__35_;
      r_30__34_ <= r_n_30__34_;
      r_30__33_ <= r_n_30__33_;
      r_30__32_ <= r_n_30__32_;
      r_30__31_ <= r_n_30__31_;
      r_30__30_ <= r_n_30__30_;
      r_30__29_ <= r_n_30__29_;
      r_30__28_ <= r_n_30__28_;
      r_30__27_ <= r_n_30__27_;
      r_30__26_ <= r_n_30__26_;
      r_30__25_ <= r_n_30__25_;
      r_30__24_ <= r_n_30__24_;
      r_30__23_ <= r_n_30__23_;
      r_30__22_ <= r_n_30__22_;
      r_30__21_ <= r_n_30__21_;
      r_30__20_ <= r_n_30__20_;
      r_30__19_ <= r_n_30__19_;
      r_30__18_ <= r_n_30__18_;
      r_30__17_ <= r_n_30__17_;
      r_30__16_ <= r_n_30__16_;
      r_30__15_ <= r_n_30__15_;
      r_30__14_ <= r_n_30__14_;
      r_30__13_ <= r_n_30__13_;
      r_30__12_ <= r_n_30__12_;
      r_30__11_ <= r_n_30__11_;
      r_30__10_ <= r_n_30__10_;
      r_30__9_ <= r_n_30__9_;
      r_30__8_ <= r_n_30__8_;
      r_30__7_ <= r_n_30__7_;
      r_30__6_ <= r_n_30__6_;
      r_30__5_ <= r_n_30__5_;
      r_30__4_ <= r_n_30__4_;
      r_30__3_ <= r_n_30__3_;
      r_30__2_ <= r_n_30__2_;
      r_30__1_ <= r_n_30__1_;
      r_30__0_ <= r_n_30__0_;
    end 
    if(N3615) begin
      r_31__63_ <= r_n_31__63_;
      r_31__62_ <= r_n_31__62_;
      r_31__61_ <= r_n_31__61_;
      r_31__60_ <= r_n_31__60_;
      r_31__59_ <= r_n_31__59_;
      r_31__58_ <= r_n_31__58_;
      r_31__57_ <= r_n_31__57_;
      r_31__56_ <= r_n_31__56_;
      r_31__55_ <= r_n_31__55_;
      r_31__54_ <= r_n_31__54_;
      r_31__53_ <= r_n_31__53_;
      r_31__52_ <= r_n_31__52_;
      r_31__51_ <= r_n_31__51_;
      r_31__50_ <= r_n_31__50_;
      r_31__49_ <= r_n_31__49_;
      r_31__48_ <= r_n_31__48_;
      r_31__47_ <= r_n_31__47_;
      r_31__46_ <= r_n_31__46_;
      r_31__45_ <= r_n_31__45_;
      r_31__44_ <= r_n_31__44_;
      r_31__43_ <= r_n_31__43_;
      r_31__42_ <= r_n_31__42_;
      r_31__41_ <= r_n_31__41_;
      r_31__40_ <= r_n_31__40_;
      r_31__39_ <= r_n_31__39_;
      r_31__38_ <= r_n_31__38_;
      r_31__37_ <= r_n_31__37_;
      r_31__36_ <= r_n_31__36_;
      r_31__35_ <= r_n_31__35_;
      r_31__34_ <= r_n_31__34_;
      r_31__33_ <= r_n_31__33_;
      r_31__32_ <= r_n_31__32_;
      r_31__31_ <= r_n_31__31_;
      r_31__30_ <= r_n_31__30_;
      r_31__29_ <= r_n_31__29_;
      r_31__28_ <= r_n_31__28_;
      r_31__27_ <= r_n_31__27_;
      r_31__26_ <= r_n_31__26_;
      r_31__25_ <= r_n_31__25_;
      r_31__24_ <= r_n_31__24_;
      r_31__23_ <= r_n_31__23_;
      r_31__22_ <= r_n_31__22_;
      r_31__21_ <= r_n_31__21_;
      r_31__20_ <= r_n_31__20_;
      r_31__19_ <= r_n_31__19_;
      r_31__18_ <= r_n_31__18_;
      r_31__17_ <= r_n_31__17_;
      r_31__16_ <= r_n_31__16_;
      r_31__15_ <= r_n_31__15_;
      r_31__14_ <= r_n_31__14_;
      r_31__13_ <= r_n_31__13_;
      r_31__12_ <= r_n_31__12_;
      r_31__11_ <= r_n_31__11_;
      r_31__10_ <= r_n_31__10_;
      r_31__9_ <= r_n_31__9_;
      r_31__8_ <= r_n_31__8_;
      r_31__7_ <= r_n_31__7_;
      r_31__6_ <= r_n_31__6_;
      r_31__5_ <= r_n_31__5_;
      r_31__4_ <= r_n_31__4_;
      r_31__3_ <= r_n_31__3_;
      r_31__2_ <= r_n_31__2_;
      r_31__1_ <= r_n_31__1_;
      r_31__0_ <= r_n_31__0_;
    end 
    if(N3616) begin
      r_32__63_ <= r_n_32__63_;
      r_32__62_ <= r_n_32__62_;
      r_32__61_ <= r_n_32__61_;
      r_32__60_ <= r_n_32__60_;
      r_32__59_ <= r_n_32__59_;
      r_32__58_ <= r_n_32__58_;
      r_32__57_ <= r_n_32__57_;
      r_32__56_ <= r_n_32__56_;
      r_32__55_ <= r_n_32__55_;
      r_32__54_ <= r_n_32__54_;
      r_32__53_ <= r_n_32__53_;
      r_32__52_ <= r_n_32__52_;
      r_32__51_ <= r_n_32__51_;
      r_32__50_ <= r_n_32__50_;
      r_32__49_ <= r_n_32__49_;
      r_32__48_ <= r_n_32__48_;
      r_32__47_ <= r_n_32__47_;
      r_32__46_ <= r_n_32__46_;
      r_32__45_ <= r_n_32__45_;
      r_32__44_ <= r_n_32__44_;
      r_32__43_ <= r_n_32__43_;
      r_32__42_ <= r_n_32__42_;
      r_32__41_ <= r_n_32__41_;
      r_32__40_ <= r_n_32__40_;
      r_32__39_ <= r_n_32__39_;
      r_32__38_ <= r_n_32__38_;
      r_32__37_ <= r_n_32__37_;
      r_32__36_ <= r_n_32__36_;
      r_32__35_ <= r_n_32__35_;
      r_32__34_ <= r_n_32__34_;
      r_32__33_ <= r_n_32__33_;
      r_32__32_ <= r_n_32__32_;
      r_32__31_ <= r_n_32__31_;
      r_32__30_ <= r_n_32__30_;
      r_32__29_ <= r_n_32__29_;
      r_32__28_ <= r_n_32__28_;
      r_32__27_ <= r_n_32__27_;
      r_32__26_ <= r_n_32__26_;
      r_32__25_ <= r_n_32__25_;
      r_32__24_ <= r_n_32__24_;
      r_32__23_ <= r_n_32__23_;
      r_32__22_ <= r_n_32__22_;
      r_32__21_ <= r_n_32__21_;
      r_32__20_ <= r_n_32__20_;
      r_32__19_ <= r_n_32__19_;
      r_32__18_ <= r_n_32__18_;
      r_32__17_ <= r_n_32__17_;
      r_32__16_ <= r_n_32__16_;
      r_32__15_ <= r_n_32__15_;
      r_32__14_ <= r_n_32__14_;
      r_32__13_ <= r_n_32__13_;
      r_32__12_ <= r_n_32__12_;
      r_32__11_ <= r_n_32__11_;
      r_32__10_ <= r_n_32__10_;
      r_32__9_ <= r_n_32__9_;
      r_32__8_ <= r_n_32__8_;
      r_32__7_ <= r_n_32__7_;
      r_32__6_ <= r_n_32__6_;
      r_32__5_ <= r_n_32__5_;
      r_32__4_ <= r_n_32__4_;
      r_32__3_ <= r_n_32__3_;
      r_32__2_ <= r_n_32__2_;
      r_32__1_ <= r_n_32__1_;
      r_32__0_ <= r_n_32__0_;
    end 
    if(N3617) begin
      r_33__63_ <= r_n_33__63_;
      r_33__62_ <= r_n_33__62_;
      r_33__61_ <= r_n_33__61_;
      r_33__60_ <= r_n_33__60_;
      r_33__59_ <= r_n_33__59_;
      r_33__58_ <= r_n_33__58_;
      r_33__57_ <= r_n_33__57_;
      r_33__56_ <= r_n_33__56_;
      r_33__55_ <= r_n_33__55_;
      r_33__54_ <= r_n_33__54_;
      r_33__53_ <= r_n_33__53_;
      r_33__52_ <= r_n_33__52_;
      r_33__51_ <= r_n_33__51_;
      r_33__50_ <= r_n_33__50_;
      r_33__49_ <= r_n_33__49_;
      r_33__48_ <= r_n_33__48_;
      r_33__47_ <= r_n_33__47_;
      r_33__46_ <= r_n_33__46_;
      r_33__45_ <= r_n_33__45_;
      r_33__44_ <= r_n_33__44_;
      r_33__43_ <= r_n_33__43_;
      r_33__42_ <= r_n_33__42_;
      r_33__41_ <= r_n_33__41_;
      r_33__40_ <= r_n_33__40_;
      r_33__39_ <= r_n_33__39_;
      r_33__38_ <= r_n_33__38_;
      r_33__37_ <= r_n_33__37_;
      r_33__36_ <= r_n_33__36_;
      r_33__35_ <= r_n_33__35_;
      r_33__34_ <= r_n_33__34_;
      r_33__33_ <= r_n_33__33_;
      r_33__32_ <= r_n_33__32_;
      r_33__31_ <= r_n_33__31_;
      r_33__30_ <= r_n_33__30_;
      r_33__29_ <= r_n_33__29_;
      r_33__28_ <= r_n_33__28_;
      r_33__27_ <= r_n_33__27_;
      r_33__26_ <= r_n_33__26_;
      r_33__25_ <= r_n_33__25_;
      r_33__24_ <= r_n_33__24_;
      r_33__23_ <= r_n_33__23_;
      r_33__22_ <= r_n_33__22_;
      r_33__21_ <= r_n_33__21_;
      r_33__20_ <= r_n_33__20_;
      r_33__19_ <= r_n_33__19_;
      r_33__18_ <= r_n_33__18_;
      r_33__17_ <= r_n_33__17_;
      r_33__16_ <= r_n_33__16_;
      r_33__15_ <= r_n_33__15_;
      r_33__14_ <= r_n_33__14_;
      r_33__13_ <= r_n_33__13_;
      r_33__12_ <= r_n_33__12_;
      r_33__11_ <= r_n_33__11_;
      r_33__10_ <= r_n_33__10_;
      r_33__9_ <= r_n_33__9_;
      r_33__8_ <= r_n_33__8_;
      r_33__7_ <= r_n_33__7_;
      r_33__6_ <= r_n_33__6_;
      r_33__5_ <= r_n_33__5_;
      r_33__4_ <= r_n_33__4_;
      r_33__3_ <= r_n_33__3_;
      r_33__2_ <= r_n_33__2_;
      r_33__1_ <= r_n_33__1_;
      r_33__0_ <= r_n_33__0_;
    end 
    if(N3618) begin
      r_34__63_ <= r_n_34__63_;
      r_34__62_ <= r_n_34__62_;
      r_34__61_ <= r_n_34__61_;
      r_34__60_ <= r_n_34__60_;
      r_34__59_ <= r_n_34__59_;
      r_34__58_ <= r_n_34__58_;
      r_34__57_ <= r_n_34__57_;
      r_34__56_ <= r_n_34__56_;
      r_34__55_ <= r_n_34__55_;
      r_34__54_ <= r_n_34__54_;
      r_34__53_ <= r_n_34__53_;
      r_34__52_ <= r_n_34__52_;
      r_34__51_ <= r_n_34__51_;
      r_34__50_ <= r_n_34__50_;
      r_34__49_ <= r_n_34__49_;
      r_34__48_ <= r_n_34__48_;
      r_34__47_ <= r_n_34__47_;
      r_34__46_ <= r_n_34__46_;
      r_34__45_ <= r_n_34__45_;
      r_34__44_ <= r_n_34__44_;
      r_34__43_ <= r_n_34__43_;
      r_34__42_ <= r_n_34__42_;
      r_34__41_ <= r_n_34__41_;
      r_34__40_ <= r_n_34__40_;
      r_34__39_ <= r_n_34__39_;
      r_34__38_ <= r_n_34__38_;
      r_34__37_ <= r_n_34__37_;
      r_34__36_ <= r_n_34__36_;
      r_34__35_ <= r_n_34__35_;
      r_34__34_ <= r_n_34__34_;
      r_34__33_ <= r_n_34__33_;
      r_34__32_ <= r_n_34__32_;
      r_34__31_ <= r_n_34__31_;
      r_34__30_ <= r_n_34__30_;
      r_34__29_ <= r_n_34__29_;
      r_34__28_ <= r_n_34__28_;
      r_34__27_ <= r_n_34__27_;
      r_34__26_ <= r_n_34__26_;
      r_34__25_ <= r_n_34__25_;
      r_34__24_ <= r_n_34__24_;
      r_34__23_ <= r_n_34__23_;
      r_34__22_ <= r_n_34__22_;
      r_34__21_ <= r_n_34__21_;
      r_34__20_ <= r_n_34__20_;
      r_34__19_ <= r_n_34__19_;
      r_34__18_ <= r_n_34__18_;
      r_34__17_ <= r_n_34__17_;
      r_34__16_ <= r_n_34__16_;
      r_34__15_ <= r_n_34__15_;
      r_34__14_ <= r_n_34__14_;
      r_34__13_ <= r_n_34__13_;
      r_34__12_ <= r_n_34__12_;
      r_34__11_ <= r_n_34__11_;
      r_34__10_ <= r_n_34__10_;
      r_34__9_ <= r_n_34__9_;
      r_34__8_ <= r_n_34__8_;
      r_34__7_ <= r_n_34__7_;
      r_34__6_ <= r_n_34__6_;
      r_34__5_ <= r_n_34__5_;
      r_34__4_ <= r_n_34__4_;
      r_34__3_ <= r_n_34__3_;
      r_34__2_ <= r_n_34__2_;
      r_34__1_ <= r_n_34__1_;
      r_34__0_ <= r_n_34__0_;
    end 
    if(N3619) begin
      r_35__63_ <= r_n_35__63_;
      r_35__62_ <= r_n_35__62_;
      r_35__61_ <= r_n_35__61_;
      r_35__60_ <= r_n_35__60_;
      r_35__59_ <= r_n_35__59_;
      r_35__58_ <= r_n_35__58_;
      r_35__57_ <= r_n_35__57_;
      r_35__56_ <= r_n_35__56_;
      r_35__55_ <= r_n_35__55_;
      r_35__54_ <= r_n_35__54_;
      r_35__53_ <= r_n_35__53_;
      r_35__52_ <= r_n_35__52_;
      r_35__51_ <= r_n_35__51_;
      r_35__50_ <= r_n_35__50_;
      r_35__49_ <= r_n_35__49_;
      r_35__48_ <= r_n_35__48_;
      r_35__47_ <= r_n_35__47_;
      r_35__46_ <= r_n_35__46_;
      r_35__45_ <= r_n_35__45_;
      r_35__44_ <= r_n_35__44_;
      r_35__43_ <= r_n_35__43_;
      r_35__42_ <= r_n_35__42_;
      r_35__41_ <= r_n_35__41_;
      r_35__40_ <= r_n_35__40_;
      r_35__39_ <= r_n_35__39_;
      r_35__38_ <= r_n_35__38_;
      r_35__37_ <= r_n_35__37_;
      r_35__36_ <= r_n_35__36_;
      r_35__35_ <= r_n_35__35_;
      r_35__34_ <= r_n_35__34_;
      r_35__33_ <= r_n_35__33_;
      r_35__32_ <= r_n_35__32_;
      r_35__31_ <= r_n_35__31_;
      r_35__30_ <= r_n_35__30_;
      r_35__29_ <= r_n_35__29_;
      r_35__28_ <= r_n_35__28_;
      r_35__27_ <= r_n_35__27_;
      r_35__26_ <= r_n_35__26_;
      r_35__25_ <= r_n_35__25_;
      r_35__24_ <= r_n_35__24_;
      r_35__23_ <= r_n_35__23_;
      r_35__22_ <= r_n_35__22_;
      r_35__21_ <= r_n_35__21_;
      r_35__20_ <= r_n_35__20_;
      r_35__19_ <= r_n_35__19_;
      r_35__18_ <= r_n_35__18_;
      r_35__17_ <= r_n_35__17_;
      r_35__16_ <= r_n_35__16_;
      r_35__15_ <= r_n_35__15_;
      r_35__14_ <= r_n_35__14_;
      r_35__13_ <= r_n_35__13_;
      r_35__12_ <= r_n_35__12_;
      r_35__11_ <= r_n_35__11_;
      r_35__10_ <= r_n_35__10_;
      r_35__9_ <= r_n_35__9_;
      r_35__8_ <= r_n_35__8_;
      r_35__7_ <= r_n_35__7_;
      r_35__6_ <= r_n_35__6_;
      r_35__5_ <= r_n_35__5_;
      r_35__4_ <= r_n_35__4_;
      r_35__3_ <= r_n_35__3_;
      r_35__2_ <= r_n_35__2_;
      r_35__1_ <= r_n_35__1_;
      r_35__0_ <= r_n_35__0_;
    end 
    if(N3620) begin
      r_36__63_ <= r_n_36__63_;
      r_36__62_ <= r_n_36__62_;
      r_36__61_ <= r_n_36__61_;
      r_36__60_ <= r_n_36__60_;
      r_36__59_ <= r_n_36__59_;
      r_36__58_ <= r_n_36__58_;
      r_36__57_ <= r_n_36__57_;
      r_36__56_ <= r_n_36__56_;
      r_36__55_ <= r_n_36__55_;
      r_36__54_ <= r_n_36__54_;
      r_36__53_ <= r_n_36__53_;
      r_36__52_ <= r_n_36__52_;
      r_36__51_ <= r_n_36__51_;
      r_36__50_ <= r_n_36__50_;
      r_36__49_ <= r_n_36__49_;
      r_36__48_ <= r_n_36__48_;
      r_36__47_ <= r_n_36__47_;
      r_36__46_ <= r_n_36__46_;
      r_36__45_ <= r_n_36__45_;
      r_36__44_ <= r_n_36__44_;
      r_36__43_ <= r_n_36__43_;
      r_36__42_ <= r_n_36__42_;
      r_36__41_ <= r_n_36__41_;
      r_36__40_ <= r_n_36__40_;
      r_36__39_ <= r_n_36__39_;
      r_36__38_ <= r_n_36__38_;
      r_36__37_ <= r_n_36__37_;
      r_36__36_ <= r_n_36__36_;
      r_36__35_ <= r_n_36__35_;
      r_36__34_ <= r_n_36__34_;
      r_36__33_ <= r_n_36__33_;
      r_36__32_ <= r_n_36__32_;
      r_36__31_ <= r_n_36__31_;
      r_36__30_ <= r_n_36__30_;
      r_36__29_ <= r_n_36__29_;
      r_36__28_ <= r_n_36__28_;
      r_36__27_ <= r_n_36__27_;
      r_36__26_ <= r_n_36__26_;
      r_36__25_ <= r_n_36__25_;
      r_36__24_ <= r_n_36__24_;
      r_36__23_ <= r_n_36__23_;
      r_36__22_ <= r_n_36__22_;
      r_36__21_ <= r_n_36__21_;
      r_36__20_ <= r_n_36__20_;
      r_36__19_ <= r_n_36__19_;
      r_36__18_ <= r_n_36__18_;
      r_36__17_ <= r_n_36__17_;
      r_36__16_ <= r_n_36__16_;
      r_36__15_ <= r_n_36__15_;
      r_36__14_ <= r_n_36__14_;
      r_36__13_ <= r_n_36__13_;
      r_36__12_ <= r_n_36__12_;
      r_36__11_ <= r_n_36__11_;
      r_36__10_ <= r_n_36__10_;
      r_36__9_ <= r_n_36__9_;
      r_36__8_ <= r_n_36__8_;
      r_36__7_ <= r_n_36__7_;
      r_36__6_ <= r_n_36__6_;
      r_36__5_ <= r_n_36__5_;
      r_36__4_ <= r_n_36__4_;
      r_36__3_ <= r_n_36__3_;
      r_36__2_ <= r_n_36__2_;
      r_36__1_ <= r_n_36__1_;
      r_36__0_ <= r_n_36__0_;
    end 
    if(N3621) begin
      r_37__63_ <= r_n_37__63_;
      r_37__62_ <= r_n_37__62_;
      r_37__61_ <= r_n_37__61_;
      r_37__60_ <= r_n_37__60_;
      r_37__59_ <= r_n_37__59_;
      r_37__58_ <= r_n_37__58_;
      r_37__57_ <= r_n_37__57_;
      r_37__56_ <= r_n_37__56_;
      r_37__55_ <= r_n_37__55_;
      r_37__54_ <= r_n_37__54_;
      r_37__53_ <= r_n_37__53_;
      r_37__52_ <= r_n_37__52_;
      r_37__51_ <= r_n_37__51_;
      r_37__50_ <= r_n_37__50_;
      r_37__49_ <= r_n_37__49_;
      r_37__48_ <= r_n_37__48_;
      r_37__47_ <= r_n_37__47_;
      r_37__46_ <= r_n_37__46_;
      r_37__45_ <= r_n_37__45_;
      r_37__44_ <= r_n_37__44_;
      r_37__43_ <= r_n_37__43_;
      r_37__42_ <= r_n_37__42_;
      r_37__41_ <= r_n_37__41_;
      r_37__40_ <= r_n_37__40_;
      r_37__39_ <= r_n_37__39_;
      r_37__38_ <= r_n_37__38_;
      r_37__37_ <= r_n_37__37_;
      r_37__36_ <= r_n_37__36_;
      r_37__35_ <= r_n_37__35_;
      r_37__34_ <= r_n_37__34_;
      r_37__33_ <= r_n_37__33_;
      r_37__32_ <= r_n_37__32_;
      r_37__31_ <= r_n_37__31_;
      r_37__30_ <= r_n_37__30_;
      r_37__29_ <= r_n_37__29_;
      r_37__28_ <= r_n_37__28_;
      r_37__27_ <= r_n_37__27_;
      r_37__26_ <= r_n_37__26_;
      r_37__25_ <= r_n_37__25_;
      r_37__24_ <= r_n_37__24_;
      r_37__23_ <= r_n_37__23_;
      r_37__22_ <= r_n_37__22_;
      r_37__21_ <= r_n_37__21_;
      r_37__20_ <= r_n_37__20_;
      r_37__19_ <= r_n_37__19_;
      r_37__18_ <= r_n_37__18_;
      r_37__17_ <= r_n_37__17_;
      r_37__16_ <= r_n_37__16_;
      r_37__15_ <= r_n_37__15_;
      r_37__14_ <= r_n_37__14_;
      r_37__13_ <= r_n_37__13_;
      r_37__12_ <= r_n_37__12_;
      r_37__11_ <= r_n_37__11_;
      r_37__10_ <= r_n_37__10_;
      r_37__9_ <= r_n_37__9_;
      r_37__8_ <= r_n_37__8_;
      r_37__7_ <= r_n_37__7_;
      r_37__6_ <= r_n_37__6_;
      r_37__5_ <= r_n_37__5_;
      r_37__4_ <= r_n_37__4_;
      r_37__3_ <= r_n_37__3_;
      r_37__2_ <= r_n_37__2_;
      r_37__1_ <= r_n_37__1_;
      r_37__0_ <= r_n_37__0_;
    end 
    if(N3622) begin
      r_38__63_ <= r_n_38__63_;
      r_38__62_ <= r_n_38__62_;
      r_38__61_ <= r_n_38__61_;
      r_38__60_ <= r_n_38__60_;
      r_38__59_ <= r_n_38__59_;
      r_38__58_ <= r_n_38__58_;
      r_38__57_ <= r_n_38__57_;
      r_38__56_ <= r_n_38__56_;
      r_38__55_ <= r_n_38__55_;
      r_38__54_ <= r_n_38__54_;
      r_38__53_ <= r_n_38__53_;
      r_38__52_ <= r_n_38__52_;
      r_38__51_ <= r_n_38__51_;
      r_38__50_ <= r_n_38__50_;
      r_38__49_ <= r_n_38__49_;
      r_38__48_ <= r_n_38__48_;
      r_38__47_ <= r_n_38__47_;
      r_38__46_ <= r_n_38__46_;
      r_38__45_ <= r_n_38__45_;
      r_38__44_ <= r_n_38__44_;
      r_38__43_ <= r_n_38__43_;
      r_38__42_ <= r_n_38__42_;
      r_38__41_ <= r_n_38__41_;
      r_38__40_ <= r_n_38__40_;
      r_38__39_ <= r_n_38__39_;
      r_38__38_ <= r_n_38__38_;
      r_38__37_ <= r_n_38__37_;
      r_38__36_ <= r_n_38__36_;
      r_38__35_ <= r_n_38__35_;
      r_38__34_ <= r_n_38__34_;
      r_38__33_ <= r_n_38__33_;
      r_38__32_ <= r_n_38__32_;
      r_38__31_ <= r_n_38__31_;
      r_38__30_ <= r_n_38__30_;
      r_38__29_ <= r_n_38__29_;
      r_38__28_ <= r_n_38__28_;
      r_38__27_ <= r_n_38__27_;
      r_38__26_ <= r_n_38__26_;
      r_38__25_ <= r_n_38__25_;
      r_38__24_ <= r_n_38__24_;
      r_38__23_ <= r_n_38__23_;
      r_38__22_ <= r_n_38__22_;
      r_38__21_ <= r_n_38__21_;
      r_38__20_ <= r_n_38__20_;
      r_38__19_ <= r_n_38__19_;
      r_38__18_ <= r_n_38__18_;
      r_38__17_ <= r_n_38__17_;
      r_38__16_ <= r_n_38__16_;
      r_38__15_ <= r_n_38__15_;
      r_38__14_ <= r_n_38__14_;
      r_38__13_ <= r_n_38__13_;
      r_38__12_ <= r_n_38__12_;
      r_38__11_ <= r_n_38__11_;
      r_38__10_ <= r_n_38__10_;
      r_38__9_ <= r_n_38__9_;
      r_38__8_ <= r_n_38__8_;
      r_38__7_ <= r_n_38__7_;
      r_38__6_ <= r_n_38__6_;
      r_38__5_ <= r_n_38__5_;
      r_38__4_ <= r_n_38__4_;
      r_38__3_ <= r_n_38__3_;
      r_38__2_ <= r_n_38__2_;
      r_38__1_ <= r_n_38__1_;
      r_38__0_ <= r_n_38__0_;
    end 
    if(N3623) begin
      r_39__63_ <= r_n_39__63_;
      r_39__62_ <= r_n_39__62_;
      r_39__61_ <= r_n_39__61_;
      r_39__60_ <= r_n_39__60_;
      r_39__59_ <= r_n_39__59_;
      r_39__58_ <= r_n_39__58_;
      r_39__57_ <= r_n_39__57_;
      r_39__56_ <= r_n_39__56_;
      r_39__55_ <= r_n_39__55_;
      r_39__54_ <= r_n_39__54_;
      r_39__53_ <= r_n_39__53_;
      r_39__52_ <= r_n_39__52_;
      r_39__51_ <= r_n_39__51_;
      r_39__50_ <= r_n_39__50_;
      r_39__49_ <= r_n_39__49_;
      r_39__48_ <= r_n_39__48_;
      r_39__47_ <= r_n_39__47_;
      r_39__46_ <= r_n_39__46_;
      r_39__45_ <= r_n_39__45_;
      r_39__44_ <= r_n_39__44_;
      r_39__43_ <= r_n_39__43_;
      r_39__42_ <= r_n_39__42_;
      r_39__41_ <= r_n_39__41_;
      r_39__40_ <= r_n_39__40_;
      r_39__39_ <= r_n_39__39_;
      r_39__38_ <= r_n_39__38_;
      r_39__37_ <= r_n_39__37_;
      r_39__36_ <= r_n_39__36_;
      r_39__35_ <= r_n_39__35_;
      r_39__34_ <= r_n_39__34_;
      r_39__33_ <= r_n_39__33_;
      r_39__32_ <= r_n_39__32_;
      r_39__31_ <= r_n_39__31_;
      r_39__30_ <= r_n_39__30_;
      r_39__29_ <= r_n_39__29_;
      r_39__28_ <= r_n_39__28_;
      r_39__27_ <= r_n_39__27_;
      r_39__26_ <= r_n_39__26_;
      r_39__25_ <= r_n_39__25_;
      r_39__24_ <= r_n_39__24_;
      r_39__23_ <= r_n_39__23_;
      r_39__22_ <= r_n_39__22_;
      r_39__21_ <= r_n_39__21_;
      r_39__20_ <= r_n_39__20_;
      r_39__19_ <= r_n_39__19_;
      r_39__18_ <= r_n_39__18_;
      r_39__17_ <= r_n_39__17_;
      r_39__16_ <= r_n_39__16_;
      r_39__15_ <= r_n_39__15_;
      r_39__14_ <= r_n_39__14_;
      r_39__13_ <= r_n_39__13_;
      r_39__12_ <= r_n_39__12_;
      r_39__11_ <= r_n_39__11_;
      r_39__10_ <= r_n_39__10_;
      r_39__9_ <= r_n_39__9_;
      r_39__8_ <= r_n_39__8_;
      r_39__7_ <= r_n_39__7_;
      r_39__6_ <= r_n_39__6_;
      r_39__5_ <= r_n_39__5_;
      r_39__4_ <= r_n_39__4_;
      r_39__3_ <= r_n_39__3_;
      r_39__2_ <= r_n_39__2_;
      r_39__1_ <= r_n_39__1_;
      r_39__0_ <= r_n_39__0_;
    end 
    if(N3624) begin
      r_40__63_ <= r_n_40__63_;
      r_40__62_ <= r_n_40__62_;
      r_40__61_ <= r_n_40__61_;
      r_40__60_ <= r_n_40__60_;
      r_40__59_ <= r_n_40__59_;
      r_40__58_ <= r_n_40__58_;
      r_40__57_ <= r_n_40__57_;
      r_40__56_ <= r_n_40__56_;
      r_40__55_ <= r_n_40__55_;
      r_40__54_ <= r_n_40__54_;
      r_40__53_ <= r_n_40__53_;
      r_40__52_ <= r_n_40__52_;
      r_40__51_ <= r_n_40__51_;
      r_40__50_ <= r_n_40__50_;
      r_40__49_ <= r_n_40__49_;
      r_40__48_ <= r_n_40__48_;
      r_40__47_ <= r_n_40__47_;
      r_40__46_ <= r_n_40__46_;
      r_40__45_ <= r_n_40__45_;
      r_40__44_ <= r_n_40__44_;
      r_40__43_ <= r_n_40__43_;
      r_40__42_ <= r_n_40__42_;
      r_40__41_ <= r_n_40__41_;
      r_40__40_ <= r_n_40__40_;
      r_40__39_ <= r_n_40__39_;
      r_40__38_ <= r_n_40__38_;
      r_40__37_ <= r_n_40__37_;
      r_40__36_ <= r_n_40__36_;
      r_40__35_ <= r_n_40__35_;
      r_40__34_ <= r_n_40__34_;
      r_40__33_ <= r_n_40__33_;
      r_40__32_ <= r_n_40__32_;
      r_40__31_ <= r_n_40__31_;
      r_40__30_ <= r_n_40__30_;
      r_40__29_ <= r_n_40__29_;
      r_40__28_ <= r_n_40__28_;
      r_40__27_ <= r_n_40__27_;
      r_40__26_ <= r_n_40__26_;
      r_40__25_ <= r_n_40__25_;
      r_40__24_ <= r_n_40__24_;
      r_40__23_ <= r_n_40__23_;
      r_40__22_ <= r_n_40__22_;
      r_40__21_ <= r_n_40__21_;
      r_40__20_ <= r_n_40__20_;
      r_40__19_ <= r_n_40__19_;
      r_40__18_ <= r_n_40__18_;
      r_40__17_ <= r_n_40__17_;
      r_40__16_ <= r_n_40__16_;
      r_40__15_ <= r_n_40__15_;
      r_40__14_ <= r_n_40__14_;
      r_40__13_ <= r_n_40__13_;
      r_40__12_ <= r_n_40__12_;
      r_40__11_ <= r_n_40__11_;
      r_40__10_ <= r_n_40__10_;
      r_40__9_ <= r_n_40__9_;
      r_40__8_ <= r_n_40__8_;
      r_40__7_ <= r_n_40__7_;
      r_40__6_ <= r_n_40__6_;
      r_40__5_ <= r_n_40__5_;
      r_40__4_ <= r_n_40__4_;
      r_40__3_ <= r_n_40__3_;
      r_40__2_ <= r_n_40__2_;
      r_40__1_ <= r_n_40__1_;
      r_40__0_ <= r_n_40__0_;
    end 
    if(N3625) begin
      r_41__63_ <= r_n_41__63_;
      r_41__62_ <= r_n_41__62_;
      r_41__61_ <= r_n_41__61_;
      r_41__60_ <= r_n_41__60_;
      r_41__59_ <= r_n_41__59_;
      r_41__58_ <= r_n_41__58_;
      r_41__57_ <= r_n_41__57_;
      r_41__56_ <= r_n_41__56_;
      r_41__55_ <= r_n_41__55_;
      r_41__54_ <= r_n_41__54_;
      r_41__53_ <= r_n_41__53_;
      r_41__52_ <= r_n_41__52_;
      r_41__51_ <= r_n_41__51_;
      r_41__50_ <= r_n_41__50_;
      r_41__49_ <= r_n_41__49_;
      r_41__48_ <= r_n_41__48_;
      r_41__47_ <= r_n_41__47_;
      r_41__46_ <= r_n_41__46_;
      r_41__45_ <= r_n_41__45_;
      r_41__44_ <= r_n_41__44_;
      r_41__43_ <= r_n_41__43_;
      r_41__42_ <= r_n_41__42_;
      r_41__41_ <= r_n_41__41_;
      r_41__40_ <= r_n_41__40_;
      r_41__39_ <= r_n_41__39_;
      r_41__38_ <= r_n_41__38_;
      r_41__37_ <= r_n_41__37_;
      r_41__36_ <= r_n_41__36_;
      r_41__35_ <= r_n_41__35_;
      r_41__34_ <= r_n_41__34_;
      r_41__33_ <= r_n_41__33_;
      r_41__32_ <= r_n_41__32_;
      r_41__31_ <= r_n_41__31_;
      r_41__30_ <= r_n_41__30_;
      r_41__29_ <= r_n_41__29_;
      r_41__28_ <= r_n_41__28_;
      r_41__27_ <= r_n_41__27_;
      r_41__26_ <= r_n_41__26_;
      r_41__25_ <= r_n_41__25_;
      r_41__24_ <= r_n_41__24_;
      r_41__23_ <= r_n_41__23_;
      r_41__22_ <= r_n_41__22_;
      r_41__21_ <= r_n_41__21_;
      r_41__20_ <= r_n_41__20_;
      r_41__19_ <= r_n_41__19_;
      r_41__18_ <= r_n_41__18_;
      r_41__17_ <= r_n_41__17_;
      r_41__16_ <= r_n_41__16_;
      r_41__15_ <= r_n_41__15_;
      r_41__14_ <= r_n_41__14_;
      r_41__13_ <= r_n_41__13_;
      r_41__12_ <= r_n_41__12_;
      r_41__11_ <= r_n_41__11_;
      r_41__10_ <= r_n_41__10_;
      r_41__9_ <= r_n_41__9_;
      r_41__8_ <= r_n_41__8_;
      r_41__7_ <= r_n_41__7_;
      r_41__6_ <= r_n_41__6_;
      r_41__5_ <= r_n_41__5_;
      r_41__4_ <= r_n_41__4_;
      r_41__3_ <= r_n_41__3_;
      r_41__2_ <= r_n_41__2_;
      r_41__1_ <= r_n_41__1_;
      r_41__0_ <= r_n_41__0_;
    end 
    if(N3626) begin
      r_42__63_ <= r_n_42__63_;
      r_42__62_ <= r_n_42__62_;
      r_42__61_ <= r_n_42__61_;
      r_42__60_ <= r_n_42__60_;
      r_42__59_ <= r_n_42__59_;
      r_42__58_ <= r_n_42__58_;
      r_42__57_ <= r_n_42__57_;
      r_42__56_ <= r_n_42__56_;
      r_42__55_ <= r_n_42__55_;
      r_42__54_ <= r_n_42__54_;
      r_42__53_ <= r_n_42__53_;
      r_42__52_ <= r_n_42__52_;
      r_42__51_ <= r_n_42__51_;
      r_42__50_ <= r_n_42__50_;
      r_42__49_ <= r_n_42__49_;
      r_42__48_ <= r_n_42__48_;
      r_42__47_ <= r_n_42__47_;
      r_42__46_ <= r_n_42__46_;
      r_42__45_ <= r_n_42__45_;
      r_42__44_ <= r_n_42__44_;
      r_42__43_ <= r_n_42__43_;
      r_42__42_ <= r_n_42__42_;
      r_42__41_ <= r_n_42__41_;
      r_42__40_ <= r_n_42__40_;
      r_42__39_ <= r_n_42__39_;
      r_42__38_ <= r_n_42__38_;
      r_42__37_ <= r_n_42__37_;
      r_42__36_ <= r_n_42__36_;
      r_42__35_ <= r_n_42__35_;
      r_42__34_ <= r_n_42__34_;
      r_42__33_ <= r_n_42__33_;
      r_42__32_ <= r_n_42__32_;
      r_42__31_ <= r_n_42__31_;
      r_42__30_ <= r_n_42__30_;
      r_42__29_ <= r_n_42__29_;
      r_42__28_ <= r_n_42__28_;
      r_42__27_ <= r_n_42__27_;
      r_42__26_ <= r_n_42__26_;
      r_42__25_ <= r_n_42__25_;
      r_42__24_ <= r_n_42__24_;
      r_42__23_ <= r_n_42__23_;
      r_42__22_ <= r_n_42__22_;
      r_42__21_ <= r_n_42__21_;
      r_42__20_ <= r_n_42__20_;
      r_42__19_ <= r_n_42__19_;
      r_42__18_ <= r_n_42__18_;
      r_42__17_ <= r_n_42__17_;
      r_42__16_ <= r_n_42__16_;
      r_42__15_ <= r_n_42__15_;
      r_42__14_ <= r_n_42__14_;
      r_42__13_ <= r_n_42__13_;
      r_42__12_ <= r_n_42__12_;
      r_42__11_ <= r_n_42__11_;
      r_42__10_ <= r_n_42__10_;
      r_42__9_ <= r_n_42__9_;
      r_42__8_ <= r_n_42__8_;
      r_42__7_ <= r_n_42__7_;
      r_42__6_ <= r_n_42__6_;
      r_42__5_ <= r_n_42__5_;
      r_42__4_ <= r_n_42__4_;
      r_42__3_ <= r_n_42__3_;
      r_42__2_ <= r_n_42__2_;
      r_42__1_ <= r_n_42__1_;
      r_42__0_ <= r_n_42__0_;
    end 
    if(N3627) begin
      r_43__63_ <= r_n_43__63_;
      r_43__62_ <= r_n_43__62_;
      r_43__61_ <= r_n_43__61_;
      r_43__60_ <= r_n_43__60_;
      r_43__59_ <= r_n_43__59_;
      r_43__58_ <= r_n_43__58_;
      r_43__57_ <= r_n_43__57_;
      r_43__56_ <= r_n_43__56_;
      r_43__55_ <= r_n_43__55_;
      r_43__54_ <= r_n_43__54_;
      r_43__53_ <= r_n_43__53_;
      r_43__52_ <= r_n_43__52_;
      r_43__51_ <= r_n_43__51_;
      r_43__50_ <= r_n_43__50_;
      r_43__49_ <= r_n_43__49_;
      r_43__48_ <= r_n_43__48_;
      r_43__47_ <= r_n_43__47_;
      r_43__46_ <= r_n_43__46_;
      r_43__45_ <= r_n_43__45_;
      r_43__44_ <= r_n_43__44_;
      r_43__43_ <= r_n_43__43_;
      r_43__42_ <= r_n_43__42_;
      r_43__41_ <= r_n_43__41_;
      r_43__40_ <= r_n_43__40_;
      r_43__39_ <= r_n_43__39_;
      r_43__38_ <= r_n_43__38_;
      r_43__37_ <= r_n_43__37_;
      r_43__36_ <= r_n_43__36_;
      r_43__35_ <= r_n_43__35_;
      r_43__34_ <= r_n_43__34_;
      r_43__33_ <= r_n_43__33_;
      r_43__32_ <= r_n_43__32_;
      r_43__31_ <= r_n_43__31_;
      r_43__30_ <= r_n_43__30_;
      r_43__29_ <= r_n_43__29_;
      r_43__28_ <= r_n_43__28_;
      r_43__27_ <= r_n_43__27_;
      r_43__26_ <= r_n_43__26_;
      r_43__25_ <= r_n_43__25_;
      r_43__24_ <= r_n_43__24_;
      r_43__23_ <= r_n_43__23_;
      r_43__22_ <= r_n_43__22_;
      r_43__21_ <= r_n_43__21_;
      r_43__20_ <= r_n_43__20_;
      r_43__19_ <= r_n_43__19_;
      r_43__18_ <= r_n_43__18_;
      r_43__17_ <= r_n_43__17_;
      r_43__16_ <= r_n_43__16_;
      r_43__15_ <= r_n_43__15_;
      r_43__14_ <= r_n_43__14_;
      r_43__13_ <= r_n_43__13_;
      r_43__12_ <= r_n_43__12_;
      r_43__11_ <= r_n_43__11_;
      r_43__10_ <= r_n_43__10_;
      r_43__9_ <= r_n_43__9_;
      r_43__8_ <= r_n_43__8_;
      r_43__7_ <= r_n_43__7_;
      r_43__6_ <= r_n_43__6_;
      r_43__5_ <= r_n_43__5_;
      r_43__4_ <= r_n_43__4_;
      r_43__3_ <= r_n_43__3_;
      r_43__2_ <= r_n_43__2_;
      r_43__1_ <= r_n_43__1_;
      r_43__0_ <= r_n_43__0_;
    end 
    if(N3628) begin
      r_44__63_ <= r_n_44__63_;
      r_44__62_ <= r_n_44__62_;
      r_44__61_ <= r_n_44__61_;
      r_44__60_ <= r_n_44__60_;
      r_44__59_ <= r_n_44__59_;
      r_44__58_ <= r_n_44__58_;
      r_44__57_ <= r_n_44__57_;
      r_44__56_ <= r_n_44__56_;
      r_44__55_ <= r_n_44__55_;
      r_44__54_ <= r_n_44__54_;
      r_44__53_ <= r_n_44__53_;
      r_44__52_ <= r_n_44__52_;
      r_44__51_ <= r_n_44__51_;
      r_44__50_ <= r_n_44__50_;
      r_44__49_ <= r_n_44__49_;
      r_44__48_ <= r_n_44__48_;
      r_44__47_ <= r_n_44__47_;
      r_44__46_ <= r_n_44__46_;
      r_44__45_ <= r_n_44__45_;
      r_44__44_ <= r_n_44__44_;
      r_44__43_ <= r_n_44__43_;
      r_44__42_ <= r_n_44__42_;
      r_44__41_ <= r_n_44__41_;
      r_44__40_ <= r_n_44__40_;
      r_44__39_ <= r_n_44__39_;
      r_44__38_ <= r_n_44__38_;
      r_44__37_ <= r_n_44__37_;
      r_44__36_ <= r_n_44__36_;
      r_44__35_ <= r_n_44__35_;
      r_44__34_ <= r_n_44__34_;
      r_44__33_ <= r_n_44__33_;
      r_44__32_ <= r_n_44__32_;
      r_44__31_ <= r_n_44__31_;
      r_44__30_ <= r_n_44__30_;
      r_44__29_ <= r_n_44__29_;
      r_44__28_ <= r_n_44__28_;
      r_44__27_ <= r_n_44__27_;
      r_44__26_ <= r_n_44__26_;
      r_44__25_ <= r_n_44__25_;
      r_44__24_ <= r_n_44__24_;
      r_44__23_ <= r_n_44__23_;
      r_44__22_ <= r_n_44__22_;
      r_44__21_ <= r_n_44__21_;
      r_44__20_ <= r_n_44__20_;
      r_44__19_ <= r_n_44__19_;
      r_44__18_ <= r_n_44__18_;
      r_44__17_ <= r_n_44__17_;
      r_44__16_ <= r_n_44__16_;
      r_44__15_ <= r_n_44__15_;
      r_44__14_ <= r_n_44__14_;
      r_44__13_ <= r_n_44__13_;
      r_44__12_ <= r_n_44__12_;
      r_44__11_ <= r_n_44__11_;
      r_44__10_ <= r_n_44__10_;
      r_44__9_ <= r_n_44__9_;
      r_44__8_ <= r_n_44__8_;
      r_44__7_ <= r_n_44__7_;
      r_44__6_ <= r_n_44__6_;
      r_44__5_ <= r_n_44__5_;
      r_44__4_ <= r_n_44__4_;
      r_44__3_ <= r_n_44__3_;
      r_44__2_ <= r_n_44__2_;
      r_44__1_ <= r_n_44__1_;
      r_44__0_ <= r_n_44__0_;
    end 
    if(N3629) begin
      r_45__63_ <= r_n_45__63_;
      r_45__62_ <= r_n_45__62_;
      r_45__61_ <= r_n_45__61_;
      r_45__60_ <= r_n_45__60_;
      r_45__59_ <= r_n_45__59_;
      r_45__58_ <= r_n_45__58_;
      r_45__57_ <= r_n_45__57_;
      r_45__56_ <= r_n_45__56_;
      r_45__55_ <= r_n_45__55_;
      r_45__54_ <= r_n_45__54_;
      r_45__53_ <= r_n_45__53_;
      r_45__52_ <= r_n_45__52_;
      r_45__51_ <= r_n_45__51_;
      r_45__50_ <= r_n_45__50_;
      r_45__49_ <= r_n_45__49_;
      r_45__48_ <= r_n_45__48_;
      r_45__47_ <= r_n_45__47_;
      r_45__46_ <= r_n_45__46_;
      r_45__45_ <= r_n_45__45_;
      r_45__44_ <= r_n_45__44_;
      r_45__43_ <= r_n_45__43_;
      r_45__42_ <= r_n_45__42_;
      r_45__41_ <= r_n_45__41_;
      r_45__40_ <= r_n_45__40_;
      r_45__39_ <= r_n_45__39_;
      r_45__38_ <= r_n_45__38_;
      r_45__37_ <= r_n_45__37_;
      r_45__36_ <= r_n_45__36_;
      r_45__35_ <= r_n_45__35_;
      r_45__34_ <= r_n_45__34_;
      r_45__33_ <= r_n_45__33_;
      r_45__32_ <= r_n_45__32_;
      r_45__31_ <= r_n_45__31_;
      r_45__30_ <= r_n_45__30_;
      r_45__29_ <= r_n_45__29_;
      r_45__28_ <= r_n_45__28_;
      r_45__27_ <= r_n_45__27_;
      r_45__26_ <= r_n_45__26_;
      r_45__25_ <= r_n_45__25_;
      r_45__24_ <= r_n_45__24_;
      r_45__23_ <= r_n_45__23_;
      r_45__22_ <= r_n_45__22_;
      r_45__21_ <= r_n_45__21_;
      r_45__20_ <= r_n_45__20_;
      r_45__19_ <= r_n_45__19_;
      r_45__18_ <= r_n_45__18_;
      r_45__17_ <= r_n_45__17_;
      r_45__16_ <= r_n_45__16_;
      r_45__15_ <= r_n_45__15_;
      r_45__14_ <= r_n_45__14_;
      r_45__13_ <= r_n_45__13_;
      r_45__12_ <= r_n_45__12_;
      r_45__11_ <= r_n_45__11_;
      r_45__10_ <= r_n_45__10_;
      r_45__9_ <= r_n_45__9_;
      r_45__8_ <= r_n_45__8_;
      r_45__7_ <= r_n_45__7_;
      r_45__6_ <= r_n_45__6_;
      r_45__5_ <= r_n_45__5_;
      r_45__4_ <= r_n_45__4_;
      r_45__3_ <= r_n_45__3_;
      r_45__2_ <= r_n_45__2_;
      r_45__1_ <= r_n_45__1_;
      r_45__0_ <= r_n_45__0_;
    end 
    if(N3630) begin
      r_46__63_ <= r_n_46__63_;
      r_46__62_ <= r_n_46__62_;
      r_46__61_ <= r_n_46__61_;
      r_46__60_ <= r_n_46__60_;
      r_46__59_ <= r_n_46__59_;
      r_46__58_ <= r_n_46__58_;
      r_46__57_ <= r_n_46__57_;
      r_46__56_ <= r_n_46__56_;
      r_46__55_ <= r_n_46__55_;
      r_46__54_ <= r_n_46__54_;
      r_46__53_ <= r_n_46__53_;
      r_46__52_ <= r_n_46__52_;
      r_46__51_ <= r_n_46__51_;
      r_46__50_ <= r_n_46__50_;
      r_46__49_ <= r_n_46__49_;
      r_46__48_ <= r_n_46__48_;
      r_46__47_ <= r_n_46__47_;
      r_46__46_ <= r_n_46__46_;
      r_46__45_ <= r_n_46__45_;
      r_46__44_ <= r_n_46__44_;
      r_46__43_ <= r_n_46__43_;
      r_46__42_ <= r_n_46__42_;
      r_46__41_ <= r_n_46__41_;
      r_46__40_ <= r_n_46__40_;
      r_46__39_ <= r_n_46__39_;
      r_46__38_ <= r_n_46__38_;
      r_46__37_ <= r_n_46__37_;
      r_46__36_ <= r_n_46__36_;
      r_46__35_ <= r_n_46__35_;
      r_46__34_ <= r_n_46__34_;
      r_46__33_ <= r_n_46__33_;
      r_46__32_ <= r_n_46__32_;
      r_46__31_ <= r_n_46__31_;
      r_46__30_ <= r_n_46__30_;
      r_46__29_ <= r_n_46__29_;
      r_46__28_ <= r_n_46__28_;
      r_46__27_ <= r_n_46__27_;
      r_46__26_ <= r_n_46__26_;
      r_46__25_ <= r_n_46__25_;
      r_46__24_ <= r_n_46__24_;
      r_46__23_ <= r_n_46__23_;
      r_46__22_ <= r_n_46__22_;
      r_46__21_ <= r_n_46__21_;
      r_46__20_ <= r_n_46__20_;
      r_46__19_ <= r_n_46__19_;
      r_46__18_ <= r_n_46__18_;
      r_46__17_ <= r_n_46__17_;
      r_46__16_ <= r_n_46__16_;
      r_46__15_ <= r_n_46__15_;
      r_46__14_ <= r_n_46__14_;
      r_46__13_ <= r_n_46__13_;
      r_46__12_ <= r_n_46__12_;
      r_46__11_ <= r_n_46__11_;
      r_46__10_ <= r_n_46__10_;
      r_46__9_ <= r_n_46__9_;
      r_46__8_ <= r_n_46__8_;
      r_46__7_ <= r_n_46__7_;
      r_46__6_ <= r_n_46__6_;
      r_46__5_ <= r_n_46__5_;
      r_46__4_ <= r_n_46__4_;
      r_46__3_ <= r_n_46__3_;
      r_46__2_ <= r_n_46__2_;
      r_46__1_ <= r_n_46__1_;
      r_46__0_ <= r_n_46__0_;
    end 
    if(N3631) begin
      r_47__63_ <= r_n_47__63_;
      r_47__62_ <= r_n_47__62_;
      r_47__61_ <= r_n_47__61_;
      r_47__60_ <= r_n_47__60_;
      r_47__59_ <= r_n_47__59_;
      r_47__58_ <= r_n_47__58_;
      r_47__57_ <= r_n_47__57_;
      r_47__56_ <= r_n_47__56_;
      r_47__55_ <= r_n_47__55_;
      r_47__54_ <= r_n_47__54_;
      r_47__53_ <= r_n_47__53_;
      r_47__52_ <= r_n_47__52_;
      r_47__51_ <= r_n_47__51_;
      r_47__50_ <= r_n_47__50_;
      r_47__49_ <= r_n_47__49_;
      r_47__48_ <= r_n_47__48_;
      r_47__47_ <= r_n_47__47_;
      r_47__46_ <= r_n_47__46_;
      r_47__45_ <= r_n_47__45_;
      r_47__44_ <= r_n_47__44_;
      r_47__43_ <= r_n_47__43_;
      r_47__42_ <= r_n_47__42_;
      r_47__41_ <= r_n_47__41_;
      r_47__40_ <= r_n_47__40_;
      r_47__39_ <= r_n_47__39_;
      r_47__38_ <= r_n_47__38_;
      r_47__37_ <= r_n_47__37_;
      r_47__36_ <= r_n_47__36_;
      r_47__35_ <= r_n_47__35_;
      r_47__34_ <= r_n_47__34_;
      r_47__33_ <= r_n_47__33_;
      r_47__32_ <= r_n_47__32_;
      r_47__31_ <= r_n_47__31_;
      r_47__30_ <= r_n_47__30_;
      r_47__29_ <= r_n_47__29_;
      r_47__28_ <= r_n_47__28_;
      r_47__27_ <= r_n_47__27_;
      r_47__26_ <= r_n_47__26_;
      r_47__25_ <= r_n_47__25_;
      r_47__24_ <= r_n_47__24_;
      r_47__23_ <= r_n_47__23_;
      r_47__22_ <= r_n_47__22_;
      r_47__21_ <= r_n_47__21_;
      r_47__20_ <= r_n_47__20_;
      r_47__19_ <= r_n_47__19_;
      r_47__18_ <= r_n_47__18_;
      r_47__17_ <= r_n_47__17_;
      r_47__16_ <= r_n_47__16_;
      r_47__15_ <= r_n_47__15_;
      r_47__14_ <= r_n_47__14_;
      r_47__13_ <= r_n_47__13_;
      r_47__12_ <= r_n_47__12_;
      r_47__11_ <= r_n_47__11_;
      r_47__10_ <= r_n_47__10_;
      r_47__9_ <= r_n_47__9_;
      r_47__8_ <= r_n_47__8_;
      r_47__7_ <= r_n_47__7_;
      r_47__6_ <= r_n_47__6_;
      r_47__5_ <= r_n_47__5_;
      r_47__4_ <= r_n_47__4_;
      r_47__3_ <= r_n_47__3_;
      r_47__2_ <= r_n_47__2_;
      r_47__1_ <= r_n_47__1_;
      r_47__0_ <= r_n_47__0_;
    end 
    if(N3632) begin
      r_48__63_ <= r_n_48__63_;
      r_48__62_ <= r_n_48__62_;
      r_48__61_ <= r_n_48__61_;
      r_48__60_ <= r_n_48__60_;
      r_48__59_ <= r_n_48__59_;
      r_48__58_ <= r_n_48__58_;
      r_48__57_ <= r_n_48__57_;
      r_48__56_ <= r_n_48__56_;
      r_48__55_ <= r_n_48__55_;
      r_48__54_ <= r_n_48__54_;
      r_48__53_ <= r_n_48__53_;
      r_48__52_ <= r_n_48__52_;
      r_48__51_ <= r_n_48__51_;
      r_48__50_ <= r_n_48__50_;
      r_48__49_ <= r_n_48__49_;
      r_48__48_ <= r_n_48__48_;
      r_48__47_ <= r_n_48__47_;
      r_48__46_ <= r_n_48__46_;
      r_48__45_ <= r_n_48__45_;
      r_48__44_ <= r_n_48__44_;
      r_48__43_ <= r_n_48__43_;
      r_48__42_ <= r_n_48__42_;
      r_48__41_ <= r_n_48__41_;
      r_48__40_ <= r_n_48__40_;
      r_48__39_ <= r_n_48__39_;
      r_48__38_ <= r_n_48__38_;
      r_48__37_ <= r_n_48__37_;
      r_48__36_ <= r_n_48__36_;
      r_48__35_ <= r_n_48__35_;
      r_48__34_ <= r_n_48__34_;
      r_48__33_ <= r_n_48__33_;
      r_48__32_ <= r_n_48__32_;
      r_48__31_ <= r_n_48__31_;
      r_48__30_ <= r_n_48__30_;
      r_48__29_ <= r_n_48__29_;
      r_48__28_ <= r_n_48__28_;
      r_48__27_ <= r_n_48__27_;
      r_48__26_ <= r_n_48__26_;
      r_48__25_ <= r_n_48__25_;
      r_48__24_ <= r_n_48__24_;
      r_48__23_ <= r_n_48__23_;
      r_48__22_ <= r_n_48__22_;
      r_48__21_ <= r_n_48__21_;
      r_48__20_ <= r_n_48__20_;
      r_48__19_ <= r_n_48__19_;
      r_48__18_ <= r_n_48__18_;
      r_48__17_ <= r_n_48__17_;
      r_48__16_ <= r_n_48__16_;
      r_48__15_ <= r_n_48__15_;
      r_48__14_ <= r_n_48__14_;
      r_48__13_ <= r_n_48__13_;
      r_48__12_ <= r_n_48__12_;
      r_48__11_ <= r_n_48__11_;
      r_48__10_ <= r_n_48__10_;
      r_48__9_ <= r_n_48__9_;
      r_48__8_ <= r_n_48__8_;
      r_48__7_ <= r_n_48__7_;
      r_48__6_ <= r_n_48__6_;
      r_48__5_ <= r_n_48__5_;
      r_48__4_ <= r_n_48__4_;
      r_48__3_ <= r_n_48__3_;
      r_48__2_ <= r_n_48__2_;
      r_48__1_ <= r_n_48__1_;
      r_48__0_ <= r_n_48__0_;
    end 
    if(N3633) begin
      r_49__63_ <= r_n_49__63_;
      r_49__62_ <= r_n_49__62_;
      r_49__61_ <= r_n_49__61_;
      r_49__60_ <= r_n_49__60_;
      r_49__59_ <= r_n_49__59_;
      r_49__58_ <= r_n_49__58_;
      r_49__57_ <= r_n_49__57_;
      r_49__56_ <= r_n_49__56_;
      r_49__55_ <= r_n_49__55_;
      r_49__54_ <= r_n_49__54_;
      r_49__53_ <= r_n_49__53_;
      r_49__52_ <= r_n_49__52_;
      r_49__51_ <= r_n_49__51_;
      r_49__50_ <= r_n_49__50_;
      r_49__49_ <= r_n_49__49_;
      r_49__48_ <= r_n_49__48_;
      r_49__47_ <= r_n_49__47_;
      r_49__46_ <= r_n_49__46_;
      r_49__45_ <= r_n_49__45_;
      r_49__44_ <= r_n_49__44_;
      r_49__43_ <= r_n_49__43_;
      r_49__42_ <= r_n_49__42_;
      r_49__41_ <= r_n_49__41_;
      r_49__40_ <= r_n_49__40_;
      r_49__39_ <= r_n_49__39_;
      r_49__38_ <= r_n_49__38_;
      r_49__37_ <= r_n_49__37_;
      r_49__36_ <= r_n_49__36_;
      r_49__35_ <= r_n_49__35_;
      r_49__34_ <= r_n_49__34_;
      r_49__33_ <= r_n_49__33_;
      r_49__32_ <= r_n_49__32_;
      r_49__31_ <= r_n_49__31_;
      r_49__30_ <= r_n_49__30_;
      r_49__29_ <= r_n_49__29_;
      r_49__28_ <= r_n_49__28_;
      r_49__27_ <= r_n_49__27_;
      r_49__26_ <= r_n_49__26_;
      r_49__25_ <= r_n_49__25_;
      r_49__24_ <= r_n_49__24_;
      r_49__23_ <= r_n_49__23_;
      r_49__22_ <= r_n_49__22_;
      r_49__21_ <= r_n_49__21_;
      r_49__20_ <= r_n_49__20_;
      r_49__19_ <= r_n_49__19_;
      r_49__18_ <= r_n_49__18_;
      r_49__17_ <= r_n_49__17_;
      r_49__16_ <= r_n_49__16_;
      r_49__15_ <= r_n_49__15_;
      r_49__14_ <= r_n_49__14_;
      r_49__13_ <= r_n_49__13_;
      r_49__12_ <= r_n_49__12_;
      r_49__11_ <= r_n_49__11_;
      r_49__10_ <= r_n_49__10_;
      r_49__9_ <= r_n_49__9_;
      r_49__8_ <= r_n_49__8_;
      r_49__7_ <= r_n_49__7_;
      r_49__6_ <= r_n_49__6_;
      r_49__5_ <= r_n_49__5_;
      r_49__4_ <= r_n_49__4_;
      r_49__3_ <= r_n_49__3_;
      r_49__2_ <= r_n_49__2_;
      r_49__1_ <= r_n_49__1_;
      r_49__0_ <= r_n_49__0_;
    end 
    if(N3634) begin
      r_50__63_ <= r_n_50__63_;
      r_50__62_ <= r_n_50__62_;
      r_50__61_ <= r_n_50__61_;
      r_50__60_ <= r_n_50__60_;
      r_50__59_ <= r_n_50__59_;
      r_50__58_ <= r_n_50__58_;
      r_50__57_ <= r_n_50__57_;
      r_50__56_ <= r_n_50__56_;
      r_50__55_ <= r_n_50__55_;
      r_50__54_ <= r_n_50__54_;
      r_50__53_ <= r_n_50__53_;
      r_50__52_ <= r_n_50__52_;
      r_50__51_ <= r_n_50__51_;
      r_50__50_ <= r_n_50__50_;
      r_50__49_ <= r_n_50__49_;
      r_50__48_ <= r_n_50__48_;
      r_50__47_ <= r_n_50__47_;
      r_50__46_ <= r_n_50__46_;
      r_50__45_ <= r_n_50__45_;
      r_50__44_ <= r_n_50__44_;
      r_50__43_ <= r_n_50__43_;
      r_50__42_ <= r_n_50__42_;
      r_50__41_ <= r_n_50__41_;
      r_50__40_ <= r_n_50__40_;
      r_50__39_ <= r_n_50__39_;
      r_50__38_ <= r_n_50__38_;
      r_50__37_ <= r_n_50__37_;
      r_50__36_ <= r_n_50__36_;
      r_50__35_ <= r_n_50__35_;
      r_50__34_ <= r_n_50__34_;
      r_50__33_ <= r_n_50__33_;
      r_50__32_ <= r_n_50__32_;
      r_50__31_ <= r_n_50__31_;
      r_50__30_ <= r_n_50__30_;
      r_50__29_ <= r_n_50__29_;
      r_50__28_ <= r_n_50__28_;
      r_50__27_ <= r_n_50__27_;
      r_50__26_ <= r_n_50__26_;
      r_50__25_ <= r_n_50__25_;
      r_50__24_ <= r_n_50__24_;
      r_50__23_ <= r_n_50__23_;
      r_50__22_ <= r_n_50__22_;
      r_50__21_ <= r_n_50__21_;
      r_50__20_ <= r_n_50__20_;
      r_50__19_ <= r_n_50__19_;
      r_50__18_ <= r_n_50__18_;
      r_50__17_ <= r_n_50__17_;
      r_50__16_ <= r_n_50__16_;
      r_50__15_ <= r_n_50__15_;
      r_50__14_ <= r_n_50__14_;
      r_50__13_ <= r_n_50__13_;
      r_50__12_ <= r_n_50__12_;
      r_50__11_ <= r_n_50__11_;
      r_50__10_ <= r_n_50__10_;
      r_50__9_ <= r_n_50__9_;
      r_50__8_ <= r_n_50__8_;
      r_50__7_ <= r_n_50__7_;
      r_50__6_ <= r_n_50__6_;
      r_50__5_ <= r_n_50__5_;
      r_50__4_ <= r_n_50__4_;
      r_50__3_ <= r_n_50__3_;
      r_50__2_ <= r_n_50__2_;
      r_50__1_ <= r_n_50__1_;
      r_50__0_ <= r_n_50__0_;
    end 
    if(N3635) begin
      r_51__63_ <= r_n_51__63_;
      r_51__62_ <= r_n_51__62_;
      r_51__61_ <= r_n_51__61_;
      r_51__60_ <= r_n_51__60_;
      r_51__59_ <= r_n_51__59_;
      r_51__58_ <= r_n_51__58_;
      r_51__57_ <= r_n_51__57_;
      r_51__56_ <= r_n_51__56_;
      r_51__55_ <= r_n_51__55_;
      r_51__54_ <= r_n_51__54_;
      r_51__53_ <= r_n_51__53_;
      r_51__52_ <= r_n_51__52_;
      r_51__51_ <= r_n_51__51_;
      r_51__50_ <= r_n_51__50_;
      r_51__49_ <= r_n_51__49_;
      r_51__48_ <= r_n_51__48_;
      r_51__47_ <= r_n_51__47_;
      r_51__46_ <= r_n_51__46_;
      r_51__45_ <= r_n_51__45_;
      r_51__44_ <= r_n_51__44_;
      r_51__43_ <= r_n_51__43_;
      r_51__42_ <= r_n_51__42_;
      r_51__41_ <= r_n_51__41_;
      r_51__40_ <= r_n_51__40_;
      r_51__39_ <= r_n_51__39_;
      r_51__38_ <= r_n_51__38_;
      r_51__37_ <= r_n_51__37_;
      r_51__36_ <= r_n_51__36_;
      r_51__35_ <= r_n_51__35_;
      r_51__34_ <= r_n_51__34_;
      r_51__33_ <= r_n_51__33_;
      r_51__32_ <= r_n_51__32_;
      r_51__31_ <= r_n_51__31_;
      r_51__30_ <= r_n_51__30_;
      r_51__29_ <= r_n_51__29_;
      r_51__28_ <= r_n_51__28_;
      r_51__27_ <= r_n_51__27_;
      r_51__26_ <= r_n_51__26_;
      r_51__25_ <= r_n_51__25_;
      r_51__24_ <= r_n_51__24_;
      r_51__23_ <= r_n_51__23_;
      r_51__22_ <= r_n_51__22_;
      r_51__21_ <= r_n_51__21_;
      r_51__20_ <= r_n_51__20_;
      r_51__19_ <= r_n_51__19_;
      r_51__18_ <= r_n_51__18_;
      r_51__17_ <= r_n_51__17_;
      r_51__16_ <= r_n_51__16_;
      r_51__15_ <= r_n_51__15_;
      r_51__14_ <= r_n_51__14_;
      r_51__13_ <= r_n_51__13_;
      r_51__12_ <= r_n_51__12_;
      r_51__11_ <= r_n_51__11_;
      r_51__10_ <= r_n_51__10_;
      r_51__9_ <= r_n_51__9_;
      r_51__8_ <= r_n_51__8_;
      r_51__7_ <= r_n_51__7_;
      r_51__6_ <= r_n_51__6_;
      r_51__5_ <= r_n_51__5_;
      r_51__4_ <= r_n_51__4_;
      r_51__3_ <= r_n_51__3_;
      r_51__2_ <= r_n_51__2_;
      r_51__1_ <= r_n_51__1_;
      r_51__0_ <= r_n_51__0_;
    end 
    if(N3636) begin
      r_52__63_ <= r_n_52__63_;
      r_52__62_ <= r_n_52__62_;
      r_52__61_ <= r_n_52__61_;
      r_52__60_ <= r_n_52__60_;
      r_52__59_ <= r_n_52__59_;
      r_52__58_ <= r_n_52__58_;
      r_52__57_ <= r_n_52__57_;
      r_52__56_ <= r_n_52__56_;
      r_52__55_ <= r_n_52__55_;
      r_52__54_ <= r_n_52__54_;
      r_52__53_ <= r_n_52__53_;
      r_52__52_ <= r_n_52__52_;
      r_52__51_ <= r_n_52__51_;
      r_52__50_ <= r_n_52__50_;
      r_52__49_ <= r_n_52__49_;
      r_52__48_ <= r_n_52__48_;
      r_52__47_ <= r_n_52__47_;
      r_52__46_ <= r_n_52__46_;
      r_52__45_ <= r_n_52__45_;
      r_52__44_ <= r_n_52__44_;
      r_52__43_ <= r_n_52__43_;
      r_52__42_ <= r_n_52__42_;
      r_52__41_ <= r_n_52__41_;
      r_52__40_ <= r_n_52__40_;
      r_52__39_ <= r_n_52__39_;
      r_52__38_ <= r_n_52__38_;
      r_52__37_ <= r_n_52__37_;
      r_52__36_ <= r_n_52__36_;
      r_52__35_ <= r_n_52__35_;
      r_52__34_ <= r_n_52__34_;
      r_52__33_ <= r_n_52__33_;
      r_52__32_ <= r_n_52__32_;
      r_52__31_ <= r_n_52__31_;
      r_52__30_ <= r_n_52__30_;
      r_52__29_ <= r_n_52__29_;
      r_52__28_ <= r_n_52__28_;
      r_52__27_ <= r_n_52__27_;
      r_52__26_ <= r_n_52__26_;
      r_52__25_ <= r_n_52__25_;
      r_52__24_ <= r_n_52__24_;
      r_52__23_ <= r_n_52__23_;
      r_52__22_ <= r_n_52__22_;
      r_52__21_ <= r_n_52__21_;
      r_52__20_ <= r_n_52__20_;
      r_52__19_ <= r_n_52__19_;
      r_52__18_ <= r_n_52__18_;
      r_52__17_ <= r_n_52__17_;
      r_52__16_ <= r_n_52__16_;
      r_52__15_ <= r_n_52__15_;
      r_52__14_ <= r_n_52__14_;
      r_52__13_ <= r_n_52__13_;
      r_52__12_ <= r_n_52__12_;
      r_52__11_ <= r_n_52__11_;
      r_52__10_ <= r_n_52__10_;
      r_52__9_ <= r_n_52__9_;
      r_52__8_ <= r_n_52__8_;
      r_52__7_ <= r_n_52__7_;
      r_52__6_ <= r_n_52__6_;
      r_52__5_ <= r_n_52__5_;
      r_52__4_ <= r_n_52__4_;
      r_52__3_ <= r_n_52__3_;
      r_52__2_ <= r_n_52__2_;
      r_52__1_ <= r_n_52__1_;
      r_52__0_ <= r_n_52__0_;
    end 
    if(N3637) begin
      r_53__63_ <= r_n_53__63_;
      r_53__62_ <= r_n_53__62_;
      r_53__61_ <= r_n_53__61_;
      r_53__60_ <= r_n_53__60_;
      r_53__59_ <= r_n_53__59_;
      r_53__58_ <= r_n_53__58_;
      r_53__57_ <= r_n_53__57_;
      r_53__56_ <= r_n_53__56_;
      r_53__55_ <= r_n_53__55_;
      r_53__54_ <= r_n_53__54_;
      r_53__53_ <= r_n_53__53_;
      r_53__52_ <= r_n_53__52_;
      r_53__51_ <= r_n_53__51_;
      r_53__50_ <= r_n_53__50_;
      r_53__49_ <= r_n_53__49_;
      r_53__48_ <= r_n_53__48_;
      r_53__47_ <= r_n_53__47_;
      r_53__46_ <= r_n_53__46_;
      r_53__45_ <= r_n_53__45_;
      r_53__44_ <= r_n_53__44_;
      r_53__43_ <= r_n_53__43_;
      r_53__42_ <= r_n_53__42_;
      r_53__41_ <= r_n_53__41_;
      r_53__40_ <= r_n_53__40_;
      r_53__39_ <= r_n_53__39_;
      r_53__38_ <= r_n_53__38_;
      r_53__37_ <= r_n_53__37_;
      r_53__36_ <= r_n_53__36_;
      r_53__35_ <= r_n_53__35_;
      r_53__34_ <= r_n_53__34_;
      r_53__33_ <= r_n_53__33_;
      r_53__32_ <= r_n_53__32_;
      r_53__31_ <= r_n_53__31_;
      r_53__30_ <= r_n_53__30_;
      r_53__29_ <= r_n_53__29_;
      r_53__28_ <= r_n_53__28_;
      r_53__27_ <= r_n_53__27_;
      r_53__26_ <= r_n_53__26_;
      r_53__25_ <= r_n_53__25_;
      r_53__24_ <= r_n_53__24_;
      r_53__23_ <= r_n_53__23_;
      r_53__22_ <= r_n_53__22_;
      r_53__21_ <= r_n_53__21_;
      r_53__20_ <= r_n_53__20_;
      r_53__19_ <= r_n_53__19_;
      r_53__18_ <= r_n_53__18_;
      r_53__17_ <= r_n_53__17_;
      r_53__16_ <= r_n_53__16_;
      r_53__15_ <= r_n_53__15_;
      r_53__14_ <= r_n_53__14_;
      r_53__13_ <= r_n_53__13_;
      r_53__12_ <= r_n_53__12_;
      r_53__11_ <= r_n_53__11_;
      r_53__10_ <= r_n_53__10_;
      r_53__9_ <= r_n_53__9_;
      r_53__8_ <= r_n_53__8_;
      r_53__7_ <= r_n_53__7_;
      r_53__6_ <= r_n_53__6_;
      r_53__5_ <= r_n_53__5_;
      r_53__4_ <= r_n_53__4_;
      r_53__3_ <= r_n_53__3_;
      r_53__2_ <= r_n_53__2_;
      r_53__1_ <= r_n_53__1_;
      r_53__0_ <= r_n_53__0_;
    end 
    if(N3638) begin
      r_54__63_ <= r_n_54__63_;
      r_54__62_ <= r_n_54__62_;
      r_54__61_ <= r_n_54__61_;
      r_54__60_ <= r_n_54__60_;
      r_54__59_ <= r_n_54__59_;
      r_54__58_ <= r_n_54__58_;
      r_54__57_ <= r_n_54__57_;
      r_54__56_ <= r_n_54__56_;
      r_54__55_ <= r_n_54__55_;
      r_54__54_ <= r_n_54__54_;
      r_54__53_ <= r_n_54__53_;
      r_54__52_ <= r_n_54__52_;
      r_54__51_ <= r_n_54__51_;
      r_54__50_ <= r_n_54__50_;
      r_54__49_ <= r_n_54__49_;
      r_54__48_ <= r_n_54__48_;
      r_54__47_ <= r_n_54__47_;
      r_54__46_ <= r_n_54__46_;
      r_54__45_ <= r_n_54__45_;
      r_54__44_ <= r_n_54__44_;
      r_54__43_ <= r_n_54__43_;
      r_54__42_ <= r_n_54__42_;
      r_54__41_ <= r_n_54__41_;
      r_54__40_ <= r_n_54__40_;
      r_54__39_ <= r_n_54__39_;
      r_54__38_ <= r_n_54__38_;
      r_54__37_ <= r_n_54__37_;
      r_54__36_ <= r_n_54__36_;
      r_54__35_ <= r_n_54__35_;
      r_54__34_ <= r_n_54__34_;
      r_54__33_ <= r_n_54__33_;
      r_54__32_ <= r_n_54__32_;
      r_54__31_ <= r_n_54__31_;
      r_54__30_ <= r_n_54__30_;
      r_54__29_ <= r_n_54__29_;
      r_54__28_ <= r_n_54__28_;
      r_54__27_ <= r_n_54__27_;
      r_54__26_ <= r_n_54__26_;
      r_54__25_ <= r_n_54__25_;
      r_54__24_ <= r_n_54__24_;
      r_54__23_ <= r_n_54__23_;
      r_54__22_ <= r_n_54__22_;
      r_54__21_ <= r_n_54__21_;
      r_54__20_ <= r_n_54__20_;
      r_54__19_ <= r_n_54__19_;
      r_54__18_ <= r_n_54__18_;
      r_54__17_ <= r_n_54__17_;
      r_54__16_ <= r_n_54__16_;
      r_54__15_ <= r_n_54__15_;
      r_54__14_ <= r_n_54__14_;
      r_54__13_ <= r_n_54__13_;
      r_54__12_ <= r_n_54__12_;
      r_54__11_ <= r_n_54__11_;
      r_54__10_ <= r_n_54__10_;
      r_54__9_ <= r_n_54__9_;
      r_54__8_ <= r_n_54__8_;
      r_54__7_ <= r_n_54__7_;
      r_54__6_ <= r_n_54__6_;
      r_54__5_ <= r_n_54__5_;
      r_54__4_ <= r_n_54__4_;
      r_54__3_ <= r_n_54__3_;
      r_54__2_ <= r_n_54__2_;
      r_54__1_ <= r_n_54__1_;
      r_54__0_ <= r_n_54__0_;
    end 
    if(N3639) begin
      r_55__63_ <= r_n_55__63_;
      r_55__62_ <= r_n_55__62_;
      r_55__61_ <= r_n_55__61_;
      r_55__60_ <= r_n_55__60_;
      r_55__59_ <= r_n_55__59_;
      r_55__58_ <= r_n_55__58_;
      r_55__57_ <= r_n_55__57_;
      r_55__56_ <= r_n_55__56_;
      r_55__55_ <= r_n_55__55_;
      r_55__54_ <= r_n_55__54_;
      r_55__53_ <= r_n_55__53_;
      r_55__52_ <= r_n_55__52_;
      r_55__51_ <= r_n_55__51_;
      r_55__50_ <= r_n_55__50_;
      r_55__49_ <= r_n_55__49_;
      r_55__48_ <= r_n_55__48_;
      r_55__47_ <= r_n_55__47_;
      r_55__46_ <= r_n_55__46_;
      r_55__45_ <= r_n_55__45_;
      r_55__44_ <= r_n_55__44_;
      r_55__43_ <= r_n_55__43_;
      r_55__42_ <= r_n_55__42_;
      r_55__41_ <= r_n_55__41_;
      r_55__40_ <= r_n_55__40_;
      r_55__39_ <= r_n_55__39_;
      r_55__38_ <= r_n_55__38_;
      r_55__37_ <= r_n_55__37_;
      r_55__36_ <= r_n_55__36_;
      r_55__35_ <= r_n_55__35_;
      r_55__34_ <= r_n_55__34_;
      r_55__33_ <= r_n_55__33_;
      r_55__32_ <= r_n_55__32_;
      r_55__31_ <= r_n_55__31_;
      r_55__30_ <= r_n_55__30_;
      r_55__29_ <= r_n_55__29_;
      r_55__28_ <= r_n_55__28_;
      r_55__27_ <= r_n_55__27_;
      r_55__26_ <= r_n_55__26_;
      r_55__25_ <= r_n_55__25_;
      r_55__24_ <= r_n_55__24_;
      r_55__23_ <= r_n_55__23_;
      r_55__22_ <= r_n_55__22_;
      r_55__21_ <= r_n_55__21_;
      r_55__20_ <= r_n_55__20_;
      r_55__19_ <= r_n_55__19_;
      r_55__18_ <= r_n_55__18_;
      r_55__17_ <= r_n_55__17_;
      r_55__16_ <= r_n_55__16_;
      r_55__15_ <= r_n_55__15_;
      r_55__14_ <= r_n_55__14_;
      r_55__13_ <= r_n_55__13_;
      r_55__12_ <= r_n_55__12_;
      r_55__11_ <= r_n_55__11_;
      r_55__10_ <= r_n_55__10_;
      r_55__9_ <= r_n_55__9_;
      r_55__8_ <= r_n_55__8_;
      r_55__7_ <= r_n_55__7_;
      r_55__6_ <= r_n_55__6_;
      r_55__5_ <= r_n_55__5_;
      r_55__4_ <= r_n_55__4_;
      r_55__3_ <= r_n_55__3_;
      r_55__2_ <= r_n_55__2_;
      r_55__1_ <= r_n_55__1_;
      r_55__0_ <= r_n_55__0_;
    end 
    if(N3640) begin
      r_56__63_ <= r_n_56__63_;
      r_56__62_ <= r_n_56__62_;
      r_56__61_ <= r_n_56__61_;
      r_56__60_ <= r_n_56__60_;
      r_56__59_ <= r_n_56__59_;
      r_56__58_ <= r_n_56__58_;
      r_56__57_ <= r_n_56__57_;
      r_56__56_ <= r_n_56__56_;
      r_56__55_ <= r_n_56__55_;
      r_56__54_ <= r_n_56__54_;
      r_56__53_ <= r_n_56__53_;
      r_56__52_ <= r_n_56__52_;
      r_56__51_ <= r_n_56__51_;
      r_56__50_ <= r_n_56__50_;
      r_56__49_ <= r_n_56__49_;
      r_56__48_ <= r_n_56__48_;
      r_56__47_ <= r_n_56__47_;
      r_56__46_ <= r_n_56__46_;
      r_56__45_ <= r_n_56__45_;
      r_56__44_ <= r_n_56__44_;
      r_56__43_ <= r_n_56__43_;
      r_56__42_ <= r_n_56__42_;
      r_56__41_ <= r_n_56__41_;
      r_56__40_ <= r_n_56__40_;
      r_56__39_ <= r_n_56__39_;
      r_56__38_ <= r_n_56__38_;
      r_56__37_ <= r_n_56__37_;
      r_56__36_ <= r_n_56__36_;
      r_56__35_ <= r_n_56__35_;
      r_56__34_ <= r_n_56__34_;
      r_56__33_ <= r_n_56__33_;
      r_56__32_ <= r_n_56__32_;
      r_56__31_ <= r_n_56__31_;
      r_56__30_ <= r_n_56__30_;
      r_56__29_ <= r_n_56__29_;
      r_56__28_ <= r_n_56__28_;
      r_56__27_ <= r_n_56__27_;
      r_56__26_ <= r_n_56__26_;
      r_56__25_ <= r_n_56__25_;
      r_56__24_ <= r_n_56__24_;
      r_56__23_ <= r_n_56__23_;
      r_56__22_ <= r_n_56__22_;
      r_56__21_ <= r_n_56__21_;
      r_56__20_ <= r_n_56__20_;
      r_56__19_ <= r_n_56__19_;
      r_56__18_ <= r_n_56__18_;
      r_56__17_ <= r_n_56__17_;
      r_56__16_ <= r_n_56__16_;
      r_56__15_ <= r_n_56__15_;
      r_56__14_ <= r_n_56__14_;
      r_56__13_ <= r_n_56__13_;
      r_56__12_ <= r_n_56__12_;
      r_56__11_ <= r_n_56__11_;
      r_56__10_ <= r_n_56__10_;
      r_56__9_ <= r_n_56__9_;
      r_56__8_ <= r_n_56__8_;
      r_56__7_ <= r_n_56__7_;
      r_56__6_ <= r_n_56__6_;
      r_56__5_ <= r_n_56__5_;
      r_56__4_ <= r_n_56__4_;
      r_56__3_ <= r_n_56__3_;
      r_56__2_ <= r_n_56__2_;
      r_56__1_ <= r_n_56__1_;
      r_56__0_ <= r_n_56__0_;
    end 
    if(N3641) begin
      r_57__63_ <= r_n_57__63_;
      r_57__62_ <= r_n_57__62_;
      r_57__61_ <= r_n_57__61_;
      r_57__60_ <= r_n_57__60_;
      r_57__59_ <= r_n_57__59_;
      r_57__58_ <= r_n_57__58_;
      r_57__57_ <= r_n_57__57_;
      r_57__56_ <= r_n_57__56_;
      r_57__55_ <= r_n_57__55_;
      r_57__54_ <= r_n_57__54_;
      r_57__53_ <= r_n_57__53_;
      r_57__52_ <= r_n_57__52_;
      r_57__51_ <= r_n_57__51_;
      r_57__50_ <= r_n_57__50_;
      r_57__49_ <= r_n_57__49_;
      r_57__48_ <= r_n_57__48_;
      r_57__47_ <= r_n_57__47_;
      r_57__46_ <= r_n_57__46_;
      r_57__45_ <= r_n_57__45_;
      r_57__44_ <= r_n_57__44_;
      r_57__43_ <= r_n_57__43_;
      r_57__42_ <= r_n_57__42_;
      r_57__41_ <= r_n_57__41_;
      r_57__40_ <= r_n_57__40_;
      r_57__39_ <= r_n_57__39_;
      r_57__38_ <= r_n_57__38_;
      r_57__37_ <= r_n_57__37_;
      r_57__36_ <= r_n_57__36_;
      r_57__35_ <= r_n_57__35_;
      r_57__34_ <= r_n_57__34_;
      r_57__33_ <= r_n_57__33_;
      r_57__32_ <= r_n_57__32_;
      r_57__31_ <= r_n_57__31_;
      r_57__30_ <= r_n_57__30_;
      r_57__29_ <= r_n_57__29_;
      r_57__28_ <= r_n_57__28_;
      r_57__27_ <= r_n_57__27_;
      r_57__26_ <= r_n_57__26_;
      r_57__25_ <= r_n_57__25_;
      r_57__24_ <= r_n_57__24_;
      r_57__23_ <= r_n_57__23_;
      r_57__22_ <= r_n_57__22_;
      r_57__21_ <= r_n_57__21_;
      r_57__20_ <= r_n_57__20_;
      r_57__19_ <= r_n_57__19_;
      r_57__18_ <= r_n_57__18_;
      r_57__17_ <= r_n_57__17_;
      r_57__16_ <= r_n_57__16_;
      r_57__15_ <= r_n_57__15_;
      r_57__14_ <= r_n_57__14_;
      r_57__13_ <= r_n_57__13_;
      r_57__12_ <= r_n_57__12_;
      r_57__11_ <= r_n_57__11_;
      r_57__10_ <= r_n_57__10_;
      r_57__9_ <= r_n_57__9_;
      r_57__8_ <= r_n_57__8_;
      r_57__7_ <= r_n_57__7_;
      r_57__6_ <= r_n_57__6_;
      r_57__5_ <= r_n_57__5_;
      r_57__4_ <= r_n_57__4_;
      r_57__3_ <= r_n_57__3_;
      r_57__2_ <= r_n_57__2_;
      r_57__1_ <= r_n_57__1_;
      r_57__0_ <= r_n_57__0_;
    end 
    if(N3642) begin
      r_58__63_ <= r_n_58__63_;
      r_58__62_ <= r_n_58__62_;
      r_58__61_ <= r_n_58__61_;
      r_58__60_ <= r_n_58__60_;
      r_58__59_ <= r_n_58__59_;
      r_58__58_ <= r_n_58__58_;
      r_58__57_ <= r_n_58__57_;
      r_58__56_ <= r_n_58__56_;
      r_58__55_ <= r_n_58__55_;
      r_58__54_ <= r_n_58__54_;
      r_58__53_ <= r_n_58__53_;
      r_58__52_ <= r_n_58__52_;
      r_58__51_ <= r_n_58__51_;
      r_58__50_ <= r_n_58__50_;
      r_58__49_ <= r_n_58__49_;
      r_58__48_ <= r_n_58__48_;
      r_58__47_ <= r_n_58__47_;
      r_58__46_ <= r_n_58__46_;
      r_58__45_ <= r_n_58__45_;
      r_58__44_ <= r_n_58__44_;
      r_58__43_ <= r_n_58__43_;
      r_58__42_ <= r_n_58__42_;
      r_58__41_ <= r_n_58__41_;
      r_58__40_ <= r_n_58__40_;
      r_58__39_ <= r_n_58__39_;
      r_58__38_ <= r_n_58__38_;
      r_58__37_ <= r_n_58__37_;
      r_58__36_ <= r_n_58__36_;
      r_58__35_ <= r_n_58__35_;
      r_58__34_ <= r_n_58__34_;
      r_58__33_ <= r_n_58__33_;
      r_58__32_ <= r_n_58__32_;
      r_58__31_ <= r_n_58__31_;
      r_58__30_ <= r_n_58__30_;
      r_58__29_ <= r_n_58__29_;
      r_58__28_ <= r_n_58__28_;
      r_58__27_ <= r_n_58__27_;
      r_58__26_ <= r_n_58__26_;
      r_58__25_ <= r_n_58__25_;
      r_58__24_ <= r_n_58__24_;
      r_58__23_ <= r_n_58__23_;
      r_58__22_ <= r_n_58__22_;
      r_58__21_ <= r_n_58__21_;
      r_58__20_ <= r_n_58__20_;
      r_58__19_ <= r_n_58__19_;
      r_58__18_ <= r_n_58__18_;
      r_58__17_ <= r_n_58__17_;
      r_58__16_ <= r_n_58__16_;
      r_58__15_ <= r_n_58__15_;
      r_58__14_ <= r_n_58__14_;
      r_58__13_ <= r_n_58__13_;
      r_58__12_ <= r_n_58__12_;
      r_58__11_ <= r_n_58__11_;
      r_58__10_ <= r_n_58__10_;
      r_58__9_ <= r_n_58__9_;
      r_58__8_ <= r_n_58__8_;
      r_58__7_ <= r_n_58__7_;
      r_58__6_ <= r_n_58__6_;
      r_58__5_ <= r_n_58__5_;
      r_58__4_ <= r_n_58__4_;
      r_58__3_ <= r_n_58__3_;
      r_58__2_ <= r_n_58__2_;
      r_58__1_ <= r_n_58__1_;
      r_58__0_ <= r_n_58__0_;
    end 
    if(N3643) begin
      r_59__63_ <= r_n_59__63_;
      r_59__62_ <= r_n_59__62_;
      r_59__61_ <= r_n_59__61_;
      r_59__60_ <= r_n_59__60_;
      r_59__59_ <= r_n_59__59_;
      r_59__58_ <= r_n_59__58_;
      r_59__57_ <= r_n_59__57_;
      r_59__56_ <= r_n_59__56_;
      r_59__55_ <= r_n_59__55_;
      r_59__54_ <= r_n_59__54_;
      r_59__53_ <= r_n_59__53_;
      r_59__52_ <= r_n_59__52_;
      r_59__51_ <= r_n_59__51_;
      r_59__50_ <= r_n_59__50_;
      r_59__49_ <= r_n_59__49_;
      r_59__48_ <= r_n_59__48_;
      r_59__47_ <= r_n_59__47_;
      r_59__46_ <= r_n_59__46_;
      r_59__45_ <= r_n_59__45_;
      r_59__44_ <= r_n_59__44_;
      r_59__43_ <= r_n_59__43_;
      r_59__42_ <= r_n_59__42_;
      r_59__41_ <= r_n_59__41_;
      r_59__40_ <= r_n_59__40_;
      r_59__39_ <= r_n_59__39_;
      r_59__38_ <= r_n_59__38_;
      r_59__37_ <= r_n_59__37_;
      r_59__36_ <= r_n_59__36_;
      r_59__35_ <= r_n_59__35_;
      r_59__34_ <= r_n_59__34_;
      r_59__33_ <= r_n_59__33_;
      r_59__32_ <= r_n_59__32_;
      r_59__31_ <= r_n_59__31_;
      r_59__30_ <= r_n_59__30_;
      r_59__29_ <= r_n_59__29_;
      r_59__28_ <= r_n_59__28_;
      r_59__27_ <= r_n_59__27_;
      r_59__26_ <= r_n_59__26_;
      r_59__25_ <= r_n_59__25_;
      r_59__24_ <= r_n_59__24_;
      r_59__23_ <= r_n_59__23_;
      r_59__22_ <= r_n_59__22_;
      r_59__21_ <= r_n_59__21_;
      r_59__20_ <= r_n_59__20_;
      r_59__19_ <= r_n_59__19_;
      r_59__18_ <= r_n_59__18_;
      r_59__17_ <= r_n_59__17_;
      r_59__16_ <= r_n_59__16_;
      r_59__15_ <= r_n_59__15_;
      r_59__14_ <= r_n_59__14_;
      r_59__13_ <= r_n_59__13_;
      r_59__12_ <= r_n_59__12_;
      r_59__11_ <= r_n_59__11_;
      r_59__10_ <= r_n_59__10_;
      r_59__9_ <= r_n_59__9_;
      r_59__8_ <= r_n_59__8_;
      r_59__7_ <= r_n_59__7_;
      r_59__6_ <= r_n_59__6_;
      r_59__5_ <= r_n_59__5_;
      r_59__4_ <= r_n_59__4_;
      r_59__3_ <= r_n_59__3_;
      r_59__2_ <= r_n_59__2_;
      r_59__1_ <= r_n_59__1_;
      r_59__0_ <= r_n_59__0_;
    end 
    if(N3644) begin
      r_60__63_ <= r_n_60__63_;
      r_60__62_ <= r_n_60__62_;
      r_60__61_ <= r_n_60__61_;
      r_60__60_ <= r_n_60__60_;
      r_60__59_ <= r_n_60__59_;
      r_60__58_ <= r_n_60__58_;
      r_60__57_ <= r_n_60__57_;
      r_60__56_ <= r_n_60__56_;
      r_60__55_ <= r_n_60__55_;
      r_60__54_ <= r_n_60__54_;
      r_60__53_ <= r_n_60__53_;
      r_60__52_ <= r_n_60__52_;
      r_60__51_ <= r_n_60__51_;
      r_60__50_ <= r_n_60__50_;
      r_60__49_ <= r_n_60__49_;
      r_60__48_ <= r_n_60__48_;
      r_60__47_ <= r_n_60__47_;
      r_60__46_ <= r_n_60__46_;
      r_60__45_ <= r_n_60__45_;
      r_60__44_ <= r_n_60__44_;
      r_60__43_ <= r_n_60__43_;
      r_60__42_ <= r_n_60__42_;
      r_60__41_ <= r_n_60__41_;
      r_60__40_ <= r_n_60__40_;
      r_60__39_ <= r_n_60__39_;
      r_60__38_ <= r_n_60__38_;
      r_60__37_ <= r_n_60__37_;
      r_60__36_ <= r_n_60__36_;
      r_60__35_ <= r_n_60__35_;
      r_60__34_ <= r_n_60__34_;
      r_60__33_ <= r_n_60__33_;
      r_60__32_ <= r_n_60__32_;
      r_60__31_ <= r_n_60__31_;
      r_60__30_ <= r_n_60__30_;
      r_60__29_ <= r_n_60__29_;
      r_60__28_ <= r_n_60__28_;
      r_60__27_ <= r_n_60__27_;
      r_60__26_ <= r_n_60__26_;
      r_60__25_ <= r_n_60__25_;
      r_60__24_ <= r_n_60__24_;
      r_60__23_ <= r_n_60__23_;
      r_60__22_ <= r_n_60__22_;
      r_60__21_ <= r_n_60__21_;
      r_60__20_ <= r_n_60__20_;
      r_60__19_ <= r_n_60__19_;
      r_60__18_ <= r_n_60__18_;
      r_60__17_ <= r_n_60__17_;
      r_60__16_ <= r_n_60__16_;
      r_60__15_ <= r_n_60__15_;
      r_60__14_ <= r_n_60__14_;
      r_60__13_ <= r_n_60__13_;
      r_60__12_ <= r_n_60__12_;
      r_60__11_ <= r_n_60__11_;
      r_60__10_ <= r_n_60__10_;
      r_60__9_ <= r_n_60__9_;
      r_60__8_ <= r_n_60__8_;
      r_60__7_ <= r_n_60__7_;
      r_60__6_ <= r_n_60__6_;
      r_60__5_ <= r_n_60__5_;
      r_60__4_ <= r_n_60__4_;
      r_60__3_ <= r_n_60__3_;
      r_60__2_ <= r_n_60__2_;
      r_60__1_ <= r_n_60__1_;
      r_60__0_ <= r_n_60__0_;
    end 
    if(N3645) begin
      r_61__63_ <= r_n_61__63_;
      r_61__62_ <= r_n_61__62_;
      r_61__61_ <= r_n_61__61_;
      r_61__60_ <= r_n_61__60_;
      r_61__59_ <= r_n_61__59_;
      r_61__58_ <= r_n_61__58_;
      r_61__57_ <= r_n_61__57_;
      r_61__56_ <= r_n_61__56_;
      r_61__55_ <= r_n_61__55_;
      r_61__54_ <= r_n_61__54_;
      r_61__53_ <= r_n_61__53_;
      r_61__52_ <= r_n_61__52_;
      r_61__51_ <= r_n_61__51_;
      r_61__50_ <= r_n_61__50_;
      r_61__49_ <= r_n_61__49_;
      r_61__48_ <= r_n_61__48_;
      r_61__47_ <= r_n_61__47_;
      r_61__46_ <= r_n_61__46_;
      r_61__45_ <= r_n_61__45_;
      r_61__44_ <= r_n_61__44_;
      r_61__43_ <= r_n_61__43_;
      r_61__42_ <= r_n_61__42_;
      r_61__41_ <= r_n_61__41_;
      r_61__40_ <= r_n_61__40_;
      r_61__39_ <= r_n_61__39_;
      r_61__38_ <= r_n_61__38_;
      r_61__37_ <= r_n_61__37_;
      r_61__36_ <= r_n_61__36_;
      r_61__35_ <= r_n_61__35_;
      r_61__34_ <= r_n_61__34_;
      r_61__33_ <= r_n_61__33_;
      r_61__32_ <= r_n_61__32_;
      r_61__31_ <= r_n_61__31_;
      r_61__30_ <= r_n_61__30_;
      r_61__29_ <= r_n_61__29_;
      r_61__28_ <= r_n_61__28_;
      r_61__27_ <= r_n_61__27_;
      r_61__26_ <= r_n_61__26_;
      r_61__25_ <= r_n_61__25_;
      r_61__24_ <= r_n_61__24_;
      r_61__23_ <= r_n_61__23_;
      r_61__22_ <= r_n_61__22_;
      r_61__21_ <= r_n_61__21_;
      r_61__20_ <= r_n_61__20_;
      r_61__19_ <= r_n_61__19_;
      r_61__18_ <= r_n_61__18_;
      r_61__17_ <= r_n_61__17_;
      r_61__16_ <= r_n_61__16_;
      r_61__15_ <= r_n_61__15_;
      r_61__14_ <= r_n_61__14_;
      r_61__13_ <= r_n_61__13_;
      r_61__12_ <= r_n_61__12_;
      r_61__11_ <= r_n_61__11_;
      r_61__10_ <= r_n_61__10_;
      r_61__9_ <= r_n_61__9_;
      r_61__8_ <= r_n_61__8_;
      r_61__7_ <= r_n_61__7_;
      r_61__6_ <= r_n_61__6_;
      r_61__5_ <= r_n_61__5_;
      r_61__4_ <= r_n_61__4_;
      r_61__3_ <= r_n_61__3_;
      r_61__2_ <= r_n_61__2_;
      r_61__1_ <= r_n_61__1_;
      r_61__0_ <= r_n_61__0_;
    end 
    if(N3646) begin
      r_62__63_ <= r_n_62__63_;
      r_62__62_ <= r_n_62__62_;
      r_62__61_ <= r_n_62__61_;
      r_62__60_ <= r_n_62__60_;
      r_62__59_ <= r_n_62__59_;
      r_62__58_ <= r_n_62__58_;
      r_62__57_ <= r_n_62__57_;
      r_62__56_ <= r_n_62__56_;
      r_62__55_ <= r_n_62__55_;
      r_62__54_ <= r_n_62__54_;
      r_62__53_ <= r_n_62__53_;
      r_62__52_ <= r_n_62__52_;
      r_62__51_ <= r_n_62__51_;
      r_62__50_ <= r_n_62__50_;
      r_62__49_ <= r_n_62__49_;
      r_62__48_ <= r_n_62__48_;
      r_62__47_ <= r_n_62__47_;
      r_62__46_ <= r_n_62__46_;
      r_62__45_ <= r_n_62__45_;
      r_62__44_ <= r_n_62__44_;
      r_62__43_ <= r_n_62__43_;
      r_62__42_ <= r_n_62__42_;
      r_62__41_ <= r_n_62__41_;
      r_62__40_ <= r_n_62__40_;
      r_62__39_ <= r_n_62__39_;
      r_62__38_ <= r_n_62__38_;
      r_62__37_ <= r_n_62__37_;
      r_62__36_ <= r_n_62__36_;
      r_62__35_ <= r_n_62__35_;
      r_62__34_ <= r_n_62__34_;
      r_62__33_ <= r_n_62__33_;
      r_62__32_ <= r_n_62__32_;
      r_62__31_ <= r_n_62__31_;
      r_62__30_ <= r_n_62__30_;
      r_62__29_ <= r_n_62__29_;
      r_62__28_ <= r_n_62__28_;
      r_62__27_ <= r_n_62__27_;
      r_62__26_ <= r_n_62__26_;
      r_62__25_ <= r_n_62__25_;
      r_62__24_ <= r_n_62__24_;
      r_62__23_ <= r_n_62__23_;
      r_62__22_ <= r_n_62__22_;
      r_62__21_ <= r_n_62__21_;
      r_62__20_ <= r_n_62__20_;
      r_62__19_ <= r_n_62__19_;
      r_62__18_ <= r_n_62__18_;
      r_62__17_ <= r_n_62__17_;
      r_62__16_ <= r_n_62__16_;
      r_62__15_ <= r_n_62__15_;
      r_62__14_ <= r_n_62__14_;
      r_62__13_ <= r_n_62__13_;
      r_62__12_ <= r_n_62__12_;
      r_62__11_ <= r_n_62__11_;
      r_62__10_ <= r_n_62__10_;
      r_62__9_ <= r_n_62__9_;
      r_62__8_ <= r_n_62__8_;
      r_62__7_ <= r_n_62__7_;
      r_62__6_ <= r_n_62__6_;
      r_62__5_ <= r_n_62__5_;
      r_62__4_ <= r_n_62__4_;
      r_62__3_ <= r_n_62__3_;
      r_62__2_ <= r_n_62__2_;
      r_62__1_ <= r_n_62__1_;
      r_62__0_ <= r_n_62__0_;
    end 
    if(N3647) begin
      r_63__63_ <= r_n_63__63_;
      r_63__62_ <= r_n_63__62_;
      r_63__61_ <= r_n_63__61_;
      r_63__60_ <= r_n_63__60_;
      r_63__59_ <= r_n_63__59_;
      r_63__58_ <= r_n_63__58_;
      r_63__57_ <= r_n_63__57_;
      r_63__56_ <= r_n_63__56_;
      r_63__55_ <= r_n_63__55_;
      r_63__54_ <= r_n_63__54_;
      r_63__53_ <= r_n_63__53_;
      r_63__52_ <= r_n_63__52_;
      r_63__51_ <= r_n_63__51_;
      r_63__50_ <= r_n_63__50_;
      r_63__49_ <= r_n_63__49_;
      r_63__48_ <= r_n_63__48_;
      r_63__47_ <= r_n_63__47_;
      r_63__46_ <= r_n_63__46_;
      r_63__45_ <= r_n_63__45_;
      r_63__44_ <= r_n_63__44_;
      r_63__43_ <= r_n_63__43_;
      r_63__42_ <= r_n_63__42_;
      r_63__41_ <= r_n_63__41_;
      r_63__40_ <= r_n_63__40_;
      r_63__39_ <= r_n_63__39_;
      r_63__38_ <= r_n_63__38_;
      r_63__37_ <= r_n_63__37_;
      r_63__36_ <= r_n_63__36_;
      r_63__35_ <= r_n_63__35_;
      r_63__34_ <= r_n_63__34_;
      r_63__33_ <= r_n_63__33_;
      r_63__32_ <= r_n_63__32_;
      r_63__31_ <= r_n_63__31_;
      r_63__30_ <= r_n_63__30_;
      r_63__29_ <= r_n_63__29_;
      r_63__28_ <= r_n_63__28_;
      r_63__27_ <= r_n_63__27_;
      r_63__26_ <= r_n_63__26_;
      r_63__25_ <= r_n_63__25_;
      r_63__24_ <= r_n_63__24_;
      r_63__23_ <= r_n_63__23_;
      r_63__22_ <= r_n_63__22_;
      r_63__21_ <= r_n_63__21_;
      r_63__20_ <= r_n_63__20_;
      r_63__19_ <= r_n_63__19_;
      r_63__18_ <= r_n_63__18_;
      r_63__17_ <= r_n_63__17_;
      r_63__16_ <= r_n_63__16_;
      r_63__15_ <= r_n_63__15_;
      r_63__14_ <= r_n_63__14_;
      r_63__13_ <= r_n_63__13_;
      r_63__12_ <= r_n_63__12_;
      r_63__11_ <= r_n_63__11_;
      r_63__10_ <= r_n_63__10_;
      r_63__9_ <= r_n_63__9_;
      r_63__8_ <= r_n_63__8_;
      r_63__7_ <= r_n_63__7_;
      r_63__6_ <= r_n_63__6_;
      r_63__5_ <= r_n_63__5_;
      r_63__4_ <= r_n_63__4_;
      r_63__3_ <= r_n_63__3_;
      r_63__2_ <= r_n_63__2_;
      r_63__1_ <= r_n_63__1_;
      r_63__0_ <= r_n_63__0_;
    end 
    if(N3648) begin
      r_64__63_ <= r_n_64__63_;
      r_64__62_ <= r_n_64__62_;
      r_64__61_ <= r_n_64__61_;
      r_64__60_ <= r_n_64__60_;
      r_64__59_ <= r_n_64__59_;
      r_64__58_ <= r_n_64__58_;
      r_64__57_ <= r_n_64__57_;
      r_64__56_ <= r_n_64__56_;
      r_64__55_ <= r_n_64__55_;
      r_64__54_ <= r_n_64__54_;
      r_64__53_ <= r_n_64__53_;
      r_64__52_ <= r_n_64__52_;
      r_64__51_ <= r_n_64__51_;
      r_64__50_ <= r_n_64__50_;
      r_64__49_ <= r_n_64__49_;
      r_64__48_ <= r_n_64__48_;
      r_64__47_ <= r_n_64__47_;
      r_64__46_ <= r_n_64__46_;
      r_64__45_ <= r_n_64__45_;
      r_64__44_ <= r_n_64__44_;
      r_64__43_ <= r_n_64__43_;
      r_64__42_ <= r_n_64__42_;
      r_64__41_ <= r_n_64__41_;
      r_64__40_ <= r_n_64__40_;
      r_64__39_ <= r_n_64__39_;
      r_64__38_ <= r_n_64__38_;
      r_64__37_ <= r_n_64__37_;
      r_64__36_ <= r_n_64__36_;
      r_64__35_ <= r_n_64__35_;
      r_64__34_ <= r_n_64__34_;
      r_64__33_ <= r_n_64__33_;
      r_64__32_ <= r_n_64__32_;
      r_64__31_ <= r_n_64__31_;
      r_64__30_ <= r_n_64__30_;
      r_64__29_ <= r_n_64__29_;
      r_64__28_ <= r_n_64__28_;
      r_64__27_ <= r_n_64__27_;
      r_64__26_ <= r_n_64__26_;
      r_64__25_ <= r_n_64__25_;
      r_64__24_ <= r_n_64__24_;
      r_64__23_ <= r_n_64__23_;
      r_64__22_ <= r_n_64__22_;
      r_64__21_ <= r_n_64__21_;
      r_64__20_ <= r_n_64__20_;
      r_64__19_ <= r_n_64__19_;
      r_64__18_ <= r_n_64__18_;
      r_64__17_ <= r_n_64__17_;
      r_64__16_ <= r_n_64__16_;
      r_64__15_ <= r_n_64__15_;
      r_64__14_ <= r_n_64__14_;
      r_64__13_ <= r_n_64__13_;
      r_64__12_ <= r_n_64__12_;
      r_64__11_ <= r_n_64__11_;
      r_64__10_ <= r_n_64__10_;
      r_64__9_ <= r_n_64__9_;
      r_64__8_ <= r_n_64__8_;
      r_64__7_ <= r_n_64__7_;
      r_64__6_ <= r_n_64__6_;
      r_64__5_ <= r_n_64__5_;
      r_64__4_ <= r_n_64__4_;
      r_64__3_ <= r_n_64__3_;
      r_64__2_ <= r_n_64__2_;
      r_64__1_ <= r_n_64__1_;
      r_64__0_ <= r_n_64__0_;
    end 
    if(N3649) begin
      r_65__63_ <= r_n_65__63_;
      r_65__62_ <= r_n_65__62_;
      r_65__61_ <= r_n_65__61_;
      r_65__60_ <= r_n_65__60_;
      r_65__59_ <= r_n_65__59_;
      r_65__58_ <= r_n_65__58_;
      r_65__57_ <= r_n_65__57_;
      r_65__56_ <= r_n_65__56_;
      r_65__55_ <= r_n_65__55_;
      r_65__54_ <= r_n_65__54_;
      r_65__53_ <= r_n_65__53_;
      r_65__52_ <= r_n_65__52_;
      r_65__51_ <= r_n_65__51_;
      r_65__50_ <= r_n_65__50_;
      r_65__49_ <= r_n_65__49_;
      r_65__48_ <= r_n_65__48_;
      r_65__47_ <= r_n_65__47_;
      r_65__46_ <= r_n_65__46_;
      r_65__45_ <= r_n_65__45_;
      r_65__44_ <= r_n_65__44_;
      r_65__43_ <= r_n_65__43_;
      r_65__42_ <= r_n_65__42_;
      r_65__41_ <= r_n_65__41_;
      r_65__40_ <= r_n_65__40_;
      r_65__39_ <= r_n_65__39_;
      r_65__38_ <= r_n_65__38_;
      r_65__37_ <= r_n_65__37_;
      r_65__36_ <= r_n_65__36_;
      r_65__35_ <= r_n_65__35_;
      r_65__34_ <= r_n_65__34_;
      r_65__33_ <= r_n_65__33_;
      r_65__32_ <= r_n_65__32_;
      r_65__31_ <= r_n_65__31_;
      r_65__30_ <= r_n_65__30_;
      r_65__29_ <= r_n_65__29_;
      r_65__28_ <= r_n_65__28_;
      r_65__27_ <= r_n_65__27_;
      r_65__26_ <= r_n_65__26_;
      r_65__25_ <= r_n_65__25_;
      r_65__24_ <= r_n_65__24_;
      r_65__23_ <= r_n_65__23_;
      r_65__22_ <= r_n_65__22_;
      r_65__21_ <= r_n_65__21_;
      r_65__20_ <= r_n_65__20_;
      r_65__19_ <= r_n_65__19_;
      r_65__18_ <= r_n_65__18_;
      r_65__17_ <= r_n_65__17_;
      r_65__16_ <= r_n_65__16_;
      r_65__15_ <= r_n_65__15_;
      r_65__14_ <= r_n_65__14_;
      r_65__13_ <= r_n_65__13_;
      r_65__12_ <= r_n_65__12_;
      r_65__11_ <= r_n_65__11_;
      r_65__10_ <= r_n_65__10_;
      r_65__9_ <= r_n_65__9_;
      r_65__8_ <= r_n_65__8_;
      r_65__7_ <= r_n_65__7_;
      r_65__6_ <= r_n_65__6_;
      r_65__5_ <= r_n_65__5_;
      r_65__4_ <= r_n_65__4_;
      r_65__3_ <= r_n_65__3_;
      r_65__2_ <= r_n_65__2_;
      r_65__1_ <= r_n_65__1_;
      r_65__0_ <= r_n_65__0_;
    end 
    if(N3650) begin
      r_66__63_ <= r_n_66__63_;
      r_66__62_ <= r_n_66__62_;
      r_66__61_ <= r_n_66__61_;
      r_66__60_ <= r_n_66__60_;
      r_66__59_ <= r_n_66__59_;
      r_66__58_ <= r_n_66__58_;
      r_66__57_ <= r_n_66__57_;
      r_66__56_ <= r_n_66__56_;
      r_66__55_ <= r_n_66__55_;
      r_66__54_ <= r_n_66__54_;
      r_66__53_ <= r_n_66__53_;
      r_66__52_ <= r_n_66__52_;
      r_66__51_ <= r_n_66__51_;
      r_66__50_ <= r_n_66__50_;
      r_66__49_ <= r_n_66__49_;
      r_66__48_ <= r_n_66__48_;
      r_66__47_ <= r_n_66__47_;
      r_66__46_ <= r_n_66__46_;
      r_66__45_ <= r_n_66__45_;
      r_66__44_ <= r_n_66__44_;
      r_66__43_ <= r_n_66__43_;
      r_66__42_ <= r_n_66__42_;
      r_66__41_ <= r_n_66__41_;
      r_66__40_ <= r_n_66__40_;
      r_66__39_ <= r_n_66__39_;
      r_66__38_ <= r_n_66__38_;
      r_66__37_ <= r_n_66__37_;
      r_66__36_ <= r_n_66__36_;
      r_66__35_ <= r_n_66__35_;
      r_66__34_ <= r_n_66__34_;
      r_66__33_ <= r_n_66__33_;
      r_66__32_ <= r_n_66__32_;
      r_66__31_ <= r_n_66__31_;
      r_66__30_ <= r_n_66__30_;
      r_66__29_ <= r_n_66__29_;
      r_66__28_ <= r_n_66__28_;
      r_66__27_ <= r_n_66__27_;
      r_66__26_ <= r_n_66__26_;
      r_66__25_ <= r_n_66__25_;
      r_66__24_ <= r_n_66__24_;
      r_66__23_ <= r_n_66__23_;
      r_66__22_ <= r_n_66__22_;
      r_66__21_ <= r_n_66__21_;
      r_66__20_ <= r_n_66__20_;
      r_66__19_ <= r_n_66__19_;
      r_66__18_ <= r_n_66__18_;
      r_66__17_ <= r_n_66__17_;
      r_66__16_ <= r_n_66__16_;
      r_66__15_ <= r_n_66__15_;
      r_66__14_ <= r_n_66__14_;
      r_66__13_ <= r_n_66__13_;
      r_66__12_ <= r_n_66__12_;
      r_66__11_ <= r_n_66__11_;
      r_66__10_ <= r_n_66__10_;
      r_66__9_ <= r_n_66__9_;
      r_66__8_ <= r_n_66__8_;
      r_66__7_ <= r_n_66__7_;
      r_66__6_ <= r_n_66__6_;
      r_66__5_ <= r_n_66__5_;
      r_66__4_ <= r_n_66__4_;
      r_66__3_ <= r_n_66__3_;
      r_66__2_ <= r_n_66__2_;
      r_66__1_ <= r_n_66__1_;
      r_66__0_ <= r_n_66__0_;
    end 
    if(N3651) begin
      r_67__63_ <= r_n_67__63_;
      r_67__62_ <= r_n_67__62_;
      r_67__61_ <= r_n_67__61_;
      r_67__60_ <= r_n_67__60_;
      r_67__59_ <= r_n_67__59_;
      r_67__58_ <= r_n_67__58_;
      r_67__57_ <= r_n_67__57_;
      r_67__56_ <= r_n_67__56_;
      r_67__55_ <= r_n_67__55_;
      r_67__54_ <= r_n_67__54_;
      r_67__53_ <= r_n_67__53_;
      r_67__52_ <= r_n_67__52_;
      r_67__51_ <= r_n_67__51_;
      r_67__50_ <= r_n_67__50_;
      r_67__49_ <= r_n_67__49_;
      r_67__48_ <= r_n_67__48_;
      r_67__47_ <= r_n_67__47_;
      r_67__46_ <= r_n_67__46_;
      r_67__45_ <= r_n_67__45_;
      r_67__44_ <= r_n_67__44_;
      r_67__43_ <= r_n_67__43_;
      r_67__42_ <= r_n_67__42_;
      r_67__41_ <= r_n_67__41_;
      r_67__40_ <= r_n_67__40_;
      r_67__39_ <= r_n_67__39_;
      r_67__38_ <= r_n_67__38_;
      r_67__37_ <= r_n_67__37_;
      r_67__36_ <= r_n_67__36_;
      r_67__35_ <= r_n_67__35_;
      r_67__34_ <= r_n_67__34_;
      r_67__33_ <= r_n_67__33_;
      r_67__32_ <= r_n_67__32_;
      r_67__31_ <= r_n_67__31_;
      r_67__30_ <= r_n_67__30_;
      r_67__29_ <= r_n_67__29_;
      r_67__28_ <= r_n_67__28_;
      r_67__27_ <= r_n_67__27_;
      r_67__26_ <= r_n_67__26_;
      r_67__25_ <= r_n_67__25_;
      r_67__24_ <= r_n_67__24_;
      r_67__23_ <= r_n_67__23_;
      r_67__22_ <= r_n_67__22_;
      r_67__21_ <= r_n_67__21_;
      r_67__20_ <= r_n_67__20_;
      r_67__19_ <= r_n_67__19_;
      r_67__18_ <= r_n_67__18_;
      r_67__17_ <= r_n_67__17_;
      r_67__16_ <= r_n_67__16_;
      r_67__15_ <= r_n_67__15_;
      r_67__14_ <= r_n_67__14_;
      r_67__13_ <= r_n_67__13_;
      r_67__12_ <= r_n_67__12_;
      r_67__11_ <= r_n_67__11_;
      r_67__10_ <= r_n_67__10_;
      r_67__9_ <= r_n_67__9_;
      r_67__8_ <= r_n_67__8_;
      r_67__7_ <= r_n_67__7_;
      r_67__6_ <= r_n_67__6_;
      r_67__5_ <= r_n_67__5_;
      r_67__4_ <= r_n_67__4_;
      r_67__3_ <= r_n_67__3_;
      r_67__2_ <= r_n_67__2_;
      r_67__1_ <= r_n_67__1_;
      r_67__0_ <= r_n_67__0_;
    end 
    if(N3652) begin
      r_68__63_ <= r_n_68__63_;
      r_68__62_ <= r_n_68__62_;
      r_68__61_ <= r_n_68__61_;
      r_68__60_ <= r_n_68__60_;
      r_68__59_ <= r_n_68__59_;
      r_68__58_ <= r_n_68__58_;
      r_68__57_ <= r_n_68__57_;
      r_68__56_ <= r_n_68__56_;
      r_68__55_ <= r_n_68__55_;
      r_68__54_ <= r_n_68__54_;
      r_68__53_ <= r_n_68__53_;
      r_68__52_ <= r_n_68__52_;
      r_68__51_ <= r_n_68__51_;
      r_68__50_ <= r_n_68__50_;
      r_68__49_ <= r_n_68__49_;
      r_68__48_ <= r_n_68__48_;
      r_68__47_ <= r_n_68__47_;
      r_68__46_ <= r_n_68__46_;
      r_68__45_ <= r_n_68__45_;
      r_68__44_ <= r_n_68__44_;
      r_68__43_ <= r_n_68__43_;
      r_68__42_ <= r_n_68__42_;
      r_68__41_ <= r_n_68__41_;
      r_68__40_ <= r_n_68__40_;
      r_68__39_ <= r_n_68__39_;
      r_68__38_ <= r_n_68__38_;
      r_68__37_ <= r_n_68__37_;
      r_68__36_ <= r_n_68__36_;
      r_68__35_ <= r_n_68__35_;
      r_68__34_ <= r_n_68__34_;
      r_68__33_ <= r_n_68__33_;
      r_68__32_ <= r_n_68__32_;
      r_68__31_ <= r_n_68__31_;
      r_68__30_ <= r_n_68__30_;
      r_68__29_ <= r_n_68__29_;
      r_68__28_ <= r_n_68__28_;
      r_68__27_ <= r_n_68__27_;
      r_68__26_ <= r_n_68__26_;
      r_68__25_ <= r_n_68__25_;
      r_68__24_ <= r_n_68__24_;
      r_68__23_ <= r_n_68__23_;
      r_68__22_ <= r_n_68__22_;
      r_68__21_ <= r_n_68__21_;
      r_68__20_ <= r_n_68__20_;
      r_68__19_ <= r_n_68__19_;
      r_68__18_ <= r_n_68__18_;
      r_68__17_ <= r_n_68__17_;
      r_68__16_ <= r_n_68__16_;
      r_68__15_ <= r_n_68__15_;
      r_68__14_ <= r_n_68__14_;
      r_68__13_ <= r_n_68__13_;
      r_68__12_ <= r_n_68__12_;
      r_68__11_ <= r_n_68__11_;
      r_68__10_ <= r_n_68__10_;
      r_68__9_ <= r_n_68__9_;
      r_68__8_ <= r_n_68__8_;
      r_68__7_ <= r_n_68__7_;
      r_68__6_ <= r_n_68__6_;
      r_68__5_ <= r_n_68__5_;
      r_68__4_ <= r_n_68__4_;
      r_68__3_ <= r_n_68__3_;
      r_68__2_ <= r_n_68__2_;
      r_68__1_ <= r_n_68__1_;
      r_68__0_ <= r_n_68__0_;
    end 
    if(N3653) begin
      r_69__63_ <= r_n_69__63_;
      r_69__62_ <= r_n_69__62_;
      r_69__61_ <= r_n_69__61_;
      r_69__60_ <= r_n_69__60_;
      r_69__59_ <= r_n_69__59_;
      r_69__58_ <= r_n_69__58_;
      r_69__57_ <= r_n_69__57_;
      r_69__56_ <= r_n_69__56_;
      r_69__55_ <= r_n_69__55_;
      r_69__54_ <= r_n_69__54_;
      r_69__53_ <= r_n_69__53_;
      r_69__52_ <= r_n_69__52_;
      r_69__51_ <= r_n_69__51_;
      r_69__50_ <= r_n_69__50_;
      r_69__49_ <= r_n_69__49_;
      r_69__48_ <= r_n_69__48_;
      r_69__47_ <= r_n_69__47_;
      r_69__46_ <= r_n_69__46_;
      r_69__45_ <= r_n_69__45_;
      r_69__44_ <= r_n_69__44_;
      r_69__43_ <= r_n_69__43_;
      r_69__42_ <= r_n_69__42_;
      r_69__41_ <= r_n_69__41_;
      r_69__40_ <= r_n_69__40_;
      r_69__39_ <= r_n_69__39_;
      r_69__38_ <= r_n_69__38_;
      r_69__37_ <= r_n_69__37_;
      r_69__36_ <= r_n_69__36_;
      r_69__35_ <= r_n_69__35_;
      r_69__34_ <= r_n_69__34_;
      r_69__33_ <= r_n_69__33_;
      r_69__32_ <= r_n_69__32_;
      r_69__31_ <= r_n_69__31_;
      r_69__30_ <= r_n_69__30_;
      r_69__29_ <= r_n_69__29_;
      r_69__28_ <= r_n_69__28_;
      r_69__27_ <= r_n_69__27_;
      r_69__26_ <= r_n_69__26_;
      r_69__25_ <= r_n_69__25_;
      r_69__24_ <= r_n_69__24_;
      r_69__23_ <= r_n_69__23_;
      r_69__22_ <= r_n_69__22_;
      r_69__21_ <= r_n_69__21_;
      r_69__20_ <= r_n_69__20_;
      r_69__19_ <= r_n_69__19_;
      r_69__18_ <= r_n_69__18_;
      r_69__17_ <= r_n_69__17_;
      r_69__16_ <= r_n_69__16_;
      r_69__15_ <= r_n_69__15_;
      r_69__14_ <= r_n_69__14_;
      r_69__13_ <= r_n_69__13_;
      r_69__12_ <= r_n_69__12_;
      r_69__11_ <= r_n_69__11_;
      r_69__10_ <= r_n_69__10_;
      r_69__9_ <= r_n_69__9_;
      r_69__8_ <= r_n_69__8_;
      r_69__7_ <= r_n_69__7_;
      r_69__6_ <= r_n_69__6_;
      r_69__5_ <= r_n_69__5_;
      r_69__4_ <= r_n_69__4_;
      r_69__3_ <= r_n_69__3_;
      r_69__2_ <= r_n_69__2_;
      r_69__1_ <= r_n_69__1_;
      r_69__0_ <= r_n_69__0_;
    end 
    if(N3654) begin
      r_70__63_ <= r_n_70__63_;
      r_70__62_ <= r_n_70__62_;
      r_70__61_ <= r_n_70__61_;
      r_70__60_ <= r_n_70__60_;
      r_70__59_ <= r_n_70__59_;
      r_70__58_ <= r_n_70__58_;
      r_70__57_ <= r_n_70__57_;
      r_70__56_ <= r_n_70__56_;
      r_70__55_ <= r_n_70__55_;
      r_70__54_ <= r_n_70__54_;
      r_70__53_ <= r_n_70__53_;
      r_70__52_ <= r_n_70__52_;
      r_70__51_ <= r_n_70__51_;
      r_70__50_ <= r_n_70__50_;
      r_70__49_ <= r_n_70__49_;
      r_70__48_ <= r_n_70__48_;
      r_70__47_ <= r_n_70__47_;
      r_70__46_ <= r_n_70__46_;
      r_70__45_ <= r_n_70__45_;
      r_70__44_ <= r_n_70__44_;
      r_70__43_ <= r_n_70__43_;
      r_70__42_ <= r_n_70__42_;
      r_70__41_ <= r_n_70__41_;
      r_70__40_ <= r_n_70__40_;
      r_70__39_ <= r_n_70__39_;
      r_70__38_ <= r_n_70__38_;
      r_70__37_ <= r_n_70__37_;
      r_70__36_ <= r_n_70__36_;
      r_70__35_ <= r_n_70__35_;
      r_70__34_ <= r_n_70__34_;
      r_70__33_ <= r_n_70__33_;
      r_70__32_ <= r_n_70__32_;
      r_70__31_ <= r_n_70__31_;
      r_70__30_ <= r_n_70__30_;
      r_70__29_ <= r_n_70__29_;
      r_70__28_ <= r_n_70__28_;
      r_70__27_ <= r_n_70__27_;
      r_70__26_ <= r_n_70__26_;
      r_70__25_ <= r_n_70__25_;
      r_70__24_ <= r_n_70__24_;
      r_70__23_ <= r_n_70__23_;
      r_70__22_ <= r_n_70__22_;
      r_70__21_ <= r_n_70__21_;
      r_70__20_ <= r_n_70__20_;
      r_70__19_ <= r_n_70__19_;
      r_70__18_ <= r_n_70__18_;
      r_70__17_ <= r_n_70__17_;
      r_70__16_ <= r_n_70__16_;
      r_70__15_ <= r_n_70__15_;
      r_70__14_ <= r_n_70__14_;
      r_70__13_ <= r_n_70__13_;
      r_70__12_ <= r_n_70__12_;
      r_70__11_ <= r_n_70__11_;
      r_70__10_ <= r_n_70__10_;
      r_70__9_ <= r_n_70__9_;
      r_70__8_ <= r_n_70__8_;
      r_70__7_ <= r_n_70__7_;
      r_70__6_ <= r_n_70__6_;
      r_70__5_ <= r_n_70__5_;
      r_70__4_ <= r_n_70__4_;
      r_70__3_ <= r_n_70__3_;
      r_70__2_ <= r_n_70__2_;
      r_70__1_ <= r_n_70__1_;
      r_70__0_ <= r_n_70__0_;
    end 
    if(N3655) begin
      r_71__63_ <= r_n_71__63_;
      r_71__62_ <= r_n_71__62_;
      r_71__61_ <= r_n_71__61_;
      r_71__60_ <= r_n_71__60_;
      r_71__59_ <= r_n_71__59_;
      r_71__58_ <= r_n_71__58_;
      r_71__57_ <= r_n_71__57_;
      r_71__56_ <= r_n_71__56_;
      r_71__55_ <= r_n_71__55_;
      r_71__54_ <= r_n_71__54_;
      r_71__53_ <= r_n_71__53_;
      r_71__52_ <= r_n_71__52_;
      r_71__51_ <= r_n_71__51_;
      r_71__50_ <= r_n_71__50_;
      r_71__49_ <= r_n_71__49_;
      r_71__48_ <= r_n_71__48_;
      r_71__47_ <= r_n_71__47_;
      r_71__46_ <= r_n_71__46_;
      r_71__45_ <= r_n_71__45_;
      r_71__44_ <= r_n_71__44_;
      r_71__43_ <= r_n_71__43_;
      r_71__42_ <= r_n_71__42_;
      r_71__41_ <= r_n_71__41_;
      r_71__40_ <= r_n_71__40_;
      r_71__39_ <= r_n_71__39_;
      r_71__38_ <= r_n_71__38_;
      r_71__37_ <= r_n_71__37_;
      r_71__36_ <= r_n_71__36_;
      r_71__35_ <= r_n_71__35_;
      r_71__34_ <= r_n_71__34_;
      r_71__33_ <= r_n_71__33_;
      r_71__32_ <= r_n_71__32_;
      r_71__31_ <= r_n_71__31_;
      r_71__30_ <= r_n_71__30_;
      r_71__29_ <= r_n_71__29_;
      r_71__28_ <= r_n_71__28_;
      r_71__27_ <= r_n_71__27_;
      r_71__26_ <= r_n_71__26_;
      r_71__25_ <= r_n_71__25_;
      r_71__24_ <= r_n_71__24_;
      r_71__23_ <= r_n_71__23_;
      r_71__22_ <= r_n_71__22_;
      r_71__21_ <= r_n_71__21_;
      r_71__20_ <= r_n_71__20_;
      r_71__19_ <= r_n_71__19_;
      r_71__18_ <= r_n_71__18_;
      r_71__17_ <= r_n_71__17_;
      r_71__16_ <= r_n_71__16_;
      r_71__15_ <= r_n_71__15_;
      r_71__14_ <= r_n_71__14_;
      r_71__13_ <= r_n_71__13_;
      r_71__12_ <= r_n_71__12_;
      r_71__11_ <= r_n_71__11_;
      r_71__10_ <= r_n_71__10_;
      r_71__9_ <= r_n_71__9_;
      r_71__8_ <= r_n_71__8_;
      r_71__7_ <= r_n_71__7_;
      r_71__6_ <= r_n_71__6_;
      r_71__5_ <= r_n_71__5_;
      r_71__4_ <= r_n_71__4_;
      r_71__3_ <= r_n_71__3_;
      r_71__2_ <= r_n_71__2_;
      r_71__1_ <= r_n_71__1_;
      r_71__0_ <= r_n_71__0_;
    end 
    if(N3656) begin
      r_72__63_ <= r_n_72__63_;
      r_72__62_ <= r_n_72__62_;
      r_72__61_ <= r_n_72__61_;
      r_72__60_ <= r_n_72__60_;
      r_72__59_ <= r_n_72__59_;
      r_72__58_ <= r_n_72__58_;
      r_72__57_ <= r_n_72__57_;
      r_72__56_ <= r_n_72__56_;
      r_72__55_ <= r_n_72__55_;
      r_72__54_ <= r_n_72__54_;
      r_72__53_ <= r_n_72__53_;
      r_72__52_ <= r_n_72__52_;
      r_72__51_ <= r_n_72__51_;
      r_72__50_ <= r_n_72__50_;
      r_72__49_ <= r_n_72__49_;
      r_72__48_ <= r_n_72__48_;
      r_72__47_ <= r_n_72__47_;
      r_72__46_ <= r_n_72__46_;
      r_72__45_ <= r_n_72__45_;
      r_72__44_ <= r_n_72__44_;
      r_72__43_ <= r_n_72__43_;
      r_72__42_ <= r_n_72__42_;
      r_72__41_ <= r_n_72__41_;
      r_72__40_ <= r_n_72__40_;
      r_72__39_ <= r_n_72__39_;
      r_72__38_ <= r_n_72__38_;
      r_72__37_ <= r_n_72__37_;
      r_72__36_ <= r_n_72__36_;
      r_72__35_ <= r_n_72__35_;
      r_72__34_ <= r_n_72__34_;
      r_72__33_ <= r_n_72__33_;
      r_72__32_ <= r_n_72__32_;
      r_72__31_ <= r_n_72__31_;
      r_72__30_ <= r_n_72__30_;
      r_72__29_ <= r_n_72__29_;
      r_72__28_ <= r_n_72__28_;
      r_72__27_ <= r_n_72__27_;
      r_72__26_ <= r_n_72__26_;
      r_72__25_ <= r_n_72__25_;
      r_72__24_ <= r_n_72__24_;
      r_72__23_ <= r_n_72__23_;
      r_72__22_ <= r_n_72__22_;
      r_72__21_ <= r_n_72__21_;
      r_72__20_ <= r_n_72__20_;
      r_72__19_ <= r_n_72__19_;
      r_72__18_ <= r_n_72__18_;
      r_72__17_ <= r_n_72__17_;
      r_72__16_ <= r_n_72__16_;
      r_72__15_ <= r_n_72__15_;
      r_72__14_ <= r_n_72__14_;
      r_72__13_ <= r_n_72__13_;
      r_72__12_ <= r_n_72__12_;
      r_72__11_ <= r_n_72__11_;
      r_72__10_ <= r_n_72__10_;
      r_72__9_ <= r_n_72__9_;
      r_72__8_ <= r_n_72__8_;
      r_72__7_ <= r_n_72__7_;
      r_72__6_ <= r_n_72__6_;
      r_72__5_ <= r_n_72__5_;
      r_72__4_ <= r_n_72__4_;
      r_72__3_ <= r_n_72__3_;
      r_72__2_ <= r_n_72__2_;
      r_72__1_ <= r_n_72__1_;
      r_72__0_ <= r_n_72__0_;
    end 
    if(N3657) begin
      r_73__63_ <= r_n_73__63_;
      r_73__62_ <= r_n_73__62_;
      r_73__61_ <= r_n_73__61_;
      r_73__60_ <= r_n_73__60_;
      r_73__59_ <= r_n_73__59_;
      r_73__58_ <= r_n_73__58_;
      r_73__57_ <= r_n_73__57_;
      r_73__56_ <= r_n_73__56_;
      r_73__55_ <= r_n_73__55_;
      r_73__54_ <= r_n_73__54_;
      r_73__53_ <= r_n_73__53_;
      r_73__52_ <= r_n_73__52_;
      r_73__51_ <= r_n_73__51_;
      r_73__50_ <= r_n_73__50_;
      r_73__49_ <= r_n_73__49_;
      r_73__48_ <= r_n_73__48_;
      r_73__47_ <= r_n_73__47_;
      r_73__46_ <= r_n_73__46_;
      r_73__45_ <= r_n_73__45_;
      r_73__44_ <= r_n_73__44_;
      r_73__43_ <= r_n_73__43_;
      r_73__42_ <= r_n_73__42_;
      r_73__41_ <= r_n_73__41_;
      r_73__40_ <= r_n_73__40_;
      r_73__39_ <= r_n_73__39_;
      r_73__38_ <= r_n_73__38_;
      r_73__37_ <= r_n_73__37_;
      r_73__36_ <= r_n_73__36_;
      r_73__35_ <= r_n_73__35_;
      r_73__34_ <= r_n_73__34_;
      r_73__33_ <= r_n_73__33_;
      r_73__32_ <= r_n_73__32_;
      r_73__31_ <= r_n_73__31_;
      r_73__30_ <= r_n_73__30_;
      r_73__29_ <= r_n_73__29_;
      r_73__28_ <= r_n_73__28_;
      r_73__27_ <= r_n_73__27_;
      r_73__26_ <= r_n_73__26_;
      r_73__25_ <= r_n_73__25_;
      r_73__24_ <= r_n_73__24_;
      r_73__23_ <= r_n_73__23_;
      r_73__22_ <= r_n_73__22_;
      r_73__21_ <= r_n_73__21_;
      r_73__20_ <= r_n_73__20_;
      r_73__19_ <= r_n_73__19_;
      r_73__18_ <= r_n_73__18_;
      r_73__17_ <= r_n_73__17_;
      r_73__16_ <= r_n_73__16_;
      r_73__15_ <= r_n_73__15_;
      r_73__14_ <= r_n_73__14_;
      r_73__13_ <= r_n_73__13_;
      r_73__12_ <= r_n_73__12_;
      r_73__11_ <= r_n_73__11_;
      r_73__10_ <= r_n_73__10_;
      r_73__9_ <= r_n_73__9_;
      r_73__8_ <= r_n_73__8_;
      r_73__7_ <= r_n_73__7_;
      r_73__6_ <= r_n_73__6_;
      r_73__5_ <= r_n_73__5_;
      r_73__4_ <= r_n_73__4_;
      r_73__3_ <= r_n_73__3_;
      r_73__2_ <= r_n_73__2_;
      r_73__1_ <= r_n_73__1_;
      r_73__0_ <= r_n_73__0_;
    end 
    if(N3658) begin
      r_74__63_ <= r_n_74__63_;
      r_74__62_ <= r_n_74__62_;
      r_74__61_ <= r_n_74__61_;
      r_74__60_ <= r_n_74__60_;
      r_74__59_ <= r_n_74__59_;
      r_74__58_ <= r_n_74__58_;
      r_74__57_ <= r_n_74__57_;
      r_74__56_ <= r_n_74__56_;
      r_74__55_ <= r_n_74__55_;
      r_74__54_ <= r_n_74__54_;
      r_74__53_ <= r_n_74__53_;
      r_74__52_ <= r_n_74__52_;
      r_74__51_ <= r_n_74__51_;
      r_74__50_ <= r_n_74__50_;
      r_74__49_ <= r_n_74__49_;
      r_74__48_ <= r_n_74__48_;
      r_74__47_ <= r_n_74__47_;
      r_74__46_ <= r_n_74__46_;
      r_74__45_ <= r_n_74__45_;
      r_74__44_ <= r_n_74__44_;
      r_74__43_ <= r_n_74__43_;
      r_74__42_ <= r_n_74__42_;
      r_74__41_ <= r_n_74__41_;
      r_74__40_ <= r_n_74__40_;
      r_74__39_ <= r_n_74__39_;
      r_74__38_ <= r_n_74__38_;
      r_74__37_ <= r_n_74__37_;
      r_74__36_ <= r_n_74__36_;
      r_74__35_ <= r_n_74__35_;
      r_74__34_ <= r_n_74__34_;
      r_74__33_ <= r_n_74__33_;
      r_74__32_ <= r_n_74__32_;
      r_74__31_ <= r_n_74__31_;
      r_74__30_ <= r_n_74__30_;
      r_74__29_ <= r_n_74__29_;
      r_74__28_ <= r_n_74__28_;
      r_74__27_ <= r_n_74__27_;
      r_74__26_ <= r_n_74__26_;
      r_74__25_ <= r_n_74__25_;
      r_74__24_ <= r_n_74__24_;
      r_74__23_ <= r_n_74__23_;
      r_74__22_ <= r_n_74__22_;
      r_74__21_ <= r_n_74__21_;
      r_74__20_ <= r_n_74__20_;
      r_74__19_ <= r_n_74__19_;
      r_74__18_ <= r_n_74__18_;
      r_74__17_ <= r_n_74__17_;
      r_74__16_ <= r_n_74__16_;
      r_74__15_ <= r_n_74__15_;
      r_74__14_ <= r_n_74__14_;
      r_74__13_ <= r_n_74__13_;
      r_74__12_ <= r_n_74__12_;
      r_74__11_ <= r_n_74__11_;
      r_74__10_ <= r_n_74__10_;
      r_74__9_ <= r_n_74__9_;
      r_74__8_ <= r_n_74__8_;
      r_74__7_ <= r_n_74__7_;
      r_74__6_ <= r_n_74__6_;
      r_74__5_ <= r_n_74__5_;
      r_74__4_ <= r_n_74__4_;
      r_74__3_ <= r_n_74__3_;
      r_74__2_ <= r_n_74__2_;
      r_74__1_ <= r_n_74__1_;
      r_74__0_ <= r_n_74__0_;
    end 
    if(N3659) begin
      r_75__63_ <= r_n_75__63_;
      r_75__62_ <= r_n_75__62_;
      r_75__61_ <= r_n_75__61_;
      r_75__60_ <= r_n_75__60_;
      r_75__59_ <= r_n_75__59_;
      r_75__58_ <= r_n_75__58_;
      r_75__57_ <= r_n_75__57_;
      r_75__56_ <= r_n_75__56_;
      r_75__55_ <= r_n_75__55_;
      r_75__54_ <= r_n_75__54_;
      r_75__53_ <= r_n_75__53_;
      r_75__52_ <= r_n_75__52_;
      r_75__51_ <= r_n_75__51_;
      r_75__50_ <= r_n_75__50_;
      r_75__49_ <= r_n_75__49_;
      r_75__48_ <= r_n_75__48_;
      r_75__47_ <= r_n_75__47_;
      r_75__46_ <= r_n_75__46_;
      r_75__45_ <= r_n_75__45_;
      r_75__44_ <= r_n_75__44_;
      r_75__43_ <= r_n_75__43_;
      r_75__42_ <= r_n_75__42_;
      r_75__41_ <= r_n_75__41_;
      r_75__40_ <= r_n_75__40_;
      r_75__39_ <= r_n_75__39_;
      r_75__38_ <= r_n_75__38_;
      r_75__37_ <= r_n_75__37_;
      r_75__36_ <= r_n_75__36_;
      r_75__35_ <= r_n_75__35_;
      r_75__34_ <= r_n_75__34_;
      r_75__33_ <= r_n_75__33_;
      r_75__32_ <= r_n_75__32_;
      r_75__31_ <= r_n_75__31_;
      r_75__30_ <= r_n_75__30_;
      r_75__29_ <= r_n_75__29_;
      r_75__28_ <= r_n_75__28_;
      r_75__27_ <= r_n_75__27_;
      r_75__26_ <= r_n_75__26_;
      r_75__25_ <= r_n_75__25_;
      r_75__24_ <= r_n_75__24_;
      r_75__23_ <= r_n_75__23_;
      r_75__22_ <= r_n_75__22_;
      r_75__21_ <= r_n_75__21_;
      r_75__20_ <= r_n_75__20_;
      r_75__19_ <= r_n_75__19_;
      r_75__18_ <= r_n_75__18_;
      r_75__17_ <= r_n_75__17_;
      r_75__16_ <= r_n_75__16_;
      r_75__15_ <= r_n_75__15_;
      r_75__14_ <= r_n_75__14_;
      r_75__13_ <= r_n_75__13_;
      r_75__12_ <= r_n_75__12_;
      r_75__11_ <= r_n_75__11_;
      r_75__10_ <= r_n_75__10_;
      r_75__9_ <= r_n_75__9_;
      r_75__8_ <= r_n_75__8_;
      r_75__7_ <= r_n_75__7_;
      r_75__6_ <= r_n_75__6_;
      r_75__5_ <= r_n_75__5_;
      r_75__4_ <= r_n_75__4_;
      r_75__3_ <= r_n_75__3_;
      r_75__2_ <= r_n_75__2_;
      r_75__1_ <= r_n_75__1_;
      r_75__0_ <= r_n_75__0_;
    end 
    if(N3660) begin
      r_76__63_ <= r_n_76__63_;
      r_76__62_ <= r_n_76__62_;
      r_76__61_ <= r_n_76__61_;
      r_76__60_ <= r_n_76__60_;
      r_76__59_ <= r_n_76__59_;
      r_76__58_ <= r_n_76__58_;
      r_76__57_ <= r_n_76__57_;
      r_76__56_ <= r_n_76__56_;
      r_76__55_ <= r_n_76__55_;
      r_76__54_ <= r_n_76__54_;
      r_76__53_ <= r_n_76__53_;
      r_76__52_ <= r_n_76__52_;
      r_76__51_ <= r_n_76__51_;
      r_76__50_ <= r_n_76__50_;
      r_76__49_ <= r_n_76__49_;
      r_76__48_ <= r_n_76__48_;
      r_76__47_ <= r_n_76__47_;
      r_76__46_ <= r_n_76__46_;
      r_76__45_ <= r_n_76__45_;
      r_76__44_ <= r_n_76__44_;
      r_76__43_ <= r_n_76__43_;
      r_76__42_ <= r_n_76__42_;
      r_76__41_ <= r_n_76__41_;
      r_76__40_ <= r_n_76__40_;
      r_76__39_ <= r_n_76__39_;
      r_76__38_ <= r_n_76__38_;
      r_76__37_ <= r_n_76__37_;
      r_76__36_ <= r_n_76__36_;
      r_76__35_ <= r_n_76__35_;
      r_76__34_ <= r_n_76__34_;
      r_76__33_ <= r_n_76__33_;
      r_76__32_ <= r_n_76__32_;
      r_76__31_ <= r_n_76__31_;
      r_76__30_ <= r_n_76__30_;
      r_76__29_ <= r_n_76__29_;
      r_76__28_ <= r_n_76__28_;
      r_76__27_ <= r_n_76__27_;
      r_76__26_ <= r_n_76__26_;
      r_76__25_ <= r_n_76__25_;
      r_76__24_ <= r_n_76__24_;
      r_76__23_ <= r_n_76__23_;
      r_76__22_ <= r_n_76__22_;
      r_76__21_ <= r_n_76__21_;
      r_76__20_ <= r_n_76__20_;
      r_76__19_ <= r_n_76__19_;
      r_76__18_ <= r_n_76__18_;
      r_76__17_ <= r_n_76__17_;
      r_76__16_ <= r_n_76__16_;
      r_76__15_ <= r_n_76__15_;
      r_76__14_ <= r_n_76__14_;
      r_76__13_ <= r_n_76__13_;
      r_76__12_ <= r_n_76__12_;
      r_76__11_ <= r_n_76__11_;
      r_76__10_ <= r_n_76__10_;
      r_76__9_ <= r_n_76__9_;
      r_76__8_ <= r_n_76__8_;
      r_76__7_ <= r_n_76__7_;
      r_76__6_ <= r_n_76__6_;
      r_76__5_ <= r_n_76__5_;
      r_76__4_ <= r_n_76__4_;
      r_76__3_ <= r_n_76__3_;
      r_76__2_ <= r_n_76__2_;
      r_76__1_ <= r_n_76__1_;
      r_76__0_ <= r_n_76__0_;
    end 
    if(N3661) begin
      r_77__63_ <= r_n_77__63_;
      r_77__62_ <= r_n_77__62_;
      r_77__61_ <= r_n_77__61_;
      r_77__60_ <= r_n_77__60_;
      r_77__59_ <= r_n_77__59_;
      r_77__58_ <= r_n_77__58_;
      r_77__57_ <= r_n_77__57_;
      r_77__56_ <= r_n_77__56_;
      r_77__55_ <= r_n_77__55_;
      r_77__54_ <= r_n_77__54_;
      r_77__53_ <= r_n_77__53_;
      r_77__52_ <= r_n_77__52_;
      r_77__51_ <= r_n_77__51_;
      r_77__50_ <= r_n_77__50_;
      r_77__49_ <= r_n_77__49_;
      r_77__48_ <= r_n_77__48_;
      r_77__47_ <= r_n_77__47_;
      r_77__46_ <= r_n_77__46_;
      r_77__45_ <= r_n_77__45_;
      r_77__44_ <= r_n_77__44_;
      r_77__43_ <= r_n_77__43_;
      r_77__42_ <= r_n_77__42_;
      r_77__41_ <= r_n_77__41_;
      r_77__40_ <= r_n_77__40_;
      r_77__39_ <= r_n_77__39_;
      r_77__38_ <= r_n_77__38_;
      r_77__37_ <= r_n_77__37_;
      r_77__36_ <= r_n_77__36_;
      r_77__35_ <= r_n_77__35_;
      r_77__34_ <= r_n_77__34_;
      r_77__33_ <= r_n_77__33_;
      r_77__32_ <= r_n_77__32_;
      r_77__31_ <= r_n_77__31_;
      r_77__30_ <= r_n_77__30_;
      r_77__29_ <= r_n_77__29_;
      r_77__28_ <= r_n_77__28_;
      r_77__27_ <= r_n_77__27_;
      r_77__26_ <= r_n_77__26_;
      r_77__25_ <= r_n_77__25_;
      r_77__24_ <= r_n_77__24_;
      r_77__23_ <= r_n_77__23_;
      r_77__22_ <= r_n_77__22_;
      r_77__21_ <= r_n_77__21_;
      r_77__20_ <= r_n_77__20_;
      r_77__19_ <= r_n_77__19_;
      r_77__18_ <= r_n_77__18_;
      r_77__17_ <= r_n_77__17_;
      r_77__16_ <= r_n_77__16_;
      r_77__15_ <= r_n_77__15_;
      r_77__14_ <= r_n_77__14_;
      r_77__13_ <= r_n_77__13_;
      r_77__12_ <= r_n_77__12_;
      r_77__11_ <= r_n_77__11_;
      r_77__10_ <= r_n_77__10_;
      r_77__9_ <= r_n_77__9_;
      r_77__8_ <= r_n_77__8_;
      r_77__7_ <= r_n_77__7_;
      r_77__6_ <= r_n_77__6_;
      r_77__5_ <= r_n_77__5_;
      r_77__4_ <= r_n_77__4_;
      r_77__3_ <= r_n_77__3_;
      r_77__2_ <= r_n_77__2_;
      r_77__1_ <= r_n_77__1_;
      r_77__0_ <= r_n_77__0_;
    end 
    if(N3662) begin
      r_78__63_ <= r_n_78__63_;
      r_78__62_ <= r_n_78__62_;
      r_78__61_ <= r_n_78__61_;
      r_78__60_ <= r_n_78__60_;
      r_78__59_ <= r_n_78__59_;
      r_78__58_ <= r_n_78__58_;
      r_78__57_ <= r_n_78__57_;
      r_78__56_ <= r_n_78__56_;
      r_78__55_ <= r_n_78__55_;
      r_78__54_ <= r_n_78__54_;
      r_78__53_ <= r_n_78__53_;
      r_78__52_ <= r_n_78__52_;
      r_78__51_ <= r_n_78__51_;
      r_78__50_ <= r_n_78__50_;
      r_78__49_ <= r_n_78__49_;
      r_78__48_ <= r_n_78__48_;
      r_78__47_ <= r_n_78__47_;
      r_78__46_ <= r_n_78__46_;
      r_78__45_ <= r_n_78__45_;
      r_78__44_ <= r_n_78__44_;
      r_78__43_ <= r_n_78__43_;
      r_78__42_ <= r_n_78__42_;
      r_78__41_ <= r_n_78__41_;
      r_78__40_ <= r_n_78__40_;
      r_78__39_ <= r_n_78__39_;
      r_78__38_ <= r_n_78__38_;
      r_78__37_ <= r_n_78__37_;
      r_78__36_ <= r_n_78__36_;
      r_78__35_ <= r_n_78__35_;
      r_78__34_ <= r_n_78__34_;
      r_78__33_ <= r_n_78__33_;
      r_78__32_ <= r_n_78__32_;
      r_78__31_ <= r_n_78__31_;
      r_78__30_ <= r_n_78__30_;
      r_78__29_ <= r_n_78__29_;
      r_78__28_ <= r_n_78__28_;
      r_78__27_ <= r_n_78__27_;
      r_78__26_ <= r_n_78__26_;
      r_78__25_ <= r_n_78__25_;
      r_78__24_ <= r_n_78__24_;
      r_78__23_ <= r_n_78__23_;
      r_78__22_ <= r_n_78__22_;
      r_78__21_ <= r_n_78__21_;
      r_78__20_ <= r_n_78__20_;
      r_78__19_ <= r_n_78__19_;
      r_78__18_ <= r_n_78__18_;
      r_78__17_ <= r_n_78__17_;
      r_78__16_ <= r_n_78__16_;
      r_78__15_ <= r_n_78__15_;
      r_78__14_ <= r_n_78__14_;
      r_78__13_ <= r_n_78__13_;
      r_78__12_ <= r_n_78__12_;
      r_78__11_ <= r_n_78__11_;
      r_78__10_ <= r_n_78__10_;
      r_78__9_ <= r_n_78__9_;
      r_78__8_ <= r_n_78__8_;
      r_78__7_ <= r_n_78__7_;
      r_78__6_ <= r_n_78__6_;
      r_78__5_ <= r_n_78__5_;
      r_78__4_ <= r_n_78__4_;
      r_78__3_ <= r_n_78__3_;
      r_78__2_ <= r_n_78__2_;
      r_78__1_ <= r_n_78__1_;
      r_78__0_ <= r_n_78__0_;
    end 
    if(N3663) begin
      r_79__63_ <= r_n_79__63_;
      r_79__62_ <= r_n_79__62_;
      r_79__61_ <= r_n_79__61_;
      r_79__60_ <= r_n_79__60_;
      r_79__59_ <= r_n_79__59_;
      r_79__58_ <= r_n_79__58_;
      r_79__57_ <= r_n_79__57_;
      r_79__56_ <= r_n_79__56_;
      r_79__55_ <= r_n_79__55_;
      r_79__54_ <= r_n_79__54_;
      r_79__53_ <= r_n_79__53_;
      r_79__52_ <= r_n_79__52_;
      r_79__51_ <= r_n_79__51_;
      r_79__50_ <= r_n_79__50_;
      r_79__49_ <= r_n_79__49_;
      r_79__48_ <= r_n_79__48_;
      r_79__47_ <= r_n_79__47_;
      r_79__46_ <= r_n_79__46_;
      r_79__45_ <= r_n_79__45_;
      r_79__44_ <= r_n_79__44_;
      r_79__43_ <= r_n_79__43_;
      r_79__42_ <= r_n_79__42_;
      r_79__41_ <= r_n_79__41_;
      r_79__40_ <= r_n_79__40_;
      r_79__39_ <= r_n_79__39_;
      r_79__38_ <= r_n_79__38_;
      r_79__37_ <= r_n_79__37_;
      r_79__36_ <= r_n_79__36_;
      r_79__35_ <= r_n_79__35_;
      r_79__34_ <= r_n_79__34_;
      r_79__33_ <= r_n_79__33_;
      r_79__32_ <= r_n_79__32_;
      r_79__31_ <= r_n_79__31_;
      r_79__30_ <= r_n_79__30_;
      r_79__29_ <= r_n_79__29_;
      r_79__28_ <= r_n_79__28_;
      r_79__27_ <= r_n_79__27_;
      r_79__26_ <= r_n_79__26_;
      r_79__25_ <= r_n_79__25_;
      r_79__24_ <= r_n_79__24_;
      r_79__23_ <= r_n_79__23_;
      r_79__22_ <= r_n_79__22_;
      r_79__21_ <= r_n_79__21_;
      r_79__20_ <= r_n_79__20_;
      r_79__19_ <= r_n_79__19_;
      r_79__18_ <= r_n_79__18_;
      r_79__17_ <= r_n_79__17_;
      r_79__16_ <= r_n_79__16_;
      r_79__15_ <= r_n_79__15_;
      r_79__14_ <= r_n_79__14_;
      r_79__13_ <= r_n_79__13_;
      r_79__12_ <= r_n_79__12_;
      r_79__11_ <= r_n_79__11_;
      r_79__10_ <= r_n_79__10_;
      r_79__9_ <= r_n_79__9_;
      r_79__8_ <= r_n_79__8_;
      r_79__7_ <= r_n_79__7_;
      r_79__6_ <= r_n_79__6_;
      r_79__5_ <= r_n_79__5_;
      r_79__4_ <= r_n_79__4_;
      r_79__3_ <= r_n_79__3_;
      r_79__2_ <= r_n_79__2_;
      r_79__1_ <= r_n_79__1_;
      r_79__0_ <= r_n_79__0_;
    end 
    if(N3664) begin
      r_80__63_ <= r_n_80__63_;
      r_80__62_ <= r_n_80__62_;
      r_80__61_ <= r_n_80__61_;
      r_80__60_ <= r_n_80__60_;
      r_80__59_ <= r_n_80__59_;
      r_80__58_ <= r_n_80__58_;
      r_80__57_ <= r_n_80__57_;
      r_80__56_ <= r_n_80__56_;
      r_80__55_ <= r_n_80__55_;
      r_80__54_ <= r_n_80__54_;
      r_80__53_ <= r_n_80__53_;
      r_80__52_ <= r_n_80__52_;
      r_80__51_ <= r_n_80__51_;
      r_80__50_ <= r_n_80__50_;
      r_80__49_ <= r_n_80__49_;
      r_80__48_ <= r_n_80__48_;
      r_80__47_ <= r_n_80__47_;
      r_80__46_ <= r_n_80__46_;
      r_80__45_ <= r_n_80__45_;
      r_80__44_ <= r_n_80__44_;
      r_80__43_ <= r_n_80__43_;
      r_80__42_ <= r_n_80__42_;
      r_80__41_ <= r_n_80__41_;
      r_80__40_ <= r_n_80__40_;
      r_80__39_ <= r_n_80__39_;
      r_80__38_ <= r_n_80__38_;
      r_80__37_ <= r_n_80__37_;
      r_80__36_ <= r_n_80__36_;
      r_80__35_ <= r_n_80__35_;
      r_80__34_ <= r_n_80__34_;
      r_80__33_ <= r_n_80__33_;
      r_80__32_ <= r_n_80__32_;
      r_80__31_ <= r_n_80__31_;
      r_80__30_ <= r_n_80__30_;
      r_80__29_ <= r_n_80__29_;
      r_80__28_ <= r_n_80__28_;
      r_80__27_ <= r_n_80__27_;
      r_80__26_ <= r_n_80__26_;
      r_80__25_ <= r_n_80__25_;
      r_80__24_ <= r_n_80__24_;
      r_80__23_ <= r_n_80__23_;
      r_80__22_ <= r_n_80__22_;
      r_80__21_ <= r_n_80__21_;
      r_80__20_ <= r_n_80__20_;
      r_80__19_ <= r_n_80__19_;
      r_80__18_ <= r_n_80__18_;
      r_80__17_ <= r_n_80__17_;
      r_80__16_ <= r_n_80__16_;
      r_80__15_ <= r_n_80__15_;
      r_80__14_ <= r_n_80__14_;
      r_80__13_ <= r_n_80__13_;
      r_80__12_ <= r_n_80__12_;
      r_80__11_ <= r_n_80__11_;
      r_80__10_ <= r_n_80__10_;
      r_80__9_ <= r_n_80__9_;
      r_80__8_ <= r_n_80__8_;
      r_80__7_ <= r_n_80__7_;
      r_80__6_ <= r_n_80__6_;
      r_80__5_ <= r_n_80__5_;
      r_80__4_ <= r_n_80__4_;
      r_80__3_ <= r_n_80__3_;
      r_80__2_ <= r_n_80__2_;
      r_80__1_ <= r_n_80__1_;
      r_80__0_ <= r_n_80__0_;
    end 
    if(N3665) begin
      r_81__63_ <= r_n_81__63_;
      r_81__62_ <= r_n_81__62_;
      r_81__61_ <= r_n_81__61_;
      r_81__60_ <= r_n_81__60_;
      r_81__59_ <= r_n_81__59_;
      r_81__58_ <= r_n_81__58_;
      r_81__57_ <= r_n_81__57_;
      r_81__56_ <= r_n_81__56_;
      r_81__55_ <= r_n_81__55_;
      r_81__54_ <= r_n_81__54_;
      r_81__53_ <= r_n_81__53_;
      r_81__52_ <= r_n_81__52_;
      r_81__51_ <= r_n_81__51_;
      r_81__50_ <= r_n_81__50_;
      r_81__49_ <= r_n_81__49_;
      r_81__48_ <= r_n_81__48_;
      r_81__47_ <= r_n_81__47_;
      r_81__46_ <= r_n_81__46_;
      r_81__45_ <= r_n_81__45_;
      r_81__44_ <= r_n_81__44_;
      r_81__43_ <= r_n_81__43_;
      r_81__42_ <= r_n_81__42_;
      r_81__41_ <= r_n_81__41_;
      r_81__40_ <= r_n_81__40_;
      r_81__39_ <= r_n_81__39_;
      r_81__38_ <= r_n_81__38_;
      r_81__37_ <= r_n_81__37_;
      r_81__36_ <= r_n_81__36_;
      r_81__35_ <= r_n_81__35_;
      r_81__34_ <= r_n_81__34_;
      r_81__33_ <= r_n_81__33_;
      r_81__32_ <= r_n_81__32_;
      r_81__31_ <= r_n_81__31_;
      r_81__30_ <= r_n_81__30_;
      r_81__29_ <= r_n_81__29_;
      r_81__28_ <= r_n_81__28_;
      r_81__27_ <= r_n_81__27_;
      r_81__26_ <= r_n_81__26_;
      r_81__25_ <= r_n_81__25_;
      r_81__24_ <= r_n_81__24_;
      r_81__23_ <= r_n_81__23_;
      r_81__22_ <= r_n_81__22_;
      r_81__21_ <= r_n_81__21_;
      r_81__20_ <= r_n_81__20_;
      r_81__19_ <= r_n_81__19_;
      r_81__18_ <= r_n_81__18_;
      r_81__17_ <= r_n_81__17_;
      r_81__16_ <= r_n_81__16_;
      r_81__15_ <= r_n_81__15_;
      r_81__14_ <= r_n_81__14_;
      r_81__13_ <= r_n_81__13_;
      r_81__12_ <= r_n_81__12_;
      r_81__11_ <= r_n_81__11_;
      r_81__10_ <= r_n_81__10_;
      r_81__9_ <= r_n_81__9_;
      r_81__8_ <= r_n_81__8_;
      r_81__7_ <= r_n_81__7_;
      r_81__6_ <= r_n_81__6_;
      r_81__5_ <= r_n_81__5_;
      r_81__4_ <= r_n_81__4_;
      r_81__3_ <= r_n_81__3_;
      r_81__2_ <= r_n_81__2_;
      r_81__1_ <= r_n_81__1_;
      r_81__0_ <= r_n_81__0_;
    end 
    if(N3666) begin
      r_82__63_ <= r_n_82__63_;
      r_82__62_ <= r_n_82__62_;
      r_82__61_ <= r_n_82__61_;
      r_82__60_ <= r_n_82__60_;
      r_82__59_ <= r_n_82__59_;
      r_82__58_ <= r_n_82__58_;
      r_82__57_ <= r_n_82__57_;
      r_82__56_ <= r_n_82__56_;
      r_82__55_ <= r_n_82__55_;
      r_82__54_ <= r_n_82__54_;
      r_82__53_ <= r_n_82__53_;
      r_82__52_ <= r_n_82__52_;
      r_82__51_ <= r_n_82__51_;
      r_82__50_ <= r_n_82__50_;
      r_82__49_ <= r_n_82__49_;
      r_82__48_ <= r_n_82__48_;
      r_82__47_ <= r_n_82__47_;
      r_82__46_ <= r_n_82__46_;
      r_82__45_ <= r_n_82__45_;
      r_82__44_ <= r_n_82__44_;
      r_82__43_ <= r_n_82__43_;
      r_82__42_ <= r_n_82__42_;
      r_82__41_ <= r_n_82__41_;
      r_82__40_ <= r_n_82__40_;
      r_82__39_ <= r_n_82__39_;
      r_82__38_ <= r_n_82__38_;
      r_82__37_ <= r_n_82__37_;
      r_82__36_ <= r_n_82__36_;
      r_82__35_ <= r_n_82__35_;
      r_82__34_ <= r_n_82__34_;
      r_82__33_ <= r_n_82__33_;
      r_82__32_ <= r_n_82__32_;
      r_82__31_ <= r_n_82__31_;
      r_82__30_ <= r_n_82__30_;
      r_82__29_ <= r_n_82__29_;
      r_82__28_ <= r_n_82__28_;
      r_82__27_ <= r_n_82__27_;
      r_82__26_ <= r_n_82__26_;
      r_82__25_ <= r_n_82__25_;
      r_82__24_ <= r_n_82__24_;
      r_82__23_ <= r_n_82__23_;
      r_82__22_ <= r_n_82__22_;
      r_82__21_ <= r_n_82__21_;
      r_82__20_ <= r_n_82__20_;
      r_82__19_ <= r_n_82__19_;
      r_82__18_ <= r_n_82__18_;
      r_82__17_ <= r_n_82__17_;
      r_82__16_ <= r_n_82__16_;
      r_82__15_ <= r_n_82__15_;
      r_82__14_ <= r_n_82__14_;
      r_82__13_ <= r_n_82__13_;
      r_82__12_ <= r_n_82__12_;
      r_82__11_ <= r_n_82__11_;
      r_82__10_ <= r_n_82__10_;
      r_82__9_ <= r_n_82__9_;
      r_82__8_ <= r_n_82__8_;
      r_82__7_ <= r_n_82__7_;
      r_82__6_ <= r_n_82__6_;
      r_82__5_ <= r_n_82__5_;
      r_82__4_ <= r_n_82__4_;
      r_82__3_ <= r_n_82__3_;
      r_82__2_ <= r_n_82__2_;
      r_82__1_ <= r_n_82__1_;
      r_82__0_ <= r_n_82__0_;
    end 
    if(N3667) begin
      r_83__63_ <= r_n_83__63_;
      r_83__62_ <= r_n_83__62_;
      r_83__61_ <= r_n_83__61_;
      r_83__60_ <= r_n_83__60_;
      r_83__59_ <= r_n_83__59_;
      r_83__58_ <= r_n_83__58_;
      r_83__57_ <= r_n_83__57_;
      r_83__56_ <= r_n_83__56_;
      r_83__55_ <= r_n_83__55_;
      r_83__54_ <= r_n_83__54_;
      r_83__53_ <= r_n_83__53_;
      r_83__52_ <= r_n_83__52_;
      r_83__51_ <= r_n_83__51_;
      r_83__50_ <= r_n_83__50_;
      r_83__49_ <= r_n_83__49_;
      r_83__48_ <= r_n_83__48_;
      r_83__47_ <= r_n_83__47_;
      r_83__46_ <= r_n_83__46_;
      r_83__45_ <= r_n_83__45_;
      r_83__44_ <= r_n_83__44_;
      r_83__43_ <= r_n_83__43_;
      r_83__42_ <= r_n_83__42_;
      r_83__41_ <= r_n_83__41_;
      r_83__40_ <= r_n_83__40_;
      r_83__39_ <= r_n_83__39_;
      r_83__38_ <= r_n_83__38_;
      r_83__37_ <= r_n_83__37_;
      r_83__36_ <= r_n_83__36_;
      r_83__35_ <= r_n_83__35_;
      r_83__34_ <= r_n_83__34_;
      r_83__33_ <= r_n_83__33_;
      r_83__32_ <= r_n_83__32_;
      r_83__31_ <= r_n_83__31_;
      r_83__30_ <= r_n_83__30_;
      r_83__29_ <= r_n_83__29_;
      r_83__28_ <= r_n_83__28_;
      r_83__27_ <= r_n_83__27_;
      r_83__26_ <= r_n_83__26_;
      r_83__25_ <= r_n_83__25_;
      r_83__24_ <= r_n_83__24_;
      r_83__23_ <= r_n_83__23_;
      r_83__22_ <= r_n_83__22_;
      r_83__21_ <= r_n_83__21_;
      r_83__20_ <= r_n_83__20_;
      r_83__19_ <= r_n_83__19_;
      r_83__18_ <= r_n_83__18_;
      r_83__17_ <= r_n_83__17_;
      r_83__16_ <= r_n_83__16_;
      r_83__15_ <= r_n_83__15_;
      r_83__14_ <= r_n_83__14_;
      r_83__13_ <= r_n_83__13_;
      r_83__12_ <= r_n_83__12_;
      r_83__11_ <= r_n_83__11_;
      r_83__10_ <= r_n_83__10_;
      r_83__9_ <= r_n_83__9_;
      r_83__8_ <= r_n_83__8_;
      r_83__7_ <= r_n_83__7_;
      r_83__6_ <= r_n_83__6_;
      r_83__5_ <= r_n_83__5_;
      r_83__4_ <= r_n_83__4_;
      r_83__3_ <= r_n_83__3_;
      r_83__2_ <= r_n_83__2_;
      r_83__1_ <= r_n_83__1_;
      r_83__0_ <= r_n_83__0_;
    end 
    if(N3668) begin
      r_84__63_ <= r_n_84__63_;
      r_84__62_ <= r_n_84__62_;
      r_84__61_ <= r_n_84__61_;
      r_84__60_ <= r_n_84__60_;
      r_84__59_ <= r_n_84__59_;
      r_84__58_ <= r_n_84__58_;
      r_84__57_ <= r_n_84__57_;
      r_84__56_ <= r_n_84__56_;
      r_84__55_ <= r_n_84__55_;
      r_84__54_ <= r_n_84__54_;
      r_84__53_ <= r_n_84__53_;
      r_84__52_ <= r_n_84__52_;
      r_84__51_ <= r_n_84__51_;
      r_84__50_ <= r_n_84__50_;
      r_84__49_ <= r_n_84__49_;
      r_84__48_ <= r_n_84__48_;
      r_84__47_ <= r_n_84__47_;
      r_84__46_ <= r_n_84__46_;
      r_84__45_ <= r_n_84__45_;
      r_84__44_ <= r_n_84__44_;
      r_84__43_ <= r_n_84__43_;
      r_84__42_ <= r_n_84__42_;
      r_84__41_ <= r_n_84__41_;
      r_84__40_ <= r_n_84__40_;
      r_84__39_ <= r_n_84__39_;
      r_84__38_ <= r_n_84__38_;
      r_84__37_ <= r_n_84__37_;
      r_84__36_ <= r_n_84__36_;
      r_84__35_ <= r_n_84__35_;
      r_84__34_ <= r_n_84__34_;
      r_84__33_ <= r_n_84__33_;
      r_84__32_ <= r_n_84__32_;
      r_84__31_ <= r_n_84__31_;
      r_84__30_ <= r_n_84__30_;
      r_84__29_ <= r_n_84__29_;
      r_84__28_ <= r_n_84__28_;
      r_84__27_ <= r_n_84__27_;
      r_84__26_ <= r_n_84__26_;
      r_84__25_ <= r_n_84__25_;
      r_84__24_ <= r_n_84__24_;
      r_84__23_ <= r_n_84__23_;
      r_84__22_ <= r_n_84__22_;
      r_84__21_ <= r_n_84__21_;
      r_84__20_ <= r_n_84__20_;
      r_84__19_ <= r_n_84__19_;
      r_84__18_ <= r_n_84__18_;
      r_84__17_ <= r_n_84__17_;
      r_84__16_ <= r_n_84__16_;
      r_84__15_ <= r_n_84__15_;
      r_84__14_ <= r_n_84__14_;
      r_84__13_ <= r_n_84__13_;
      r_84__12_ <= r_n_84__12_;
      r_84__11_ <= r_n_84__11_;
      r_84__10_ <= r_n_84__10_;
      r_84__9_ <= r_n_84__9_;
      r_84__8_ <= r_n_84__8_;
      r_84__7_ <= r_n_84__7_;
      r_84__6_ <= r_n_84__6_;
      r_84__5_ <= r_n_84__5_;
      r_84__4_ <= r_n_84__4_;
      r_84__3_ <= r_n_84__3_;
      r_84__2_ <= r_n_84__2_;
      r_84__1_ <= r_n_84__1_;
      r_84__0_ <= r_n_84__0_;
    end 
    if(N3669) begin
      r_85__63_ <= r_n_85__63_;
      r_85__62_ <= r_n_85__62_;
      r_85__61_ <= r_n_85__61_;
      r_85__60_ <= r_n_85__60_;
      r_85__59_ <= r_n_85__59_;
      r_85__58_ <= r_n_85__58_;
      r_85__57_ <= r_n_85__57_;
      r_85__56_ <= r_n_85__56_;
      r_85__55_ <= r_n_85__55_;
      r_85__54_ <= r_n_85__54_;
      r_85__53_ <= r_n_85__53_;
      r_85__52_ <= r_n_85__52_;
      r_85__51_ <= r_n_85__51_;
      r_85__50_ <= r_n_85__50_;
      r_85__49_ <= r_n_85__49_;
      r_85__48_ <= r_n_85__48_;
      r_85__47_ <= r_n_85__47_;
      r_85__46_ <= r_n_85__46_;
      r_85__45_ <= r_n_85__45_;
      r_85__44_ <= r_n_85__44_;
      r_85__43_ <= r_n_85__43_;
      r_85__42_ <= r_n_85__42_;
      r_85__41_ <= r_n_85__41_;
      r_85__40_ <= r_n_85__40_;
      r_85__39_ <= r_n_85__39_;
      r_85__38_ <= r_n_85__38_;
      r_85__37_ <= r_n_85__37_;
      r_85__36_ <= r_n_85__36_;
      r_85__35_ <= r_n_85__35_;
      r_85__34_ <= r_n_85__34_;
      r_85__33_ <= r_n_85__33_;
      r_85__32_ <= r_n_85__32_;
      r_85__31_ <= r_n_85__31_;
      r_85__30_ <= r_n_85__30_;
      r_85__29_ <= r_n_85__29_;
      r_85__28_ <= r_n_85__28_;
      r_85__27_ <= r_n_85__27_;
      r_85__26_ <= r_n_85__26_;
      r_85__25_ <= r_n_85__25_;
      r_85__24_ <= r_n_85__24_;
      r_85__23_ <= r_n_85__23_;
      r_85__22_ <= r_n_85__22_;
      r_85__21_ <= r_n_85__21_;
      r_85__20_ <= r_n_85__20_;
      r_85__19_ <= r_n_85__19_;
      r_85__18_ <= r_n_85__18_;
      r_85__17_ <= r_n_85__17_;
      r_85__16_ <= r_n_85__16_;
      r_85__15_ <= r_n_85__15_;
      r_85__14_ <= r_n_85__14_;
      r_85__13_ <= r_n_85__13_;
      r_85__12_ <= r_n_85__12_;
      r_85__11_ <= r_n_85__11_;
      r_85__10_ <= r_n_85__10_;
      r_85__9_ <= r_n_85__9_;
      r_85__8_ <= r_n_85__8_;
      r_85__7_ <= r_n_85__7_;
      r_85__6_ <= r_n_85__6_;
      r_85__5_ <= r_n_85__5_;
      r_85__4_ <= r_n_85__4_;
      r_85__3_ <= r_n_85__3_;
      r_85__2_ <= r_n_85__2_;
      r_85__1_ <= r_n_85__1_;
      r_85__0_ <= r_n_85__0_;
    end 
    if(N3670) begin
      r_86__63_ <= r_n_86__63_;
      r_86__62_ <= r_n_86__62_;
      r_86__61_ <= r_n_86__61_;
      r_86__60_ <= r_n_86__60_;
      r_86__59_ <= r_n_86__59_;
      r_86__58_ <= r_n_86__58_;
      r_86__57_ <= r_n_86__57_;
      r_86__56_ <= r_n_86__56_;
      r_86__55_ <= r_n_86__55_;
      r_86__54_ <= r_n_86__54_;
      r_86__53_ <= r_n_86__53_;
      r_86__52_ <= r_n_86__52_;
      r_86__51_ <= r_n_86__51_;
      r_86__50_ <= r_n_86__50_;
      r_86__49_ <= r_n_86__49_;
      r_86__48_ <= r_n_86__48_;
      r_86__47_ <= r_n_86__47_;
      r_86__46_ <= r_n_86__46_;
      r_86__45_ <= r_n_86__45_;
      r_86__44_ <= r_n_86__44_;
      r_86__43_ <= r_n_86__43_;
      r_86__42_ <= r_n_86__42_;
      r_86__41_ <= r_n_86__41_;
      r_86__40_ <= r_n_86__40_;
      r_86__39_ <= r_n_86__39_;
      r_86__38_ <= r_n_86__38_;
      r_86__37_ <= r_n_86__37_;
      r_86__36_ <= r_n_86__36_;
      r_86__35_ <= r_n_86__35_;
      r_86__34_ <= r_n_86__34_;
      r_86__33_ <= r_n_86__33_;
      r_86__32_ <= r_n_86__32_;
      r_86__31_ <= r_n_86__31_;
      r_86__30_ <= r_n_86__30_;
      r_86__29_ <= r_n_86__29_;
      r_86__28_ <= r_n_86__28_;
      r_86__27_ <= r_n_86__27_;
      r_86__26_ <= r_n_86__26_;
      r_86__25_ <= r_n_86__25_;
      r_86__24_ <= r_n_86__24_;
      r_86__23_ <= r_n_86__23_;
      r_86__22_ <= r_n_86__22_;
      r_86__21_ <= r_n_86__21_;
      r_86__20_ <= r_n_86__20_;
      r_86__19_ <= r_n_86__19_;
      r_86__18_ <= r_n_86__18_;
      r_86__17_ <= r_n_86__17_;
      r_86__16_ <= r_n_86__16_;
      r_86__15_ <= r_n_86__15_;
      r_86__14_ <= r_n_86__14_;
      r_86__13_ <= r_n_86__13_;
      r_86__12_ <= r_n_86__12_;
      r_86__11_ <= r_n_86__11_;
      r_86__10_ <= r_n_86__10_;
      r_86__9_ <= r_n_86__9_;
      r_86__8_ <= r_n_86__8_;
      r_86__7_ <= r_n_86__7_;
      r_86__6_ <= r_n_86__6_;
      r_86__5_ <= r_n_86__5_;
      r_86__4_ <= r_n_86__4_;
      r_86__3_ <= r_n_86__3_;
      r_86__2_ <= r_n_86__2_;
      r_86__1_ <= r_n_86__1_;
      r_86__0_ <= r_n_86__0_;
    end 
    if(N3671) begin
      r_87__63_ <= r_n_87__63_;
      r_87__62_ <= r_n_87__62_;
      r_87__61_ <= r_n_87__61_;
      r_87__60_ <= r_n_87__60_;
      r_87__59_ <= r_n_87__59_;
      r_87__58_ <= r_n_87__58_;
      r_87__57_ <= r_n_87__57_;
      r_87__56_ <= r_n_87__56_;
      r_87__55_ <= r_n_87__55_;
      r_87__54_ <= r_n_87__54_;
      r_87__53_ <= r_n_87__53_;
      r_87__52_ <= r_n_87__52_;
      r_87__51_ <= r_n_87__51_;
      r_87__50_ <= r_n_87__50_;
      r_87__49_ <= r_n_87__49_;
      r_87__48_ <= r_n_87__48_;
      r_87__47_ <= r_n_87__47_;
      r_87__46_ <= r_n_87__46_;
      r_87__45_ <= r_n_87__45_;
      r_87__44_ <= r_n_87__44_;
      r_87__43_ <= r_n_87__43_;
      r_87__42_ <= r_n_87__42_;
      r_87__41_ <= r_n_87__41_;
      r_87__40_ <= r_n_87__40_;
      r_87__39_ <= r_n_87__39_;
      r_87__38_ <= r_n_87__38_;
      r_87__37_ <= r_n_87__37_;
      r_87__36_ <= r_n_87__36_;
      r_87__35_ <= r_n_87__35_;
      r_87__34_ <= r_n_87__34_;
      r_87__33_ <= r_n_87__33_;
      r_87__32_ <= r_n_87__32_;
      r_87__31_ <= r_n_87__31_;
      r_87__30_ <= r_n_87__30_;
      r_87__29_ <= r_n_87__29_;
      r_87__28_ <= r_n_87__28_;
      r_87__27_ <= r_n_87__27_;
      r_87__26_ <= r_n_87__26_;
      r_87__25_ <= r_n_87__25_;
      r_87__24_ <= r_n_87__24_;
      r_87__23_ <= r_n_87__23_;
      r_87__22_ <= r_n_87__22_;
      r_87__21_ <= r_n_87__21_;
      r_87__20_ <= r_n_87__20_;
      r_87__19_ <= r_n_87__19_;
      r_87__18_ <= r_n_87__18_;
      r_87__17_ <= r_n_87__17_;
      r_87__16_ <= r_n_87__16_;
      r_87__15_ <= r_n_87__15_;
      r_87__14_ <= r_n_87__14_;
      r_87__13_ <= r_n_87__13_;
      r_87__12_ <= r_n_87__12_;
      r_87__11_ <= r_n_87__11_;
      r_87__10_ <= r_n_87__10_;
      r_87__9_ <= r_n_87__9_;
      r_87__8_ <= r_n_87__8_;
      r_87__7_ <= r_n_87__7_;
      r_87__6_ <= r_n_87__6_;
      r_87__5_ <= r_n_87__5_;
      r_87__4_ <= r_n_87__4_;
      r_87__3_ <= r_n_87__3_;
      r_87__2_ <= r_n_87__2_;
      r_87__1_ <= r_n_87__1_;
      r_87__0_ <= r_n_87__0_;
    end 
    if(N3672) begin
      r_88__63_ <= r_n_88__63_;
      r_88__62_ <= r_n_88__62_;
      r_88__61_ <= r_n_88__61_;
      r_88__60_ <= r_n_88__60_;
      r_88__59_ <= r_n_88__59_;
      r_88__58_ <= r_n_88__58_;
      r_88__57_ <= r_n_88__57_;
      r_88__56_ <= r_n_88__56_;
      r_88__55_ <= r_n_88__55_;
      r_88__54_ <= r_n_88__54_;
      r_88__53_ <= r_n_88__53_;
      r_88__52_ <= r_n_88__52_;
      r_88__51_ <= r_n_88__51_;
      r_88__50_ <= r_n_88__50_;
      r_88__49_ <= r_n_88__49_;
      r_88__48_ <= r_n_88__48_;
      r_88__47_ <= r_n_88__47_;
      r_88__46_ <= r_n_88__46_;
      r_88__45_ <= r_n_88__45_;
      r_88__44_ <= r_n_88__44_;
      r_88__43_ <= r_n_88__43_;
      r_88__42_ <= r_n_88__42_;
      r_88__41_ <= r_n_88__41_;
      r_88__40_ <= r_n_88__40_;
      r_88__39_ <= r_n_88__39_;
      r_88__38_ <= r_n_88__38_;
      r_88__37_ <= r_n_88__37_;
      r_88__36_ <= r_n_88__36_;
      r_88__35_ <= r_n_88__35_;
      r_88__34_ <= r_n_88__34_;
      r_88__33_ <= r_n_88__33_;
      r_88__32_ <= r_n_88__32_;
      r_88__31_ <= r_n_88__31_;
      r_88__30_ <= r_n_88__30_;
      r_88__29_ <= r_n_88__29_;
      r_88__28_ <= r_n_88__28_;
      r_88__27_ <= r_n_88__27_;
      r_88__26_ <= r_n_88__26_;
      r_88__25_ <= r_n_88__25_;
      r_88__24_ <= r_n_88__24_;
      r_88__23_ <= r_n_88__23_;
      r_88__22_ <= r_n_88__22_;
      r_88__21_ <= r_n_88__21_;
      r_88__20_ <= r_n_88__20_;
      r_88__19_ <= r_n_88__19_;
      r_88__18_ <= r_n_88__18_;
      r_88__17_ <= r_n_88__17_;
      r_88__16_ <= r_n_88__16_;
      r_88__15_ <= r_n_88__15_;
      r_88__14_ <= r_n_88__14_;
      r_88__13_ <= r_n_88__13_;
      r_88__12_ <= r_n_88__12_;
      r_88__11_ <= r_n_88__11_;
      r_88__10_ <= r_n_88__10_;
      r_88__9_ <= r_n_88__9_;
      r_88__8_ <= r_n_88__8_;
      r_88__7_ <= r_n_88__7_;
      r_88__6_ <= r_n_88__6_;
      r_88__5_ <= r_n_88__5_;
      r_88__4_ <= r_n_88__4_;
      r_88__3_ <= r_n_88__3_;
      r_88__2_ <= r_n_88__2_;
      r_88__1_ <= r_n_88__1_;
      r_88__0_ <= r_n_88__0_;
    end 
    if(N3673) begin
      r_89__63_ <= r_n_89__63_;
      r_89__62_ <= r_n_89__62_;
      r_89__61_ <= r_n_89__61_;
      r_89__60_ <= r_n_89__60_;
      r_89__59_ <= r_n_89__59_;
      r_89__58_ <= r_n_89__58_;
      r_89__57_ <= r_n_89__57_;
      r_89__56_ <= r_n_89__56_;
      r_89__55_ <= r_n_89__55_;
      r_89__54_ <= r_n_89__54_;
      r_89__53_ <= r_n_89__53_;
      r_89__52_ <= r_n_89__52_;
      r_89__51_ <= r_n_89__51_;
      r_89__50_ <= r_n_89__50_;
      r_89__49_ <= r_n_89__49_;
      r_89__48_ <= r_n_89__48_;
      r_89__47_ <= r_n_89__47_;
      r_89__46_ <= r_n_89__46_;
      r_89__45_ <= r_n_89__45_;
      r_89__44_ <= r_n_89__44_;
      r_89__43_ <= r_n_89__43_;
      r_89__42_ <= r_n_89__42_;
      r_89__41_ <= r_n_89__41_;
      r_89__40_ <= r_n_89__40_;
      r_89__39_ <= r_n_89__39_;
      r_89__38_ <= r_n_89__38_;
      r_89__37_ <= r_n_89__37_;
      r_89__36_ <= r_n_89__36_;
      r_89__35_ <= r_n_89__35_;
      r_89__34_ <= r_n_89__34_;
      r_89__33_ <= r_n_89__33_;
      r_89__32_ <= r_n_89__32_;
      r_89__31_ <= r_n_89__31_;
      r_89__30_ <= r_n_89__30_;
      r_89__29_ <= r_n_89__29_;
      r_89__28_ <= r_n_89__28_;
      r_89__27_ <= r_n_89__27_;
      r_89__26_ <= r_n_89__26_;
      r_89__25_ <= r_n_89__25_;
      r_89__24_ <= r_n_89__24_;
      r_89__23_ <= r_n_89__23_;
      r_89__22_ <= r_n_89__22_;
      r_89__21_ <= r_n_89__21_;
      r_89__20_ <= r_n_89__20_;
      r_89__19_ <= r_n_89__19_;
      r_89__18_ <= r_n_89__18_;
      r_89__17_ <= r_n_89__17_;
      r_89__16_ <= r_n_89__16_;
      r_89__15_ <= r_n_89__15_;
      r_89__14_ <= r_n_89__14_;
      r_89__13_ <= r_n_89__13_;
      r_89__12_ <= r_n_89__12_;
      r_89__11_ <= r_n_89__11_;
      r_89__10_ <= r_n_89__10_;
      r_89__9_ <= r_n_89__9_;
      r_89__8_ <= r_n_89__8_;
      r_89__7_ <= r_n_89__7_;
      r_89__6_ <= r_n_89__6_;
      r_89__5_ <= r_n_89__5_;
      r_89__4_ <= r_n_89__4_;
      r_89__3_ <= r_n_89__3_;
      r_89__2_ <= r_n_89__2_;
      r_89__1_ <= r_n_89__1_;
      r_89__0_ <= r_n_89__0_;
    end 
    if(N3674) begin
      r_90__63_ <= r_n_90__63_;
      r_90__62_ <= r_n_90__62_;
      r_90__61_ <= r_n_90__61_;
      r_90__60_ <= r_n_90__60_;
      r_90__59_ <= r_n_90__59_;
      r_90__58_ <= r_n_90__58_;
      r_90__57_ <= r_n_90__57_;
      r_90__56_ <= r_n_90__56_;
      r_90__55_ <= r_n_90__55_;
      r_90__54_ <= r_n_90__54_;
      r_90__53_ <= r_n_90__53_;
      r_90__52_ <= r_n_90__52_;
      r_90__51_ <= r_n_90__51_;
      r_90__50_ <= r_n_90__50_;
      r_90__49_ <= r_n_90__49_;
      r_90__48_ <= r_n_90__48_;
      r_90__47_ <= r_n_90__47_;
      r_90__46_ <= r_n_90__46_;
      r_90__45_ <= r_n_90__45_;
      r_90__44_ <= r_n_90__44_;
      r_90__43_ <= r_n_90__43_;
      r_90__42_ <= r_n_90__42_;
      r_90__41_ <= r_n_90__41_;
      r_90__40_ <= r_n_90__40_;
      r_90__39_ <= r_n_90__39_;
      r_90__38_ <= r_n_90__38_;
      r_90__37_ <= r_n_90__37_;
      r_90__36_ <= r_n_90__36_;
      r_90__35_ <= r_n_90__35_;
      r_90__34_ <= r_n_90__34_;
      r_90__33_ <= r_n_90__33_;
      r_90__32_ <= r_n_90__32_;
      r_90__31_ <= r_n_90__31_;
      r_90__30_ <= r_n_90__30_;
      r_90__29_ <= r_n_90__29_;
      r_90__28_ <= r_n_90__28_;
      r_90__27_ <= r_n_90__27_;
      r_90__26_ <= r_n_90__26_;
      r_90__25_ <= r_n_90__25_;
      r_90__24_ <= r_n_90__24_;
      r_90__23_ <= r_n_90__23_;
      r_90__22_ <= r_n_90__22_;
      r_90__21_ <= r_n_90__21_;
      r_90__20_ <= r_n_90__20_;
      r_90__19_ <= r_n_90__19_;
      r_90__18_ <= r_n_90__18_;
      r_90__17_ <= r_n_90__17_;
      r_90__16_ <= r_n_90__16_;
      r_90__15_ <= r_n_90__15_;
      r_90__14_ <= r_n_90__14_;
      r_90__13_ <= r_n_90__13_;
      r_90__12_ <= r_n_90__12_;
      r_90__11_ <= r_n_90__11_;
      r_90__10_ <= r_n_90__10_;
      r_90__9_ <= r_n_90__9_;
      r_90__8_ <= r_n_90__8_;
      r_90__7_ <= r_n_90__7_;
      r_90__6_ <= r_n_90__6_;
      r_90__5_ <= r_n_90__5_;
      r_90__4_ <= r_n_90__4_;
      r_90__3_ <= r_n_90__3_;
      r_90__2_ <= r_n_90__2_;
      r_90__1_ <= r_n_90__1_;
      r_90__0_ <= r_n_90__0_;
    end 
    if(N3675) begin
      r_91__63_ <= r_n_91__63_;
      r_91__62_ <= r_n_91__62_;
      r_91__61_ <= r_n_91__61_;
      r_91__60_ <= r_n_91__60_;
      r_91__59_ <= r_n_91__59_;
      r_91__58_ <= r_n_91__58_;
      r_91__57_ <= r_n_91__57_;
      r_91__56_ <= r_n_91__56_;
      r_91__55_ <= r_n_91__55_;
      r_91__54_ <= r_n_91__54_;
      r_91__53_ <= r_n_91__53_;
      r_91__52_ <= r_n_91__52_;
      r_91__51_ <= r_n_91__51_;
      r_91__50_ <= r_n_91__50_;
      r_91__49_ <= r_n_91__49_;
      r_91__48_ <= r_n_91__48_;
      r_91__47_ <= r_n_91__47_;
      r_91__46_ <= r_n_91__46_;
      r_91__45_ <= r_n_91__45_;
      r_91__44_ <= r_n_91__44_;
      r_91__43_ <= r_n_91__43_;
      r_91__42_ <= r_n_91__42_;
      r_91__41_ <= r_n_91__41_;
      r_91__40_ <= r_n_91__40_;
      r_91__39_ <= r_n_91__39_;
      r_91__38_ <= r_n_91__38_;
      r_91__37_ <= r_n_91__37_;
      r_91__36_ <= r_n_91__36_;
      r_91__35_ <= r_n_91__35_;
      r_91__34_ <= r_n_91__34_;
      r_91__33_ <= r_n_91__33_;
      r_91__32_ <= r_n_91__32_;
      r_91__31_ <= r_n_91__31_;
      r_91__30_ <= r_n_91__30_;
      r_91__29_ <= r_n_91__29_;
      r_91__28_ <= r_n_91__28_;
      r_91__27_ <= r_n_91__27_;
      r_91__26_ <= r_n_91__26_;
      r_91__25_ <= r_n_91__25_;
      r_91__24_ <= r_n_91__24_;
      r_91__23_ <= r_n_91__23_;
      r_91__22_ <= r_n_91__22_;
      r_91__21_ <= r_n_91__21_;
      r_91__20_ <= r_n_91__20_;
      r_91__19_ <= r_n_91__19_;
      r_91__18_ <= r_n_91__18_;
      r_91__17_ <= r_n_91__17_;
      r_91__16_ <= r_n_91__16_;
      r_91__15_ <= r_n_91__15_;
      r_91__14_ <= r_n_91__14_;
      r_91__13_ <= r_n_91__13_;
      r_91__12_ <= r_n_91__12_;
      r_91__11_ <= r_n_91__11_;
      r_91__10_ <= r_n_91__10_;
      r_91__9_ <= r_n_91__9_;
      r_91__8_ <= r_n_91__8_;
      r_91__7_ <= r_n_91__7_;
      r_91__6_ <= r_n_91__6_;
      r_91__5_ <= r_n_91__5_;
      r_91__4_ <= r_n_91__4_;
      r_91__3_ <= r_n_91__3_;
      r_91__2_ <= r_n_91__2_;
      r_91__1_ <= r_n_91__1_;
      r_91__0_ <= r_n_91__0_;
    end 
    if(N3676) begin
      r_92__63_ <= r_n_92__63_;
      r_92__62_ <= r_n_92__62_;
      r_92__61_ <= r_n_92__61_;
      r_92__60_ <= r_n_92__60_;
      r_92__59_ <= r_n_92__59_;
      r_92__58_ <= r_n_92__58_;
      r_92__57_ <= r_n_92__57_;
      r_92__56_ <= r_n_92__56_;
      r_92__55_ <= r_n_92__55_;
      r_92__54_ <= r_n_92__54_;
      r_92__53_ <= r_n_92__53_;
      r_92__52_ <= r_n_92__52_;
      r_92__51_ <= r_n_92__51_;
      r_92__50_ <= r_n_92__50_;
      r_92__49_ <= r_n_92__49_;
      r_92__48_ <= r_n_92__48_;
      r_92__47_ <= r_n_92__47_;
      r_92__46_ <= r_n_92__46_;
      r_92__45_ <= r_n_92__45_;
      r_92__44_ <= r_n_92__44_;
      r_92__43_ <= r_n_92__43_;
      r_92__42_ <= r_n_92__42_;
      r_92__41_ <= r_n_92__41_;
      r_92__40_ <= r_n_92__40_;
      r_92__39_ <= r_n_92__39_;
      r_92__38_ <= r_n_92__38_;
      r_92__37_ <= r_n_92__37_;
      r_92__36_ <= r_n_92__36_;
      r_92__35_ <= r_n_92__35_;
      r_92__34_ <= r_n_92__34_;
      r_92__33_ <= r_n_92__33_;
      r_92__32_ <= r_n_92__32_;
      r_92__31_ <= r_n_92__31_;
      r_92__30_ <= r_n_92__30_;
      r_92__29_ <= r_n_92__29_;
      r_92__28_ <= r_n_92__28_;
      r_92__27_ <= r_n_92__27_;
      r_92__26_ <= r_n_92__26_;
      r_92__25_ <= r_n_92__25_;
      r_92__24_ <= r_n_92__24_;
      r_92__23_ <= r_n_92__23_;
      r_92__22_ <= r_n_92__22_;
      r_92__21_ <= r_n_92__21_;
      r_92__20_ <= r_n_92__20_;
      r_92__19_ <= r_n_92__19_;
      r_92__18_ <= r_n_92__18_;
      r_92__17_ <= r_n_92__17_;
      r_92__16_ <= r_n_92__16_;
      r_92__15_ <= r_n_92__15_;
      r_92__14_ <= r_n_92__14_;
      r_92__13_ <= r_n_92__13_;
      r_92__12_ <= r_n_92__12_;
      r_92__11_ <= r_n_92__11_;
      r_92__10_ <= r_n_92__10_;
      r_92__9_ <= r_n_92__9_;
      r_92__8_ <= r_n_92__8_;
      r_92__7_ <= r_n_92__7_;
      r_92__6_ <= r_n_92__6_;
      r_92__5_ <= r_n_92__5_;
      r_92__4_ <= r_n_92__4_;
      r_92__3_ <= r_n_92__3_;
      r_92__2_ <= r_n_92__2_;
      r_92__1_ <= r_n_92__1_;
      r_92__0_ <= r_n_92__0_;
    end 
    if(N3677) begin
      r_93__63_ <= r_n_93__63_;
      r_93__62_ <= r_n_93__62_;
      r_93__61_ <= r_n_93__61_;
      r_93__60_ <= r_n_93__60_;
      r_93__59_ <= r_n_93__59_;
      r_93__58_ <= r_n_93__58_;
      r_93__57_ <= r_n_93__57_;
      r_93__56_ <= r_n_93__56_;
      r_93__55_ <= r_n_93__55_;
      r_93__54_ <= r_n_93__54_;
      r_93__53_ <= r_n_93__53_;
      r_93__52_ <= r_n_93__52_;
      r_93__51_ <= r_n_93__51_;
      r_93__50_ <= r_n_93__50_;
      r_93__49_ <= r_n_93__49_;
      r_93__48_ <= r_n_93__48_;
      r_93__47_ <= r_n_93__47_;
      r_93__46_ <= r_n_93__46_;
      r_93__45_ <= r_n_93__45_;
      r_93__44_ <= r_n_93__44_;
      r_93__43_ <= r_n_93__43_;
      r_93__42_ <= r_n_93__42_;
      r_93__41_ <= r_n_93__41_;
      r_93__40_ <= r_n_93__40_;
      r_93__39_ <= r_n_93__39_;
      r_93__38_ <= r_n_93__38_;
      r_93__37_ <= r_n_93__37_;
      r_93__36_ <= r_n_93__36_;
      r_93__35_ <= r_n_93__35_;
      r_93__34_ <= r_n_93__34_;
      r_93__33_ <= r_n_93__33_;
      r_93__32_ <= r_n_93__32_;
      r_93__31_ <= r_n_93__31_;
      r_93__30_ <= r_n_93__30_;
      r_93__29_ <= r_n_93__29_;
      r_93__28_ <= r_n_93__28_;
      r_93__27_ <= r_n_93__27_;
      r_93__26_ <= r_n_93__26_;
      r_93__25_ <= r_n_93__25_;
      r_93__24_ <= r_n_93__24_;
      r_93__23_ <= r_n_93__23_;
      r_93__22_ <= r_n_93__22_;
      r_93__21_ <= r_n_93__21_;
      r_93__20_ <= r_n_93__20_;
      r_93__19_ <= r_n_93__19_;
      r_93__18_ <= r_n_93__18_;
      r_93__17_ <= r_n_93__17_;
      r_93__16_ <= r_n_93__16_;
      r_93__15_ <= r_n_93__15_;
      r_93__14_ <= r_n_93__14_;
      r_93__13_ <= r_n_93__13_;
      r_93__12_ <= r_n_93__12_;
      r_93__11_ <= r_n_93__11_;
      r_93__10_ <= r_n_93__10_;
      r_93__9_ <= r_n_93__9_;
      r_93__8_ <= r_n_93__8_;
      r_93__7_ <= r_n_93__7_;
      r_93__6_ <= r_n_93__6_;
      r_93__5_ <= r_n_93__5_;
      r_93__4_ <= r_n_93__4_;
      r_93__3_ <= r_n_93__3_;
      r_93__2_ <= r_n_93__2_;
      r_93__1_ <= r_n_93__1_;
      r_93__0_ <= r_n_93__0_;
    end 
    if(N3678) begin
      r_94__63_ <= r_n_94__63_;
      r_94__62_ <= r_n_94__62_;
      r_94__61_ <= r_n_94__61_;
      r_94__60_ <= r_n_94__60_;
      r_94__59_ <= r_n_94__59_;
      r_94__58_ <= r_n_94__58_;
      r_94__57_ <= r_n_94__57_;
      r_94__56_ <= r_n_94__56_;
      r_94__55_ <= r_n_94__55_;
      r_94__54_ <= r_n_94__54_;
      r_94__53_ <= r_n_94__53_;
      r_94__52_ <= r_n_94__52_;
      r_94__51_ <= r_n_94__51_;
      r_94__50_ <= r_n_94__50_;
      r_94__49_ <= r_n_94__49_;
      r_94__48_ <= r_n_94__48_;
      r_94__47_ <= r_n_94__47_;
      r_94__46_ <= r_n_94__46_;
      r_94__45_ <= r_n_94__45_;
      r_94__44_ <= r_n_94__44_;
      r_94__43_ <= r_n_94__43_;
      r_94__42_ <= r_n_94__42_;
      r_94__41_ <= r_n_94__41_;
      r_94__40_ <= r_n_94__40_;
      r_94__39_ <= r_n_94__39_;
      r_94__38_ <= r_n_94__38_;
      r_94__37_ <= r_n_94__37_;
      r_94__36_ <= r_n_94__36_;
      r_94__35_ <= r_n_94__35_;
      r_94__34_ <= r_n_94__34_;
      r_94__33_ <= r_n_94__33_;
      r_94__32_ <= r_n_94__32_;
      r_94__31_ <= r_n_94__31_;
      r_94__30_ <= r_n_94__30_;
      r_94__29_ <= r_n_94__29_;
      r_94__28_ <= r_n_94__28_;
      r_94__27_ <= r_n_94__27_;
      r_94__26_ <= r_n_94__26_;
      r_94__25_ <= r_n_94__25_;
      r_94__24_ <= r_n_94__24_;
      r_94__23_ <= r_n_94__23_;
      r_94__22_ <= r_n_94__22_;
      r_94__21_ <= r_n_94__21_;
      r_94__20_ <= r_n_94__20_;
      r_94__19_ <= r_n_94__19_;
      r_94__18_ <= r_n_94__18_;
      r_94__17_ <= r_n_94__17_;
      r_94__16_ <= r_n_94__16_;
      r_94__15_ <= r_n_94__15_;
      r_94__14_ <= r_n_94__14_;
      r_94__13_ <= r_n_94__13_;
      r_94__12_ <= r_n_94__12_;
      r_94__11_ <= r_n_94__11_;
      r_94__10_ <= r_n_94__10_;
      r_94__9_ <= r_n_94__9_;
      r_94__8_ <= r_n_94__8_;
      r_94__7_ <= r_n_94__7_;
      r_94__6_ <= r_n_94__6_;
      r_94__5_ <= r_n_94__5_;
      r_94__4_ <= r_n_94__4_;
      r_94__3_ <= r_n_94__3_;
      r_94__2_ <= r_n_94__2_;
      r_94__1_ <= r_n_94__1_;
      r_94__0_ <= r_n_94__0_;
    end 
    if(N3679) begin
      r_95__63_ <= r_n_95__63_;
      r_95__62_ <= r_n_95__62_;
      r_95__61_ <= r_n_95__61_;
      r_95__60_ <= r_n_95__60_;
      r_95__59_ <= r_n_95__59_;
      r_95__58_ <= r_n_95__58_;
      r_95__57_ <= r_n_95__57_;
      r_95__56_ <= r_n_95__56_;
      r_95__55_ <= r_n_95__55_;
      r_95__54_ <= r_n_95__54_;
      r_95__53_ <= r_n_95__53_;
      r_95__52_ <= r_n_95__52_;
      r_95__51_ <= r_n_95__51_;
      r_95__50_ <= r_n_95__50_;
      r_95__49_ <= r_n_95__49_;
      r_95__48_ <= r_n_95__48_;
      r_95__47_ <= r_n_95__47_;
      r_95__46_ <= r_n_95__46_;
      r_95__45_ <= r_n_95__45_;
      r_95__44_ <= r_n_95__44_;
      r_95__43_ <= r_n_95__43_;
      r_95__42_ <= r_n_95__42_;
      r_95__41_ <= r_n_95__41_;
      r_95__40_ <= r_n_95__40_;
      r_95__39_ <= r_n_95__39_;
      r_95__38_ <= r_n_95__38_;
      r_95__37_ <= r_n_95__37_;
      r_95__36_ <= r_n_95__36_;
      r_95__35_ <= r_n_95__35_;
      r_95__34_ <= r_n_95__34_;
      r_95__33_ <= r_n_95__33_;
      r_95__32_ <= r_n_95__32_;
      r_95__31_ <= r_n_95__31_;
      r_95__30_ <= r_n_95__30_;
      r_95__29_ <= r_n_95__29_;
      r_95__28_ <= r_n_95__28_;
      r_95__27_ <= r_n_95__27_;
      r_95__26_ <= r_n_95__26_;
      r_95__25_ <= r_n_95__25_;
      r_95__24_ <= r_n_95__24_;
      r_95__23_ <= r_n_95__23_;
      r_95__22_ <= r_n_95__22_;
      r_95__21_ <= r_n_95__21_;
      r_95__20_ <= r_n_95__20_;
      r_95__19_ <= r_n_95__19_;
      r_95__18_ <= r_n_95__18_;
      r_95__17_ <= r_n_95__17_;
      r_95__16_ <= r_n_95__16_;
      r_95__15_ <= r_n_95__15_;
      r_95__14_ <= r_n_95__14_;
      r_95__13_ <= r_n_95__13_;
      r_95__12_ <= r_n_95__12_;
      r_95__11_ <= r_n_95__11_;
      r_95__10_ <= r_n_95__10_;
      r_95__9_ <= r_n_95__9_;
      r_95__8_ <= r_n_95__8_;
      r_95__7_ <= r_n_95__7_;
      r_95__6_ <= r_n_95__6_;
      r_95__5_ <= r_n_95__5_;
      r_95__4_ <= r_n_95__4_;
      r_95__3_ <= r_n_95__3_;
      r_95__2_ <= r_n_95__2_;
      r_95__1_ <= r_n_95__1_;
      r_95__0_ <= r_n_95__0_;
    end 
    if(N3680) begin
      r_96__63_ <= r_n_96__63_;
      r_96__62_ <= r_n_96__62_;
      r_96__61_ <= r_n_96__61_;
      r_96__60_ <= r_n_96__60_;
      r_96__59_ <= r_n_96__59_;
      r_96__58_ <= r_n_96__58_;
      r_96__57_ <= r_n_96__57_;
      r_96__56_ <= r_n_96__56_;
      r_96__55_ <= r_n_96__55_;
      r_96__54_ <= r_n_96__54_;
      r_96__53_ <= r_n_96__53_;
      r_96__52_ <= r_n_96__52_;
      r_96__51_ <= r_n_96__51_;
      r_96__50_ <= r_n_96__50_;
      r_96__49_ <= r_n_96__49_;
      r_96__48_ <= r_n_96__48_;
      r_96__47_ <= r_n_96__47_;
      r_96__46_ <= r_n_96__46_;
      r_96__45_ <= r_n_96__45_;
      r_96__44_ <= r_n_96__44_;
      r_96__43_ <= r_n_96__43_;
      r_96__42_ <= r_n_96__42_;
      r_96__41_ <= r_n_96__41_;
      r_96__40_ <= r_n_96__40_;
      r_96__39_ <= r_n_96__39_;
      r_96__38_ <= r_n_96__38_;
      r_96__37_ <= r_n_96__37_;
      r_96__36_ <= r_n_96__36_;
      r_96__35_ <= r_n_96__35_;
      r_96__34_ <= r_n_96__34_;
      r_96__33_ <= r_n_96__33_;
      r_96__32_ <= r_n_96__32_;
      r_96__31_ <= r_n_96__31_;
      r_96__30_ <= r_n_96__30_;
      r_96__29_ <= r_n_96__29_;
      r_96__28_ <= r_n_96__28_;
      r_96__27_ <= r_n_96__27_;
      r_96__26_ <= r_n_96__26_;
      r_96__25_ <= r_n_96__25_;
      r_96__24_ <= r_n_96__24_;
      r_96__23_ <= r_n_96__23_;
      r_96__22_ <= r_n_96__22_;
      r_96__21_ <= r_n_96__21_;
      r_96__20_ <= r_n_96__20_;
      r_96__19_ <= r_n_96__19_;
      r_96__18_ <= r_n_96__18_;
      r_96__17_ <= r_n_96__17_;
      r_96__16_ <= r_n_96__16_;
      r_96__15_ <= r_n_96__15_;
      r_96__14_ <= r_n_96__14_;
      r_96__13_ <= r_n_96__13_;
      r_96__12_ <= r_n_96__12_;
      r_96__11_ <= r_n_96__11_;
      r_96__10_ <= r_n_96__10_;
      r_96__9_ <= r_n_96__9_;
      r_96__8_ <= r_n_96__8_;
      r_96__7_ <= r_n_96__7_;
      r_96__6_ <= r_n_96__6_;
      r_96__5_ <= r_n_96__5_;
      r_96__4_ <= r_n_96__4_;
      r_96__3_ <= r_n_96__3_;
      r_96__2_ <= r_n_96__2_;
      r_96__1_ <= r_n_96__1_;
      r_96__0_ <= r_n_96__0_;
    end 
    if(N3681) begin
      r_97__63_ <= r_n_97__63_;
      r_97__62_ <= r_n_97__62_;
      r_97__61_ <= r_n_97__61_;
      r_97__60_ <= r_n_97__60_;
      r_97__59_ <= r_n_97__59_;
      r_97__58_ <= r_n_97__58_;
      r_97__57_ <= r_n_97__57_;
      r_97__56_ <= r_n_97__56_;
      r_97__55_ <= r_n_97__55_;
      r_97__54_ <= r_n_97__54_;
      r_97__53_ <= r_n_97__53_;
      r_97__52_ <= r_n_97__52_;
      r_97__51_ <= r_n_97__51_;
      r_97__50_ <= r_n_97__50_;
      r_97__49_ <= r_n_97__49_;
      r_97__48_ <= r_n_97__48_;
      r_97__47_ <= r_n_97__47_;
      r_97__46_ <= r_n_97__46_;
      r_97__45_ <= r_n_97__45_;
      r_97__44_ <= r_n_97__44_;
      r_97__43_ <= r_n_97__43_;
      r_97__42_ <= r_n_97__42_;
      r_97__41_ <= r_n_97__41_;
      r_97__40_ <= r_n_97__40_;
      r_97__39_ <= r_n_97__39_;
      r_97__38_ <= r_n_97__38_;
      r_97__37_ <= r_n_97__37_;
      r_97__36_ <= r_n_97__36_;
      r_97__35_ <= r_n_97__35_;
      r_97__34_ <= r_n_97__34_;
      r_97__33_ <= r_n_97__33_;
      r_97__32_ <= r_n_97__32_;
      r_97__31_ <= r_n_97__31_;
      r_97__30_ <= r_n_97__30_;
      r_97__29_ <= r_n_97__29_;
      r_97__28_ <= r_n_97__28_;
      r_97__27_ <= r_n_97__27_;
      r_97__26_ <= r_n_97__26_;
      r_97__25_ <= r_n_97__25_;
      r_97__24_ <= r_n_97__24_;
      r_97__23_ <= r_n_97__23_;
      r_97__22_ <= r_n_97__22_;
      r_97__21_ <= r_n_97__21_;
      r_97__20_ <= r_n_97__20_;
      r_97__19_ <= r_n_97__19_;
      r_97__18_ <= r_n_97__18_;
      r_97__17_ <= r_n_97__17_;
      r_97__16_ <= r_n_97__16_;
      r_97__15_ <= r_n_97__15_;
      r_97__14_ <= r_n_97__14_;
      r_97__13_ <= r_n_97__13_;
      r_97__12_ <= r_n_97__12_;
      r_97__11_ <= r_n_97__11_;
      r_97__10_ <= r_n_97__10_;
      r_97__9_ <= r_n_97__9_;
      r_97__8_ <= r_n_97__8_;
      r_97__7_ <= r_n_97__7_;
      r_97__6_ <= r_n_97__6_;
      r_97__5_ <= r_n_97__5_;
      r_97__4_ <= r_n_97__4_;
      r_97__3_ <= r_n_97__3_;
      r_97__2_ <= r_n_97__2_;
      r_97__1_ <= r_n_97__1_;
      r_97__0_ <= r_n_97__0_;
    end 
    if(N3682) begin
      r_98__63_ <= r_n_98__63_;
      r_98__62_ <= r_n_98__62_;
      r_98__61_ <= r_n_98__61_;
      r_98__60_ <= r_n_98__60_;
      r_98__59_ <= r_n_98__59_;
      r_98__58_ <= r_n_98__58_;
      r_98__57_ <= r_n_98__57_;
      r_98__56_ <= r_n_98__56_;
      r_98__55_ <= r_n_98__55_;
      r_98__54_ <= r_n_98__54_;
      r_98__53_ <= r_n_98__53_;
      r_98__52_ <= r_n_98__52_;
      r_98__51_ <= r_n_98__51_;
      r_98__50_ <= r_n_98__50_;
      r_98__49_ <= r_n_98__49_;
      r_98__48_ <= r_n_98__48_;
      r_98__47_ <= r_n_98__47_;
      r_98__46_ <= r_n_98__46_;
      r_98__45_ <= r_n_98__45_;
      r_98__44_ <= r_n_98__44_;
      r_98__43_ <= r_n_98__43_;
      r_98__42_ <= r_n_98__42_;
      r_98__41_ <= r_n_98__41_;
      r_98__40_ <= r_n_98__40_;
      r_98__39_ <= r_n_98__39_;
      r_98__38_ <= r_n_98__38_;
      r_98__37_ <= r_n_98__37_;
      r_98__36_ <= r_n_98__36_;
      r_98__35_ <= r_n_98__35_;
      r_98__34_ <= r_n_98__34_;
      r_98__33_ <= r_n_98__33_;
      r_98__32_ <= r_n_98__32_;
      r_98__31_ <= r_n_98__31_;
      r_98__30_ <= r_n_98__30_;
      r_98__29_ <= r_n_98__29_;
      r_98__28_ <= r_n_98__28_;
      r_98__27_ <= r_n_98__27_;
      r_98__26_ <= r_n_98__26_;
      r_98__25_ <= r_n_98__25_;
      r_98__24_ <= r_n_98__24_;
      r_98__23_ <= r_n_98__23_;
      r_98__22_ <= r_n_98__22_;
      r_98__21_ <= r_n_98__21_;
      r_98__20_ <= r_n_98__20_;
      r_98__19_ <= r_n_98__19_;
      r_98__18_ <= r_n_98__18_;
      r_98__17_ <= r_n_98__17_;
      r_98__16_ <= r_n_98__16_;
      r_98__15_ <= r_n_98__15_;
      r_98__14_ <= r_n_98__14_;
      r_98__13_ <= r_n_98__13_;
      r_98__12_ <= r_n_98__12_;
      r_98__11_ <= r_n_98__11_;
      r_98__10_ <= r_n_98__10_;
      r_98__9_ <= r_n_98__9_;
      r_98__8_ <= r_n_98__8_;
      r_98__7_ <= r_n_98__7_;
      r_98__6_ <= r_n_98__6_;
      r_98__5_ <= r_n_98__5_;
      r_98__4_ <= r_n_98__4_;
      r_98__3_ <= r_n_98__3_;
      r_98__2_ <= r_n_98__2_;
      r_98__1_ <= r_n_98__1_;
      r_98__0_ <= r_n_98__0_;
    end 
    if(N3683) begin
      r_99__63_ <= r_n_99__63_;
      r_99__62_ <= r_n_99__62_;
      r_99__61_ <= r_n_99__61_;
      r_99__60_ <= r_n_99__60_;
      r_99__59_ <= r_n_99__59_;
      r_99__58_ <= r_n_99__58_;
      r_99__57_ <= r_n_99__57_;
      r_99__56_ <= r_n_99__56_;
      r_99__55_ <= r_n_99__55_;
      r_99__54_ <= r_n_99__54_;
      r_99__53_ <= r_n_99__53_;
      r_99__52_ <= r_n_99__52_;
      r_99__51_ <= r_n_99__51_;
      r_99__50_ <= r_n_99__50_;
      r_99__49_ <= r_n_99__49_;
      r_99__48_ <= r_n_99__48_;
      r_99__47_ <= r_n_99__47_;
      r_99__46_ <= r_n_99__46_;
      r_99__45_ <= r_n_99__45_;
      r_99__44_ <= r_n_99__44_;
      r_99__43_ <= r_n_99__43_;
      r_99__42_ <= r_n_99__42_;
      r_99__41_ <= r_n_99__41_;
      r_99__40_ <= r_n_99__40_;
      r_99__39_ <= r_n_99__39_;
      r_99__38_ <= r_n_99__38_;
      r_99__37_ <= r_n_99__37_;
      r_99__36_ <= r_n_99__36_;
      r_99__35_ <= r_n_99__35_;
      r_99__34_ <= r_n_99__34_;
      r_99__33_ <= r_n_99__33_;
      r_99__32_ <= r_n_99__32_;
      r_99__31_ <= r_n_99__31_;
      r_99__30_ <= r_n_99__30_;
      r_99__29_ <= r_n_99__29_;
      r_99__28_ <= r_n_99__28_;
      r_99__27_ <= r_n_99__27_;
      r_99__26_ <= r_n_99__26_;
      r_99__25_ <= r_n_99__25_;
      r_99__24_ <= r_n_99__24_;
      r_99__23_ <= r_n_99__23_;
      r_99__22_ <= r_n_99__22_;
      r_99__21_ <= r_n_99__21_;
      r_99__20_ <= r_n_99__20_;
      r_99__19_ <= r_n_99__19_;
      r_99__18_ <= r_n_99__18_;
      r_99__17_ <= r_n_99__17_;
      r_99__16_ <= r_n_99__16_;
      r_99__15_ <= r_n_99__15_;
      r_99__14_ <= r_n_99__14_;
      r_99__13_ <= r_n_99__13_;
      r_99__12_ <= r_n_99__12_;
      r_99__11_ <= r_n_99__11_;
      r_99__10_ <= r_n_99__10_;
      r_99__9_ <= r_n_99__9_;
      r_99__8_ <= r_n_99__8_;
      r_99__7_ <= r_n_99__7_;
      r_99__6_ <= r_n_99__6_;
      r_99__5_ <= r_n_99__5_;
      r_99__4_ <= r_n_99__4_;
      r_99__3_ <= r_n_99__3_;
      r_99__2_ <= r_n_99__2_;
      r_99__1_ <= r_n_99__1_;
      r_99__0_ <= r_n_99__0_;
    end 
    if(N3684) begin
      r_100__63_ <= r_n_100__63_;
      r_100__62_ <= r_n_100__62_;
      r_100__61_ <= r_n_100__61_;
      r_100__60_ <= r_n_100__60_;
      r_100__59_ <= r_n_100__59_;
      r_100__58_ <= r_n_100__58_;
      r_100__57_ <= r_n_100__57_;
      r_100__56_ <= r_n_100__56_;
      r_100__55_ <= r_n_100__55_;
      r_100__54_ <= r_n_100__54_;
      r_100__53_ <= r_n_100__53_;
      r_100__52_ <= r_n_100__52_;
      r_100__51_ <= r_n_100__51_;
      r_100__50_ <= r_n_100__50_;
      r_100__49_ <= r_n_100__49_;
      r_100__48_ <= r_n_100__48_;
      r_100__47_ <= r_n_100__47_;
      r_100__46_ <= r_n_100__46_;
      r_100__45_ <= r_n_100__45_;
      r_100__44_ <= r_n_100__44_;
      r_100__43_ <= r_n_100__43_;
      r_100__42_ <= r_n_100__42_;
      r_100__41_ <= r_n_100__41_;
      r_100__40_ <= r_n_100__40_;
      r_100__39_ <= r_n_100__39_;
      r_100__38_ <= r_n_100__38_;
      r_100__37_ <= r_n_100__37_;
      r_100__36_ <= r_n_100__36_;
      r_100__35_ <= r_n_100__35_;
      r_100__34_ <= r_n_100__34_;
      r_100__33_ <= r_n_100__33_;
      r_100__32_ <= r_n_100__32_;
      r_100__31_ <= r_n_100__31_;
      r_100__30_ <= r_n_100__30_;
      r_100__29_ <= r_n_100__29_;
      r_100__28_ <= r_n_100__28_;
      r_100__27_ <= r_n_100__27_;
      r_100__26_ <= r_n_100__26_;
      r_100__25_ <= r_n_100__25_;
      r_100__24_ <= r_n_100__24_;
      r_100__23_ <= r_n_100__23_;
      r_100__22_ <= r_n_100__22_;
      r_100__21_ <= r_n_100__21_;
      r_100__20_ <= r_n_100__20_;
      r_100__19_ <= r_n_100__19_;
      r_100__18_ <= r_n_100__18_;
      r_100__17_ <= r_n_100__17_;
      r_100__16_ <= r_n_100__16_;
      r_100__15_ <= r_n_100__15_;
      r_100__14_ <= r_n_100__14_;
      r_100__13_ <= r_n_100__13_;
      r_100__12_ <= r_n_100__12_;
      r_100__11_ <= r_n_100__11_;
      r_100__10_ <= r_n_100__10_;
      r_100__9_ <= r_n_100__9_;
      r_100__8_ <= r_n_100__8_;
      r_100__7_ <= r_n_100__7_;
      r_100__6_ <= r_n_100__6_;
      r_100__5_ <= r_n_100__5_;
      r_100__4_ <= r_n_100__4_;
      r_100__3_ <= r_n_100__3_;
      r_100__2_ <= r_n_100__2_;
      r_100__1_ <= r_n_100__1_;
      r_100__0_ <= r_n_100__0_;
    end 
    if(N3685) begin
      r_101__63_ <= r_n_101__63_;
      r_101__62_ <= r_n_101__62_;
      r_101__61_ <= r_n_101__61_;
      r_101__60_ <= r_n_101__60_;
      r_101__59_ <= r_n_101__59_;
      r_101__58_ <= r_n_101__58_;
      r_101__57_ <= r_n_101__57_;
      r_101__56_ <= r_n_101__56_;
      r_101__55_ <= r_n_101__55_;
      r_101__54_ <= r_n_101__54_;
      r_101__53_ <= r_n_101__53_;
      r_101__52_ <= r_n_101__52_;
      r_101__51_ <= r_n_101__51_;
      r_101__50_ <= r_n_101__50_;
      r_101__49_ <= r_n_101__49_;
      r_101__48_ <= r_n_101__48_;
      r_101__47_ <= r_n_101__47_;
      r_101__46_ <= r_n_101__46_;
      r_101__45_ <= r_n_101__45_;
      r_101__44_ <= r_n_101__44_;
      r_101__43_ <= r_n_101__43_;
      r_101__42_ <= r_n_101__42_;
      r_101__41_ <= r_n_101__41_;
      r_101__40_ <= r_n_101__40_;
      r_101__39_ <= r_n_101__39_;
      r_101__38_ <= r_n_101__38_;
      r_101__37_ <= r_n_101__37_;
      r_101__36_ <= r_n_101__36_;
      r_101__35_ <= r_n_101__35_;
      r_101__34_ <= r_n_101__34_;
      r_101__33_ <= r_n_101__33_;
      r_101__32_ <= r_n_101__32_;
      r_101__31_ <= r_n_101__31_;
      r_101__30_ <= r_n_101__30_;
      r_101__29_ <= r_n_101__29_;
      r_101__28_ <= r_n_101__28_;
      r_101__27_ <= r_n_101__27_;
      r_101__26_ <= r_n_101__26_;
      r_101__25_ <= r_n_101__25_;
      r_101__24_ <= r_n_101__24_;
      r_101__23_ <= r_n_101__23_;
      r_101__22_ <= r_n_101__22_;
      r_101__21_ <= r_n_101__21_;
      r_101__20_ <= r_n_101__20_;
      r_101__19_ <= r_n_101__19_;
      r_101__18_ <= r_n_101__18_;
      r_101__17_ <= r_n_101__17_;
      r_101__16_ <= r_n_101__16_;
      r_101__15_ <= r_n_101__15_;
      r_101__14_ <= r_n_101__14_;
      r_101__13_ <= r_n_101__13_;
      r_101__12_ <= r_n_101__12_;
      r_101__11_ <= r_n_101__11_;
      r_101__10_ <= r_n_101__10_;
      r_101__9_ <= r_n_101__9_;
      r_101__8_ <= r_n_101__8_;
      r_101__7_ <= r_n_101__7_;
      r_101__6_ <= r_n_101__6_;
      r_101__5_ <= r_n_101__5_;
      r_101__4_ <= r_n_101__4_;
      r_101__3_ <= r_n_101__3_;
      r_101__2_ <= r_n_101__2_;
      r_101__1_ <= r_n_101__1_;
      r_101__0_ <= r_n_101__0_;
    end 
    if(N3686) begin
      r_102__63_ <= r_n_102__63_;
      r_102__62_ <= r_n_102__62_;
      r_102__61_ <= r_n_102__61_;
      r_102__60_ <= r_n_102__60_;
      r_102__59_ <= r_n_102__59_;
      r_102__58_ <= r_n_102__58_;
      r_102__57_ <= r_n_102__57_;
      r_102__56_ <= r_n_102__56_;
      r_102__55_ <= r_n_102__55_;
      r_102__54_ <= r_n_102__54_;
      r_102__53_ <= r_n_102__53_;
      r_102__52_ <= r_n_102__52_;
      r_102__51_ <= r_n_102__51_;
      r_102__50_ <= r_n_102__50_;
      r_102__49_ <= r_n_102__49_;
      r_102__48_ <= r_n_102__48_;
      r_102__47_ <= r_n_102__47_;
      r_102__46_ <= r_n_102__46_;
      r_102__45_ <= r_n_102__45_;
      r_102__44_ <= r_n_102__44_;
      r_102__43_ <= r_n_102__43_;
      r_102__42_ <= r_n_102__42_;
      r_102__41_ <= r_n_102__41_;
      r_102__40_ <= r_n_102__40_;
      r_102__39_ <= r_n_102__39_;
      r_102__38_ <= r_n_102__38_;
      r_102__37_ <= r_n_102__37_;
      r_102__36_ <= r_n_102__36_;
      r_102__35_ <= r_n_102__35_;
      r_102__34_ <= r_n_102__34_;
      r_102__33_ <= r_n_102__33_;
      r_102__32_ <= r_n_102__32_;
      r_102__31_ <= r_n_102__31_;
      r_102__30_ <= r_n_102__30_;
      r_102__29_ <= r_n_102__29_;
      r_102__28_ <= r_n_102__28_;
      r_102__27_ <= r_n_102__27_;
      r_102__26_ <= r_n_102__26_;
      r_102__25_ <= r_n_102__25_;
      r_102__24_ <= r_n_102__24_;
      r_102__23_ <= r_n_102__23_;
      r_102__22_ <= r_n_102__22_;
      r_102__21_ <= r_n_102__21_;
      r_102__20_ <= r_n_102__20_;
      r_102__19_ <= r_n_102__19_;
      r_102__18_ <= r_n_102__18_;
      r_102__17_ <= r_n_102__17_;
      r_102__16_ <= r_n_102__16_;
      r_102__15_ <= r_n_102__15_;
      r_102__14_ <= r_n_102__14_;
      r_102__13_ <= r_n_102__13_;
      r_102__12_ <= r_n_102__12_;
      r_102__11_ <= r_n_102__11_;
      r_102__10_ <= r_n_102__10_;
      r_102__9_ <= r_n_102__9_;
      r_102__8_ <= r_n_102__8_;
      r_102__7_ <= r_n_102__7_;
      r_102__6_ <= r_n_102__6_;
      r_102__5_ <= r_n_102__5_;
      r_102__4_ <= r_n_102__4_;
      r_102__3_ <= r_n_102__3_;
      r_102__2_ <= r_n_102__2_;
      r_102__1_ <= r_n_102__1_;
      r_102__0_ <= r_n_102__0_;
    end 
    if(N3687) begin
      r_103__63_ <= r_n_103__63_;
      r_103__62_ <= r_n_103__62_;
      r_103__61_ <= r_n_103__61_;
      r_103__60_ <= r_n_103__60_;
      r_103__59_ <= r_n_103__59_;
      r_103__58_ <= r_n_103__58_;
      r_103__57_ <= r_n_103__57_;
      r_103__56_ <= r_n_103__56_;
      r_103__55_ <= r_n_103__55_;
      r_103__54_ <= r_n_103__54_;
      r_103__53_ <= r_n_103__53_;
      r_103__52_ <= r_n_103__52_;
      r_103__51_ <= r_n_103__51_;
      r_103__50_ <= r_n_103__50_;
      r_103__49_ <= r_n_103__49_;
      r_103__48_ <= r_n_103__48_;
      r_103__47_ <= r_n_103__47_;
      r_103__46_ <= r_n_103__46_;
      r_103__45_ <= r_n_103__45_;
      r_103__44_ <= r_n_103__44_;
      r_103__43_ <= r_n_103__43_;
      r_103__42_ <= r_n_103__42_;
      r_103__41_ <= r_n_103__41_;
      r_103__40_ <= r_n_103__40_;
      r_103__39_ <= r_n_103__39_;
      r_103__38_ <= r_n_103__38_;
      r_103__37_ <= r_n_103__37_;
      r_103__36_ <= r_n_103__36_;
      r_103__35_ <= r_n_103__35_;
      r_103__34_ <= r_n_103__34_;
      r_103__33_ <= r_n_103__33_;
      r_103__32_ <= r_n_103__32_;
      r_103__31_ <= r_n_103__31_;
      r_103__30_ <= r_n_103__30_;
      r_103__29_ <= r_n_103__29_;
      r_103__28_ <= r_n_103__28_;
      r_103__27_ <= r_n_103__27_;
      r_103__26_ <= r_n_103__26_;
      r_103__25_ <= r_n_103__25_;
      r_103__24_ <= r_n_103__24_;
      r_103__23_ <= r_n_103__23_;
      r_103__22_ <= r_n_103__22_;
      r_103__21_ <= r_n_103__21_;
      r_103__20_ <= r_n_103__20_;
      r_103__19_ <= r_n_103__19_;
      r_103__18_ <= r_n_103__18_;
      r_103__17_ <= r_n_103__17_;
      r_103__16_ <= r_n_103__16_;
      r_103__15_ <= r_n_103__15_;
      r_103__14_ <= r_n_103__14_;
      r_103__13_ <= r_n_103__13_;
      r_103__12_ <= r_n_103__12_;
      r_103__11_ <= r_n_103__11_;
      r_103__10_ <= r_n_103__10_;
      r_103__9_ <= r_n_103__9_;
      r_103__8_ <= r_n_103__8_;
      r_103__7_ <= r_n_103__7_;
      r_103__6_ <= r_n_103__6_;
      r_103__5_ <= r_n_103__5_;
      r_103__4_ <= r_n_103__4_;
      r_103__3_ <= r_n_103__3_;
      r_103__2_ <= r_n_103__2_;
      r_103__1_ <= r_n_103__1_;
      r_103__0_ <= r_n_103__0_;
    end 
    if(N3688) begin
      r_104__63_ <= r_n_104__63_;
      r_104__62_ <= r_n_104__62_;
      r_104__61_ <= r_n_104__61_;
      r_104__60_ <= r_n_104__60_;
      r_104__59_ <= r_n_104__59_;
      r_104__58_ <= r_n_104__58_;
      r_104__57_ <= r_n_104__57_;
      r_104__56_ <= r_n_104__56_;
      r_104__55_ <= r_n_104__55_;
      r_104__54_ <= r_n_104__54_;
      r_104__53_ <= r_n_104__53_;
      r_104__52_ <= r_n_104__52_;
      r_104__51_ <= r_n_104__51_;
      r_104__50_ <= r_n_104__50_;
      r_104__49_ <= r_n_104__49_;
      r_104__48_ <= r_n_104__48_;
      r_104__47_ <= r_n_104__47_;
      r_104__46_ <= r_n_104__46_;
      r_104__45_ <= r_n_104__45_;
      r_104__44_ <= r_n_104__44_;
      r_104__43_ <= r_n_104__43_;
      r_104__42_ <= r_n_104__42_;
      r_104__41_ <= r_n_104__41_;
      r_104__40_ <= r_n_104__40_;
      r_104__39_ <= r_n_104__39_;
      r_104__38_ <= r_n_104__38_;
      r_104__37_ <= r_n_104__37_;
      r_104__36_ <= r_n_104__36_;
      r_104__35_ <= r_n_104__35_;
      r_104__34_ <= r_n_104__34_;
      r_104__33_ <= r_n_104__33_;
      r_104__32_ <= r_n_104__32_;
      r_104__31_ <= r_n_104__31_;
      r_104__30_ <= r_n_104__30_;
      r_104__29_ <= r_n_104__29_;
      r_104__28_ <= r_n_104__28_;
      r_104__27_ <= r_n_104__27_;
      r_104__26_ <= r_n_104__26_;
      r_104__25_ <= r_n_104__25_;
      r_104__24_ <= r_n_104__24_;
      r_104__23_ <= r_n_104__23_;
      r_104__22_ <= r_n_104__22_;
      r_104__21_ <= r_n_104__21_;
      r_104__20_ <= r_n_104__20_;
      r_104__19_ <= r_n_104__19_;
      r_104__18_ <= r_n_104__18_;
      r_104__17_ <= r_n_104__17_;
      r_104__16_ <= r_n_104__16_;
      r_104__15_ <= r_n_104__15_;
      r_104__14_ <= r_n_104__14_;
      r_104__13_ <= r_n_104__13_;
      r_104__12_ <= r_n_104__12_;
      r_104__11_ <= r_n_104__11_;
      r_104__10_ <= r_n_104__10_;
      r_104__9_ <= r_n_104__9_;
      r_104__8_ <= r_n_104__8_;
      r_104__7_ <= r_n_104__7_;
      r_104__6_ <= r_n_104__6_;
      r_104__5_ <= r_n_104__5_;
      r_104__4_ <= r_n_104__4_;
      r_104__3_ <= r_n_104__3_;
      r_104__2_ <= r_n_104__2_;
      r_104__1_ <= r_n_104__1_;
      r_104__0_ <= r_n_104__0_;
    end 
    if(N3689) begin
      r_105__63_ <= r_n_105__63_;
      r_105__62_ <= r_n_105__62_;
      r_105__61_ <= r_n_105__61_;
      r_105__60_ <= r_n_105__60_;
      r_105__59_ <= r_n_105__59_;
      r_105__58_ <= r_n_105__58_;
      r_105__57_ <= r_n_105__57_;
      r_105__56_ <= r_n_105__56_;
      r_105__55_ <= r_n_105__55_;
      r_105__54_ <= r_n_105__54_;
      r_105__53_ <= r_n_105__53_;
      r_105__52_ <= r_n_105__52_;
      r_105__51_ <= r_n_105__51_;
      r_105__50_ <= r_n_105__50_;
      r_105__49_ <= r_n_105__49_;
      r_105__48_ <= r_n_105__48_;
      r_105__47_ <= r_n_105__47_;
      r_105__46_ <= r_n_105__46_;
      r_105__45_ <= r_n_105__45_;
      r_105__44_ <= r_n_105__44_;
      r_105__43_ <= r_n_105__43_;
      r_105__42_ <= r_n_105__42_;
      r_105__41_ <= r_n_105__41_;
      r_105__40_ <= r_n_105__40_;
      r_105__39_ <= r_n_105__39_;
      r_105__38_ <= r_n_105__38_;
      r_105__37_ <= r_n_105__37_;
      r_105__36_ <= r_n_105__36_;
      r_105__35_ <= r_n_105__35_;
      r_105__34_ <= r_n_105__34_;
      r_105__33_ <= r_n_105__33_;
      r_105__32_ <= r_n_105__32_;
      r_105__31_ <= r_n_105__31_;
      r_105__30_ <= r_n_105__30_;
      r_105__29_ <= r_n_105__29_;
      r_105__28_ <= r_n_105__28_;
      r_105__27_ <= r_n_105__27_;
      r_105__26_ <= r_n_105__26_;
      r_105__25_ <= r_n_105__25_;
      r_105__24_ <= r_n_105__24_;
      r_105__23_ <= r_n_105__23_;
      r_105__22_ <= r_n_105__22_;
      r_105__21_ <= r_n_105__21_;
      r_105__20_ <= r_n_105__20_;
      r_105__19_ <= r_n_105__19_;
      r_105__18_ <= r_n_105__18_;
      r_105__17_ <= r_n_105__17_;
      r_105__16_ <= r_n_105__16_;
      r_105__15_ <= r_n_105__15_;
      r_105__14_ <= r_n_105__14_;
      r_105__13_ <= r_n_105__13_;
      r_105__12_ <= r_n_105__12_;
      r_105__11_ <= r_n_105__11_;
      r_105__10_ <= r_n_105__10_;
      r_105__9_ <= r_n_105__9_;
      r_105__8_ <= r_n_105__8_;
      r_105__7_ <= r_n_105__7_;
      r_105__6_ <= r_n_105__6_;
      r_105__5_ <= r_n_105__5_;
      r_105__4_ <= r_n_105__4_;
      r_105__3_ <= r_n_105__3_;
      r_105__2_ <= r_n_105__2_;
      r_105__1_ <= r_n_105__1_;
      r_105__0_ <= r_n_105__0_;
    end 
    if(N3690) begin
      r_106__63_ <= r_n_106__63_;
      r_106__62_ <= r_n_106__62_;
      r_106__61_ <= r_n_106__61_;
      r_106__60_ <= r_n_106__60_;
      r_106__59_ <= r_n_106__59_;
      r_106__58_ <= r_n_106__58_;
      r_106__57_ <= r_n_106__57_;
      r_106__56_ <= r_n_106__56_;
      r_106__55_ <= r_n_106__55_;
      r_106__54_ <= r_n_106__54_;
      r_106__53_ <= r_n_106__53_;
      r_106__52_ <= r_n_106__52_;
      r_106__51_ <= r_n_106__51_;
      r_106__50_ <= r_n_106__50_;
      r_106__49_ <= r_n_106__49_;
      r_106__48_ <= r_n_106__48_;
      r_106__47_ <= r_n_106__47_;
      r_106__46_ <= r_n_106__46_;
      r_106__45_ <= r_n_106__45_;
      r_106__44_ <= r_n_106__44_;
      r_106__43_ <= r_n_106__43_;
      r_106__42_ <= r_n_106__42_;
      r_106__41_ <= r_n_106__41_;
      r_106__40_ <= r_n_106__40_;
      r_106__39_ <= r_n_106__39_;
      r_106__38_ <= r_n_106__38_;
      r_106__37_ <= r_n_106__37_;
      r_106__36_ <= r_n_106__36_;
      r_106__35_ <= r_n_106__35_;
      r_106__34_ <= r_n_106__34_;
      r_106__33_ <= r_n_106__33_;
      r_106__32_ <= r_n_106__32_;
      r_106__31_ <= r_n_106__31_;
      r_106__30_ <= r_n_106__30_;
      r_106__29_ <= r_n_106__29_;
      r_106__28_ <= r_n_106__28_;
      r_106__27_ <= r_n_106__27_;
      r_106__26_ <= r_n_106__26_;
      r_106__25_ <= r_n_106__25_;
      r_106__24_ <= r_n_106__24_;
      r_106__23_ <= r_n_106__23_;
      r_106__22_ <= r_n_106__22_;
      r_106__21_ <= r_n_106__21_;
      r_106__20_ <= r_n_106__20_;
      r_106__19_ <= r_n_106__19_;
      r_106__18_ <= r_n_106__18_;
      r_106__17_ <= r_n_106__17_;
      r_106__16_ <= r_n_106__16_;
      r_106__15_ <= r_n_106__15_;
      r_106__14_ <= r_n_106__14_;
      r_106__13_ <= r_n_106__13_;
      r_106__12_ <= r_n_106__12_;
      r_106__11_ <= r_n_106__11_;
      r_106__10_ <= r_n_106__10_;
      r_106__9_ <= r_n_106__9_;
      r_106__8_ <= r_n_106__8_;
      r_106__7_ <= r_n_106__7_;
      r_106__6_ <= r_n_106__6_;
      r_106__5_ <= r_n_106__5_;
      r_106__4_ <= r_n_106__4_;
      r_106__3_ <= r_n_106__3_;
      r_106__2_ <= r_n_106__2_;
      r_106__1_ <= r_n_106__1_;
      r_106__0_ <= r_n_106__0_;
    end 
    if(N3691) begin
      r_107__63_ <= r_n_107__63_;
      r_107__62_ <= r_n_107__62_;
      r_107__61_ <= r_n_107__61_;
      r_107__60_ <= r_n_107__60_;
      r_107__59_ <= r_n_107__59_;
      r_107__58_ <= r_n_107__58_;
      r_107__57_ <= r_n_107__57_;
      r_107__56_ <= r_n_107__56_;
      r_107__55_ <= r_n_107__55_;
      r_107__54_ <= r_n_107__54_;
      r_107__53_ <= r_n_107__53_;
      r_107__52_ <= r_n_107__52_;
      r_107__51_ <= r_n_107__51_;
      r_107__50_ <= r_n_107__50_;
      r_107__49_ <= r_n_107__49_;
      r_107__48_ <= r_n_107__48_;
      r_107__47_ <= r_n_107__47_;
      r_107__46_ <= r_n_107__46_;
      r_107__45_ <= r_n_107__45_;
      r_107__44_ <= r_n_107__44_;
      r_107__43_ <= r_n_107__43_;
      r_107__42_ <= r_n_107__42_;
      r_107__41_ <= r_n_107__41_;
      r_107__40_ <= r_n_107__40_;
      r_107__39_ <= r_n_107__39_;
      r_107__38_ <= r_n_107__38_;
      r_107__37_ <= r_n_107__37_;
      r_107__36_ <= r_n_107__36_;
      r_107__35_ <= r_n_107__35_;
      r_107__34_ <= r_n_107__34_;
      r_107__33_ <= r_n_107__33_;
      r_107__32_ <= r_n_107__32_;
      r_107__31_ <= r_n_107__31_;
      r_107__30_ <= r_n_107__30_;
      r_107__29_ <= r_n_107__29_;
      r_107__28_ <= r_n_107__28_;
      r_107__27_ <= r_n_107__27_;
      r_107__26_ <= r_n_107__26_;
      r_107__25_ <= r_n_107__25_;
      r_107__24_ <= r_n_107__24_;
      r_107__23_ <= r_n_107__23_;
      r_107__22_ <= r_n_107__22_;
      r_107__21_ <= r_n_107__21_;
      r_107__20_ <= r_n_107__20_;
      r_107__19_ <= r_n_107__19_;
      r_107__18_ <= r_n_107__18_;
      r_107__17_ <= r_n_107__17_;
      r_107__16_ <= r_n_107__16_;
      r_107__15_ <= r_n_107__15_;
      r_107__14_ <= r_n_107__14_;
      r_107__13_ <= r_n_107__13_;
      r_107__12_ <= r_n_107__12_;
      r_107__11_ <= r_n_107__11_;
      r_107__10_ <= r_n_107__10_;
      r_107__9_ <= r_n_107__9_;
      r_107__8_ <= r_n_107__8_;
      r_107__7_ <= r_n_107__7_;
      r_107__6_ <= r_n_107__6_;
      r_107__5_ <= r_n_107__5_;
      r_107__4_ <= r_n_107__4_;
      r_107__3_ <= r_n_107__3_;
      r_107__2_ <= r_n_107__2_;
      r_107__1_ <= r_n_107__1_;
      r_107__0_ <= r_n_107__0_;
    end 
    if(N3692) begin
      r_108__63_ <= r_n_108__63_;
      r_108__62_ <= r_n_108__62_;
      r_108__61_ <= r_n_108__61_;
      r_108__60_ <= r_n_108__60_;
      r_108__59_ <= r_n_108__59_;
      r_108__58_ <= r_n_108__58_;
      r_108__57_ <= r_n_108__57_;
      r_108__56_ <= r_n_108__56_;
      r_108__55_ <= r_n_108__55_;
      r_108__54_ <= r_n_108__54_;
      r_108__53_ <= r_n_108__53_;
      r_108__52_ <= r_n_108__52_;
      r_108__51_ <= r_n_108__51_;
      r_108__50_ <= r_n_108__50_;
      r_108__49_ <= r_n_108__49_;
      r_108__48_ <= r_n_108__48_;
      r_108__47_ <= r_n_108__47_;
      r_108__46_ <= r_n_108__46_;
      r_108__45_ <= r_n_108__45_;
      r_108__44_ <= r_n_108__44_;
      r_108__43_ <= r_n_108__43_;
      r_108__42_ <= r_n_108__42_;
      r_108__41_ <= r_n_108__41_;
      r_108__40_ <= r_n_108__40_;
      r_108__39_ <= r_n_108__39_;
      r_108__38_ <= r_n_108__38_;
      r_108__37_ <= r_n_108__37_;
      r_108__36_ <= r_n_108__36_;
      r_108__35_ <= r_n_108__35_;
      r_108__34_ <= r_n_108__34_;
      r_108__33_ <= r_n_108__33_;
      r_108__32_ <= r_n_108__32_;
      r_108__31_ <= r_n_108__31_;
      r_108__30_ <= r_n_108__30_;
      r_108__29_ <= r_n_108__29_;
      r_108__28_ <= r_n_108__28_;
      r_108__27_ <= r_n_108__27_;
      r_108__26_ <= r_n_108__26_;
      r_108__25_ <= r_n_108__25_;
      r_108__24_ <= r_n_108__24_;
      r_108__23_ <= r_n_108__23_;
      r_108__22_ <= r_n_108__22_;
      r_108__21_ <= r_n_108__21_;
      r_108__20_ <= r_n_108__20_;
      r_108__19_ <= r_n_108__19_;
      r_108__18_ <= r_n_108__18_;
      r_108__17_ <= r_n_108__17_;
      r_108__16_ <= r_n_108__16_;
      r_108__15_ <= r_n_108__15_;
      r_108__14_ <= r_n_108__14_;
      r_108__13_ <= r_n_108__13_;
      r_108__12_ <= r_n_108__12_;
      r_108__11_ <= r_n_108__11_;
      r_108__10_ <= r_n_108__10_;
      r_108__9_ <= r_n_108__9_;
      r_108__8_ <= r_n_108__8_;
      r_108__7_ <= r_n_108__7_;
      r_108__6_ <= r_n_108__6_;
      r_108__5_ <= r_n_108__5_;
      r_108__4_ <= r_n_108__4_;
      r_108__3_ <= r_n_108__3_;
      r_108__2_ <= r_n_108__2_;
      r_108__1_ <= r_n_108__1_;
      r_108__0_ <= r_n_108__0_;
    end 
    if(N3693) begin
      r_109__63_ <= r_n_109__63_;
      r_109__62_ <= r_n_109__62_;
      r_109__61_ <= r_n_109__61_;
      r_109__60_ <= r_n_109__60_;
      r_109__59_ <= r_n_109__59_;
      r_109__58_ <= r_n_109__58_;
      r_109__57_ <= r_n_109__57_;
      r_109__56_ <= r_n_109__56_;
      r_109__55_ <= r_n_109__55_;
      r_109__54_ <= r_n_109__54_;
      r_109__53_ <= r_n_109__53_;
      r_109__52_ <= r_n_109__52_;
      r_109__51_ <= r_n_109__51_;
      r_109__50_ <= r_n_109__50_;
      r_109__49_ <= r_n_109__49_;
      r_109__48_ <= r_n_109__48_;
      r_109__47_ <= r_n_109__47_;
      r_109__46_ <= r_n_109__46_;
      r_109__45_ <= r_n_109__45_;
      r_109__44_ <= r_n_109__44_;
      r_109__43_ <= r_n_109__43_;
      r_109__42_ <= r_n_109__42_;
      r_109__41_ <= r_n_109__41_;
      r_109__40_ <= r_n_109__40_;
      r_109__39_ <= r_n_109__39_;
      r_109__38_ <= r_n_109__38_;
      r_109__37_ <= r_n_109__37_;
      r_109__36_ <= r_n_109__36_;
      r_109__35_ <= r_n_109__35_;
      r_109__34_ <= r_n_109__34_;
      r_109__33_ <= r_n_109__33_;
      r_109__32_ <= r_n_109__32_;
      r_109__31_ <= r_n_109__31_;
      r_109__30_ <= r_n_109__30_;
      r_109__29_ <= r_n_109__29_;
      r_109__28_ <= r_n_109__28_;
      r_109__27_ <= r_n_109__27_;
      r_109__26_ <= r_n_109__26_;
      r_109__25_ <= r_n_109__25_;
      r_109__24_ <= r_n_109__24_;
      r_109__23_ <= r_n_109__23_;
      r_109__22_ <= r_n_109__22_;
      r_109__21_ <= r_n_109__21_;
      r_109__20_ <= r_n_109__20_;
      r_109__19_ <= r_n_109__19_;
      r_109__18_ <= r_n_109__18_;
      r_109__17_ <= r_n_109__17_;
      r_109__16_ <= r_n_109__16_;
      r_109__15_ <= r_n_109__15_;
      r_109__14_ <= r_n_109__14_;
      r_109__13_ <= r_n_109__13_;
      r_109__12_ <= r_n_109__12_;
      r_109__11_ <= r_n_109__11_;
      r_109__10_ <= r_n_109__10_;
      r_109__9_ <= r_n_109__9_;
      r_109__8_ <= r_n_109__8_;
      r_109__7_ <= r_n_109__7_;
      r_109__6_ <= r_n_109__6_;
      r_109__5_ <= r_n_109__5_;
      r_109__4_ <= r_n_109__4_;
      r_109__3_ <= r_n_109__3_;
      r_109__2_ <= r_n_109__2_;
      r_109__1_ <= r_n_109__1_;
      r_109__0_ <= r_n_109__0_;
    end 
    if(N3694) begin
      r_110__63_ <= r_n_110__63_;
      r_110__62_ <= r_n_110__62_;
      r_110__61_ <= r_n_110__61_;
      r_110__60_ <= r_n_110__60_;
      r_110__59_ <= r_n_110__59_;
      r_110__58_ <= r_n_110__58_;
      r_110__57_ <= r_n_110__57_;
      r_110__56_ <= r_n_110__56_;
      r_110__55_ <= r_n_110__55_;
      r_110__54_ <= r_n_110__54_;
      r_110__53_ <= r_n_110__53_;
      r_110__52_ <= r_n_110__52_;
      r_110__51_ <= r_n_110__51_;
      r_110__50_ <= r_n_110__50_;
      r_110__49_ <= r_n_110__49_;
      r_110__48_ <= r_n_110__48_;
      r_110__47_ <= r_n_110__47_;
      r_110__46_ <= r_n_110__46_;
      r_110__45_ <= r_n_110__45_;
      r_110__44_ <= r_n_110__44_;
      r_110__43_ <= r_n_110__43_;
      r_110__42_ <= r_n_110__42_;
      r_110__41_ <= r_n_110__41_;
      r_110__40_ <= r_n_110__40_;
      r_110__39_ <= r_n_110__39_;
      r_110__38_ <= r_n_110__38_;
      r_110__37_ <= r_n_110__37_;
      r_110__36_ <= r_n_110__36_;
      r_110__35_ <= r_n_110__35_;
      r_110__34_ <= r_n_110__34_;
      r_110__33_ <= r_n_110__33_;
      r_110__32_ <= r_n_110__32_;
      r_110__31_ <= r_n_110__31_;
      r_110__30_ <= r_n_110__30_;
      r_110__29_ <= r_n_110__29_;
      r_110__28_ <= r_n_110__28_;
      r_110__27_ <= r_n_110__27_;
      r_110__26_ <= r_n_110__26_;
      r_110__25_ <= r_n_110__25_;
      r_110__24_ <= r_n_110__24_;
      r_110__23_ <= r_n_110__23_;
      r_110__22_ <= r_n_110__22_;
      r_110__21_ <= r_n_110__21_;
      r_110__20_ <= r_n_110__20_;
      r_110__19_ <= r_n_110__19_;
      r_110__18_ <= r_n_110__18_;
      r_110__17_ <= r_n_110__17_;
      r_110__16_ <= r_n_110__16_;
      r_110__15_ <= r_n_110__15_;
      r_110__14_ <= r_n_110__14_;
      r_110__13_ <= r_n_110__13_;
      r_110__12_ <= r_n_110__12_;
      r_110__11_ <= r_n_110__11_;
      r_110__10_ <= r_n_110__10_;
      r_110__9_ <= r_n_110__9_;
      r_110__8_ <= r_n_110__8_;
      r_110__7_ <= r_n_110__7_;
      r_110__6_ <= r_n_110__6_;
      r_110__5_ <= r_n_110__5_;
      r_110__4_ <= r_n_110__4_;
      r_110__3_ <= r_n_110__3_;
      r_110__2_ <= r_n_110__2_;
      r_110__1_ <= r_n_110__1_;
      r_110__0_ <= r_n_110__0_;
    end 
    if(N3695) begin
      r_111__63_ <= r_n_111__63_;
      r_111__62_ <= r_n_111__62_;
      r_111__61_ <= r_n_111__61_;
      r_111__60_ <= r_n_111__60_;
      r_111__59_ <= r_n_111__59_;
      r_111__58_ <= r_n_111__58_;
      r_111__57_ <= r_n_111__57_;
      r_111__56_ <= r_n_111__56_;
      r_111__55_ <= r_n_111__55_;
      r_111__54_ <= r_n_111__54_;
      r_111__53_ <= r_n_111__53_;
      r_111__52_ <= r_n_111__52_;
      r_111__51_ <= r_n_111__51_;
      r_111__50_ <= r_n_111__50_;
      r_111__49_ <= r_n_111__49_;
      r_111__48_ <= r_n_111__48_;
      r_111__47_ <= r_n_111__47_;
      r_111__46_ <= r_n_111__46_;
      r_111__45_ <= r_n_111__45_;
      r_111__44_ <= r_n_111__44_;
      r_111__43_ <= r_n_111__43_;
      r_111__42_ <= r_n_111__42_;
      r_111__41_ <= r_n_111__41_;
      r_111__40_ <= r_n_111__40_;
      r_111__39_ <= r_n_111__39_;
      r_111__38_ <= r_n_111__38_;
      r_111__37_ <= r_n_111__37_;
      r_111__36_ <= r_n_111__36_;
      r_111__35_ <= r_n_111__35_;
      r_111__34_ <= r_n_111__34_;
      r_111__33_ <= r_n_111__33_;
      r_111__32_ <= r_n_111__32_;
      r_111__31_ <= r_n_111__31_;
      r_111__30_ <= r_n_111__30_;
      r_111__29_ <= r_n_111__29_;
      r_111__28_ <= r_n_111__28_;
      r_111__27_ <= r_n_111__27_;
      r_111__26_ <= r_n_111__26_;
      r_111__25_ <= r_n_111__25_;
      r_111__24_ <= r_n_111__24_;
      r_111__23_ <= r_n_111__23_;
      r_111__22_ <= r_n_111__22_;
      r_111__21_ <= r_n_111__21_;
      r_111__20_ <= r_n_111__20_;
      r_111__19_ <= r_n_111__19_;
      r_111__18_ <= r_n_111__18_;
      r_111__17_ <= r_n_111__17_;
      r_111__16_ <= r_n_111__16_;
      r_111__15_ <= r_n_111__15_;
      r_111__14_ <= r_n_111__14_;
      r_111__13_ <= r_n_111__13_;
      r_111__12_ <= r_n_111__12_;
      r_111__11_ <= r_n_111__11_;
      r_111__10_ <= r_n_111__10_;
      r_111__9_ <= r_n_111__9_;
      r_111__8_ <= r_n_111__8_;
      r_111__7_ <= r_n_111__7_;
      r_111__6_ <= r_n_111__6_;
      r_111__5_ <= r_n_111__5_;
      r_111__4_ <= r_n_111__4_;
      r_111__3_ <= r_n_111__3_;
      r_111__2_ <= r_n_111__2_;
      r_111__1_ <= r_n_111__1_;
      r_111__0_ <= r_n_111__0_;
    end 
    if(N3696) begin
      r_112__63_ <= r_n_112__63_;
      r_112__62_ <= r_n_112__62_;
      r_112__61_ <= r_n_112__61_;
      r_112__60_ <= r_n_112__60_;
      r_112__59_ <= r_n_112__59_;
      r_112__58_ <= r_n_112__58_;
      r_112__57_ <= r_n_112__57_;
      r_112__56_ <= r_n_112__56_;
      r_112__55_ <= r_n_112__55_;
      r_112__54_ <= r_n_112__54_;
      r_112__53_ <= r_n_112__53_;
      r_112__52_ <= r_n_112__52_;
      r_112__51_ <= r_n_112__51_;
      r_112__50_ <= r_n_112__50_;
      r_112__49_ <= r_n_112__49_;
      r_112__48_ <= r_n_112__48_;
      r_112__47_ <= r_n_112__47_;
      r_112__46_ <= r_n_112__46_;
      r_112__45_ <= r_n_112__45_;
      r_112__44_ <= r_n_112__44_;
      r_112__43_ <= r_n_112__43_;
      r_112__42_ <= r_n_112__42_;
      r_112__41_ <= r_n_112__41_;
      r_112__40_ <= r_n_112__40_;
      r_112__39_ <= r_n_112__39_;
      r_112__38_ <= r_n_112__38_;
      r_112__37_ <= r_n_112__37_;
      r_112__36_ <= r_n_112__36_;
      r_112__35_ <= r_n_112__35_;
      r_112__34_ <= r_n_112__34_;
      r_112__33_ <= r_n_112__33_;
      r_112__32_ <= r_n_112__32_;
      r_112__31_ <= r_n_112__31_;
      r_112__30_ <= r_n_112__30_;
      r_112__29_ <= r_n_112__29_;
      r_112__28_ <= r_n_112__28_;
      r_112__27_ <= r_n_112__27_;
      r_112__26_ <= r_n_112__26_;
      r_112__25_ <= r_n_112__25_;
      r_112__24_ <= r_n_112__24_;
      r_112__23_ <= r_n_112__23_;
      r_112__22_ <= r_n_112__22_;
      r_112__21_ <= r_n_112__21_;
      r_112__20_ <= r_n_112__20_;
      r_112__19_ <= r_n_112__19_;
      r_112__18_ <= r_n_112__18_;
      r_112__17_ <= r_n_112__17_;
      r_112__16_ <= r_n_112__16_;
      r_112__15_ <= r_n_112__15_;
      r_112__14_ <= r_n_112__14_;
      r_112__13_ <= r_n_112__13_;
      r_112__12_ <= r_n_112__12_;
      r_112__11_ <= r_n_112__11_;
      r_112__10_ <= r_n_112__10_;
      r_112__9_ <= r_n_112__9_;
      r_112__8_ <= r_n_112__8_;
      r_112__7_ <= r_n_112__7_;
      r_112__6_ <= r_n_112__6_;
      r_112__5_ <= r_n_112__5_;
      r_112__4_ <= r_n_112__4_;
      r_112__3_ <= r_n_112__3_;
      r_112__2_ <= r_n_112__2_;
      r_112__1_ <= r_n_112__1_;
      r_112__0_ <= r_n_112__0_;
    end 
    if(N3697) begin
      r_113__63_ <= r_n_113__63_;
      r_113__62_ <= r_n_113__62_;
      r_113__61_ <= r_n_113__61_;
      r_113__60_ <= r_n_113__60_;
      r_113__59_ <= r_n_113__59_;
      r_113__58_ <= r_n_113__58_;
      r_113__57_ <= r_n_113__57_;
      r_113__56_ <= r_n_113__56_;
      r_113__55_ <= r_n_113__55_;
      r_113__54_ <= r_n_113__54_;
      r_113__53_ <= r_n_113__53_;
      r_113__52_ <= r_n_113__52_;
      r_113__51_ <= r_n_113__51_;
      r_113__50_ <= r_n_113__50_;
      r_113__49_ <= r_n_113__49_;
      r_113__48_ <= r_n_113__48_;
      r_113__47_ <= r_n_113__47_;
      r_113__46_ <= r_n_113__46_;
      r_113__45_ <= r_n_113__45_;
      r_113__44_ <= r_n_113__44_;
      r_113__43_ <= r_n_113__43_;
      r_113__42_ <= r_n_113__42_;
      r_113__41_ <= r_n_113__41_;
      r_113__40_ <= r_n_113__40_;
      r_113__39_ <= r_n_113__39_;
      r_113__38_ <= r_n_113__38_;
      r_113__37_ <= r_n_113__37_;
      r_113__36_ <= r_n_113__36_;
      r_113__35_ <= r_n_113__35_;
      r_113__34_ <= r_n_113__34_;
      r_113__33_ <= r_n_113__33_;
      r_113__32_ <= r_n_113__32_;
      r_113__31_ <= r_n_113__31_;
      r_113__30_ <= r_n_113__30_;
      r_113__29_ <= r_n_113__29_;
      r_113__28_ <= r_n_113__28_;
      r_113__27_ <= r_n_113__27_;
      r_113__26_ <= r_n_113__26_;
      r_113__25_ <= r_n_113__25_;
      r_113__24_ <= r_n_113__24_;
      r_113__23_ <= r_n_113__23_;
      r_113__22_ <= r_n_113__22_;
      r_113__21_ <= r_n_113__21_;
      r_113__20_ <= r_n_113__20_;
      r_113__19_ <= r_n_113__19_;
      r_113__18_ <= r_n_113__18_;
      r_113__17_ <= r_n_113__17_;
      r_113__16_ <= r_n_113__16_;
      r_113__15_ <= r_n_113__15_;
      r_113__14_ <= r_n_113__14_;
      r_113__13_ <= r_n_113__13_;
      r_113__12_ <= r_n_113__12_;
      r_113__11_ <= r_n_113__11_;
      r_113__10_ <= r_n_113__10_;
      r_113__9_ <= r_n_113__9_;
      r_113__8_ <= r_n_113__8_;
      r_113__7_ <= r_n_113__7_;
      r_113__6_ <= r_n_113__6_;
      r_113__5_ <= r_n_113__5_;
      r_113__4_ <= r_n_113__4_;
      r_113__3_ <= r_n_113__3_;
      r_113__2_ <= r_n_113__2_;
      r_113__1_ <= r_n_113__1_;
      r_113__0_ <= r_n_113__0_;
    end 
    if(N3698) begin
      r_114__63_ <= r_n_114__63_;
      r_114__62_ <= r_n_114__62_;
      r_114__61_ <= r_n_114__61_;
      r_114__60_ <= r_n_114__60_;
      r_114__59_ <= r_n_114__59_;
      r_114__58_ <= r_n_114__58_;
      r_114__57_ <= r_n_114__57_;
      r_114__56_ <= r_n_114__56_;
      r_114__55_ <= r_n_114__55_;
      r_114__54_ <= r_n_114__54_;
      r_114__53_ <= r_n_114__53_;
      r_114__52_ <= r_n_114__52_;
      r_114__51_ <= r_n_114__51_;
      r_114__50_ <= r_n_114__50_;
      r_114__49_ <= r_n_114__49_;
      r_114__48_ <= r_n_114__48_;
      r_114__47_ <= r_n_114__47_;
      r_114__46_ <= r_n_114__46_;
      r_114__45_ <= r_n_114__45_;
      r_114__44_ <= r_n_114__44_;
      r_114__43_ <= r_n_114__43_;
      r_114__42_ <= r_n_114__42_;
      r_114__41_ <= r_n_114__41_;
      r_114__40_ <= r_n_114__40_;
      r_114__39_ <= r_n_114__39_;
      r_114__38_ <= r_n_114__38_;
      r_114__37_ <= r_n_114__37_;
      r_114__36_ <= r_n_114__36_;
      r_114__35_ <= r_n_114__35_;
      r_114__34_ <= r_n_114__34_;
      r_114__33_ <= r_n_114__33_;
      r_114__32_ <= r_n_114__32_;
      r_114__31_ <= r_n_114__31_;
      r_114__30_ <= r_n_114__30_;
      r_114__29_ <= r_n_114__29_;
      r_114__28_ <= r_n_114__28_;
      r_114__27_ <= r_n_114__27_;
      r_114__26_ <= r_n_114__26_;
      r_114__25_ <= r_n_114__25_;
      r_114__24_ <= r_n_114__24_;
      r_114__23_ <= r_n_114__23_;
      r_114__22_ <= r_n_114__22_;
      r_114__21_ <= r_n_114__21_;
      r_114__20_ <= r_n_114__20_;
      r_114__19_ <= r_n_114__19_;
      r_114__18_ <= r_n_114__18_;
      r_114__17_ <= r_n_114__17_;
      r_114__16_ <= r_n_114__16_;
      r_114__15_ <= r_n_114__15_;
      r_114__14_ <= r_n_114__14_;
      r_114__13_ <= r_n_114__13_;
      r_114__12_ <= r_n_114__12_;
      r_114__11_ <= r_n_114__11_;
      r_114__10_ <= r_n_114__10_;
      r_114__9_ <= r_n_114__9_;
      r_114__8_ <= r_n_114__8_;
      r_114__7_ <= r_n_114__7_;
      r_114__6_ <= r_n_114__6_;
      r_114__5_ <= r_n_114__5_;
      r_114__4_ <= r_n_114__4_;
      r_114__3_ <= r_n_114__3_;
      r_114__2_ <= r_n_114__2_;
      r_114__1_ <= r_n_114__1_;
      r_114__0_ <= r_n_114__0_;
    end 
    if(N3699) begin
      r_115__63_ <= r_n_115__63_;
      r_115__62_ <= r_n_115__62_;
      r_115__61_ <= r_n_115__61_;
      r_115__60_ <= r_n_115__60_;
      r_115__59_ <= r_n_115__59_;
      r_115__58_ <= r_n_115__58_;
      r_115__57_ <= r_n_115__57_;
      r_115__56_ <= r_n_115__56_;
      r_115__55_ <= r_n_115__55_;
      r_115__54_ <= r_n_115__54_;
      r_115__53_ <= r_n_115__53_;
      r_115__52_ <= r_n_115__52_;
      r_115__51_ <= r_n_115__51_;
      r_115__50_ <= r_n_115__50_;
      r_115__49_ <= r_n_115__49_;
      r_115__48_ <= r_n_115__48_;
      r_115__47_ <= r_n_115__47_;
      r_115__46_ <= r_n_115__46_;
      r_115__45_ <= r_n_115__45_;
      r_115__44_ <= r_n_115__44_;
      r_115__43_ <= r_n_115__43_;
      r_115__42_ <= r_n_115__42_;
      r_115__41_ <= r_n_115__41_;
      r_115__40_ <= r_n_115__40_;
      r_115__39_ <= r_n_115__39_;
      r_115__38_ <= r_n_115__38_;
      r_115__37_ <= r_n_115__37_;
      r_115__36_ <= r_n_115__36_;
      r_115__35_ <= r_n_115__35_;
      r_115__34_ <= r_n_115__34_;
      r_115__33_ <= r_n_115__33_;
      r_115__32_ <= r_n_115__32_;
      r_115__31_ <= r_n_115__31_;
      r_115__30_ <= r_n_115__30_;
      r_115__29_ <= r_n_115__29_;
      r_115__28_ <= r_n_115__28_;
      r_115__27_ <= r_n_115__27_;
      r_115__26_ <= r_n_115__26_;
      r_115__25_ <= r_n_115__25_;
      r_115__24_ <= r_n_115__24_;
      r_115__23_ <= r_n_115__23_;
      r_115__22_ <= r_n_115__22_;
      r_115__21_ <= r_n_115__21_;
      r_115__20_ <= r_n_115__20_;
      r_115__19_ <= r_n_115__19_;
      r_115__18_ <= r_n_115__18_;
      r_115__17_ <= r_n_115__17_;
      r_115__16_ <= r_n_115__16_;
      r_115__15_ <= r_n_115__15_;
      r_115__14_ <= r_n_115__14_;
      r_115__13_ <= r_n_115__13_;
      r_115__12_ <= r_n_115__12_;
      r_115__11_ <= r_n_115__11_;
      r_115__10_ <= r_n_115__10_;
      r_115__9_ <= r_n_115__9_;
      r_115__8_ <= r_n_115__8_;
      r_115__7_ <= r_n_115__7_;
      r_115__6_ <= r_n_115__6_;
      r_115__5_ <= r_n_115__5_;
      r_115__4_ <= r_n_115__4_;
      r_115__3_ <= r_n_115__3_;
      r_115__2_ <= r_n_115__2_;
      r_115__1_ <= r_n_115__1_;
      r_115__0_ <= r_n_115__0_;
    end 
    if(N3700) begin
      r_116__63_ <= r_n_116__63_;
      r_116__62_ <= r_n_116__62_;
      r_116__61_ <= r_n_116__61_;
      r_116__60_ <= r_n_116__60_;
      r_116__59_ <= r_n_116__59_;
      r_116__58_ <= r_n_116__58_;
      r_116__57_ <= r_n_116__57_;
      r_116__56_ <= r_n_116__56_;
      r_116__55_ <= r_n_116__55_;
      r_116__54_ <= r_n_116__54_;
      r_116__53_ <= r_n_116__53_;
      r_116__52_ <= r_n_116__52_;
      r_116__51_ <= r_n_116__51_;
      r_116__50_ <= r_n_116__50_;
      r_116__49_ <= r_n_116__49_;
      r_116__48_ <= r_n_116__48_;
      r_116__47_ <= r_n_116__47_;
      r_116__46_ <= r_n_116__46_;
      r_116__45_ <= r_n_116__45_;
      r_116__44_ <= r_n_116__44_;
      r_116__43_ <= r_n_116__43_;
      r_116__42_ <= r_n_116__42_;
      r_116__41_ <= r_n_116__41_;
      r_116__40_ <= r_n_116__40_;
      r_116__39_ <= r_n_116__39_;
      r_116__38_ <= r_n_116__38_;
      r_116__37_ <= r_n_116__37_;
      r_116__36_ <= r_n_116__36_;
      r_116__35_ <= r_n_116__35_;
      r_116__34_ <= r_n_116__34_;
      r_116__33_ <= r_n_116__33_;
      r_116__32_ <= r_n_116__32_;
      r_116__31_ <= r_n_116__31_;
      r_116__30_ <= r_n_116__30_;
      r_116__29_ <= r_n_116__29_;
      r_116__28_ <= r_n_116__28_;
      r_116__27_ <= r_n_116__27_;
      r_116__26_ <= r_n_116__26_;
      r_116__25_ <= r_n_116__25_;
      r_116__24_ <= r_n_116__24_;
      r_116__23_ <= r_n_116__23_;
      r_116__22_ <= r_n_116__22_;
      r_116__21_ <= r_n_116__21_;
      r_116__20_ <= r_n_116__20_;
      r_116__19_ <= r_n_116__19_;
      r_116__18_ <= r_n_116__18_;
      r_116__17_ <= r_n_116__17_;
      r_116__16_ <= r_n_116__16_;
      r_116__15_ <= r_n_116__15_;
      r_116__14_ <= r_n_116__14_;
      r_116__13_ <= r_n_116__13_;
      r_116__12_ <= r_n_116__12_;
      r_116__11_ <= r_n_116__11_;
      r_116__10_ <= r_n_116__10_;
      r_116__9_ <= r_n_116__9_;
      r_116__8_ <= r_n_116__8_;
      r_116__7_ <= r_n_116__7_;
      r_116__6_ <= r_n_116__6_;
      r_116__5_ <= r_n_116__5_;
      r_116__4_ <= r_n_116__4_;
      r_116__3_ <= r_n_116__3_;
      r_116__2_ <= r_n_116__2_;
      r_116__1_ <= r_n_116__1_;
      r_116__0_ <= r_n_116__0_;
    end 
    if(N3701) begin
      r_117__63_ <= r_n_117__63_;
      r_117__62_ <= r_n_117__62_;
      r_117__61_ <= r_n_117__61_;
      r_117__60_ <= r_n_117__60_;
      r_117__59_ <= r_n_117__59_;
      r_117__58_ <= r_n_117__58_;
      r_117__57_ <= r_n_117__57_;
      r_117__56_ <= r_n_117__56_;
      r_117__55_ <= r_n_117__55_;
      r_117__54_ <= r_n_117__54_;
      r_117__53_ <= r_n_117__53_;
      r_117__52_ <= r_n_117__52_;
      r_117__51_ <= r_n_117__51_;
      r_117__50_ <= r_n_117__50_;
      r_117__49_ <= r_n_117__49_;
      r_117__48_ <= r_n_117__48_;
      r_117__47_ <= r_n_117__47_;
      r_117__46_ <= r_n_117__46_;
      r_117__45_ <= r_n_117__45_;
      r_117__44_ <= r_n_117__44_;
      r_117__43_ <= r_n_117__43_;
      r_117__42_ <= r_n_117__42_;
      r_117__41_ <= r_n_117__41_;
      r_117__40_ <= r_n_117__40_;
      r_117__39_ <= r_n_117__39_;
      r_117__38_ <= r_n_117__38_;
      r_117__37_ <= r_n_117__37_;
      r_117__36_ <= r_n_117__36_;
      r_117__35_ <= r_n_117__35_;
      r_117__34_ <= r_n_117__34_;
      r_117__33_ <= r_n_117__33_;
      r_117__32_ <= r_n_117__32_;
      r_117__31_ <= r_n_117__31_;
      r_117__30_ <= r_n_117__30_;
      r_117__29_ <= r_n_117__29_;
      r_117__28_ <= r_n_117__28_;
      r_117__27_ <= r_n_117__27_;
      r_117__26_ <= r_n_117__26_;
      r_117__25_ <= r_n_117__25_;
      r_117__24_ <= r_n_117__24_;
      r_117__23_ <= r_n_117__23_;
      r_117__22_ <= r_n_117__22_;
      r_117__21_ <= r_n_117__21_;
      r_117__20_ <= r_n_117__20_;
      r_117__19_ <= r_n_117__19_;
      r_117__18_ <= r_n_117__18_;
      r_117__17_ <= r_n_117__17_;
      r_117__16_ <= r_n_117__16_;
      r_117__15_ <= r_n_117__15_;
      r_117__14_ <= r_n_117__14_;
      r_117__13_ <= r_n_117__13_;
      r_117__12_ <= r_n_117__12_;
      r_117__11_ <= r_n_117__11_;
      r_117__10_ <= r_n_117__10_;
      r_117__9_ <= r_n_117__9_;
      r_117__8_ <= r_n_117__8_;
      r_117__7_ <= r_n_117__7_;
      r_117__6_ <= r_n_117__6_;
      r_117__5_ <= r_n_117__5_;
      r_117__4_ <= r_n_117__4_;
      r_117__3_ <= r_n_117__3_;
      r_117__2_ <= r_n_117__2_;
      r_117__1_ <= r_n_117__1_;
      r_117__0_ <= r_n_117__0_;
    end 
    if(N3702) begin
      r_118__63_ <= r_n_118__63_;
      r_118__62_ <= r_n_118__62_;
      r_118__61_ <= r_n_118__61_;
      r_118__60_ <= r_n_118__60_;
      r_118__59_ <= r_n_118__59_;
      r_118__58_ <= r_n_118__58_;
      r_118__57_ <= r_n_118__57_;
      r_118__56_ <= r_n_118__56_;
      r_118__55_ <= r_n_118__55_;
      r_118__54_ <= r_n_118__54_;
      r_118__53_ <= r_n_118__53_;
      r_118__52_ <= r_n_118__52_;
      r_118__51_ <= r_n_118__51_;
      r_118__50_ <= r_n_118__50_;
      r_118__49_ <= r_n_118__49_;
      r_118__48_ <= r_n_118__48_;
      r_118__47_ <= r_n_118__47_;
      r_118__46_ <= r_n_118__46_;
      r_118__45_ <= r_n_118__45_;
      r_118__44_ <= r_n_118__44_;
      r_118__43_ <= r_n_118__43_;
      r_118__42_ <= r_n_118__42_;
      r_118__41_ <= r_n_118__41_;
      r_118__40_ <= r_n_118__40_;
      r_118__39_ <= r_n_118__39_;
      r_118__38_ <= r_n_118__38_;
      r_118__37_ <= r_n_118__37_;
      r_118__36_ <= r_n_118__36_;
      r_118__35_ <= r_n_118__35_;
      r_118__34_ <= r_n_118__34_;
      r_118__33_ <= r_n_118__33_;
      r_118__32_ <= r_n_118__32_;
      r_118__31_ <= r_n_118__31_;
      r_118__30_ <= r_n_118__30_;
      r_118__29_ <= r_n_118__29_;
      r_118__28_ <= r_n_118__28_;
      r_118__27_ <= r_n_118__27_;
      r_118__26_ <= r_n_118__26_;
      r_118__25_ <= r_n_118__25_;
      r_118__24_ <= r_n_118__24_;
      r_118__23_ <= r_n_118__23_;
      r_118__22_ <= r_n_118__22_;
      r_118__21_ <= r_n_118__21_;
      r_118__20_ <= r_n_118__20_;
      r_118__19_ <= r_n_118__19_;
      r_118__18_ <= r_n_118__18_;
      r_118__17_ <= r_n_118__17_;
      r_118__16_ <= r_n_118__16_;
      r_118__15_ <= r_n_118__15_;
      r_118__14_ <= r_n_118__14_;
      r_118__13_ <= r_n_118__13_;
      r_118__12_ <= r_n_118__12_;
      r_118__11_ <= r_n_118__11_;
      r_118__10_ <= r_n_118__10_;
      r_118__9_ <= r_n_118__9_;
      r_118__8_ <= r_n_118__8_;
      r_118__7_ <= r_n_118__7_;
      r_118__6_ <= r_n_118__6_;
      r_118__5_ <= r_n_118__5_;
      r_118__4_ <= r_n_118__4_;
      r_118__3_ <= r_n_118__3_;
      r_118__2_ <= r_n_118__2_;
      r_118__1_ <= r_n_118__1_;
      r_118__0_ <= r_n_118__0_;
    end 
    if(N3703) begin
      r_119__63_ <= r_n_119__63_;
      r_119__62_ <= r_n_119__62_;
      r_119__61_ <= r_n_119__61_;
      r_119__60_ <= r_n_119__60_;
      r_119__59_ <= r_n_119__59_;
      r_119__58_ <= r_n_119__58_;
      r_119__57_ <= r_n_119__57_;
      r_119__56_ <= r_n_119__56_;
      r_119__55_ <= r_n_119__55_;
      r_119__54_ <= r_n_119__54_;
      r_119__53_ <= r_n_119__53_;
      r_119__52_ <= r_n_119__52_;
      r_119__51_ <= r_n_119__51_;
      r_119__50_ <= r_n_119__50_;
      r_119__49_ <= r_n_119__49_;
      r_119__48_ <= r_n_119__48_;
      r_119__47_ <= r_n_119__47_;
      r_119__46_ <= r_n_119__46_;
      r_119__45_ <= r_n_119__45_;
      r_119__44_ <= r_n_119__44_;
      r_119__43_ <= r_n_119__43_;
      r_119__42_ <= r_n_119__42_;
      r_119__41_ <= r_n_119__41_;
      r_119__40_ <= r_n_119__40_;
      r_119__39_ <= r_n_119__39_;
      r_119__38_ <= r_n_119__38_;
      r_119__37_ <= r_n_119__37_;
      r_119__36_ <= r_n_119__36_;
      r_119__35_ <= r_n_119__35_;
      r_119__34_ <= r_n_119__34_;
      r_119__33_ <= r_n_119__33_;
      r_119__32_ <= r_n_119__32_;
      r_119__31_ <= r_n_119__31_;
      r_119__30_ <= r_n_119__30_;
      r_119__29_ <= r_n_119__29_;
      r_119__28_ <= r_n_119__28_;
      r_119__27_ <= r_n_119__27_;
      r_119__26_ <= r_n_119__26_;
      r_119__25_ <= r_n_119__25_;
      r_119__24_ <= r_n_119__24_;
      r_119__23_ <= r_n_119__23_;
      r_119__22_ <= r_n_119__22_;
      r_119__21_ <= r_n_119__21_;
      r_119__20_ <= r_n_119__20_;
      r_119__19_ <= r_n_119__19_;
      r_119__18_ <= r_n_119__18_;
      r_119__17_ <= r_n_119__17_;
      r_119__16_ <= r_n_119__16_;
      r_119__15_ <= r_n_119__15_;
      r_119__14_ <= r_n_119__14_;
      r_119__13_ <= r_n_119__13_;
      r_119__12_ <= r_n_119__12_;
      r_119__11_ <= r_n_119__11_;
      r_119__10_ <= r_n_119__10_;
      r_119__9_ <= r_n_119__9_;
      r_119__8_ <= r_n_119__8_;
      r_119__7_ <= r_n_119__7_;
      r_119__6_ <= r_n_119__6_;
      r_119__5_ <= r_n_119__5_;
      r_119__4_ <= r_n_119__4_;
      r_119__3_ <= r_n_119__3_;
      r_119__2_ <= r_n_119__2_;
      r_119__1_ <= r_n_119__1_;
      r_119__0_ <= r_n_119__0_;
    end 
    if(N3704) begin
      r_120__63_ <= r_n_120__63_;
      r_120__62_ <= r_n_120__62_;
      r_120__61_ <= r_n_120__61_;
      r_120__60_ <= r_n_120__60_;
      r_120__59_ <= r_n_120__59_;
      r_120__58_ <= r_n_120__58_;
      r_120__57_ <= r_n_120__57_;
      r_120__56_ <= r_n_120__56_;
      r_120__55_ <= r_n_120__55_;
      r_120__54_ <= r_n_120__54_;
      r_120__53_ <= r_n_120__53_;
      r_120__52_ <= r_n_120__52_;
      r_120__51_ <= r_n_120__51_;
      r_120__50_ <= r_n_120__50_;
      r_120__49_ <= r_n_120__49_;
      r_120__48_ <= r_n_120__48_;
      r_120__47_ <= r_n_120__47_;
      r_120__46_ <= r_n_120__46_;
      r_120__45_ <= r_n_120__45_;
      r_120__44_ <= r_n_120__44_;
      r_120__43_ <= r_n_120__43_;
      r_120__42_ <= r_n_120__42_;
      r_120__41_ <= r_n_120__41_;
      r_120__40_ <= r_n_120__40_;
      r_120__39_ <= r_n_120__39_;
      r_120__38_ <= r_n_120__38_;
      r_120__37_ <= r_n_120__37_;
      r_120__36_ <= r_n_120__36_;
      r_120__35_ <= r_n_120__35_;
      r_120__34_ <= r_n_120__34_;
      r_120__33_ <= r_n_120__33_;
      r_120__32_ <= r_n_120__32_;
      r_120__31_ <= r_n_120__31_;
      r_120__30_ <= r_n_120__30_;
      r_120__29_ <= r_n_120__29_;
      r_120__28_ <= r_n_120__28_;
      r_120__27_ <= r_n_120__27_;
      r_120__26_ <= r_n_120__26_;
      r_120__25_ <= r_n_120__25_;
      r_120__24_ <= r_n_120__24_;
      r_120__23_ <= r_n_120__23_;
      r_120__22_ <= r_n_120__22_;
      r_120__21_ <= r_n_120__21_;
      r_120__20_ <= r_n_120__20_;
      r_120__19_ <= r_n_120__19_;
      r_120__18_ <= r_n_120__18_;
      r_120__17_ <= r_n_120__17_;
      r_120__16_ <= r_n_120__16_;
      r_120__15_ <= r_n_120__15_;
      r_120__14_ <= r_n_120__14_;
      r_120__13_ <= r_n_120__13_;
      r_120__12_ <= r_n_120__12_;
      r_120__11_ <= r_n_120__11_;
      r_120__10_ <= r_n_120__10_;
      r_120__9_ <= r_n_120__9_;
      r_120__8_ <= r_n_120__8_;
      r_120__7_ <= r_n_120__7_;
      r_120__6_ <= r_n_120__6_;
      r_120__5_ <= r_n_120__5_;
      r_120__4_ <= r_n_120__4_;
      r_120__3_ <= r_n_120__3_;
      r_120__2_ <= r_n_120__2_;
      r_120__1_ <= r_n_120__1_;
      r_120__0_ <= r_n_120__0_;
    end 
    if(N3705) begin
      r_121__63_ <= r_n_121__63_;
      r_121__62_ <= r_n_121__62_;
      r_121__61_ <= r_n_121__61_;
      r_121__60_ <= r_n_121__60_;
      r_121__59_ <= r_n_121__59_;
      r_121__58_ <= r_n_121__58_;
      r_121__57_ <= r_n_121__57_;
      r_121__56_ <= r_n_121__56_;
      r_121__55_ <= r_n_121__55_;
      r_121__54_ <= r_n_121__54_;
      r_121__53_ <= r_n_121__53_;
      r_121__52_ <= r_n_121__52_;
      r_121__51_ <= r_n_121__51_;
      r_121__50_ <= r_n_121__50_;
      r_121__49_ <= r_n_121__49_;
      r_121__48_ <= r_n_121__48_;
      r_121__47_ <= r_n_121__47_;
      r_121__46_ <= r_n_121__46_;
      r_121__45_ <= r_n_121__45_;
      r_121__44_ <= r_n_121__44_;
      r_121__43_ <= r_n_121__43_;
      r_121__42_ <= r_n_121__42_;
      r_121__41_ <= r_n_121__41_;
      r_121__40_ <= r_n_121__40_;
      r_121__39_ <= r_n_121__39_;
      r_121__38_ <= r_n_121__38_;
      r_121__37_ <= r_n_121__37_;
      r_121__36_ <= r_n_121__36_;
      r_121__35_ <= r_n_121__35_;
      r_121__34_ <= r_n_121__34_;
      r_121__33_ <= r_n_121__33_;
      r_121__32_ <= r_n_121__32_;
      r_121__31_ <= r_n_121__31_;
      r_121__30_ <= r_n_121__30_;
      r_121__29_ <= r_n_121__29_;
      r_121__28_ <= r_n_121__28_;
      r_121__27_ <= r_n_121__27_;
      r_121__26_ <= r_n_121__26_;
      r_121__25_ <= r_n_121__25_;
      r_121__24_ <= r_n_121__24_;
      r_121__23_ <= r_n_121__23_;
      r_121__22_ <= r_n_121__22_;
      r_121__21_ <= r_n_121__21_;
      r_121__20_ <= r_n_121__20_;
      r_121__19_ <= r_n_121__19_;
      r_121__18_ <= r_n_121__18_;
      r_121__17_ <= r_n_121__17_;
      r_121__16_ <= r_n_121__16_;
      r_121__15_ <= r_n_121__15_;
      r_121__14_ <= r_n_121__14_;
      r_121__13_ <= r_n_121__13_;
      r_121__12_ <= r_n_121__12_;
      r_121__11_ <= r_n_121__11_;
      r_121__10_ <= r_n_121__10_;
      r_121__9_ <= r_n_121__9_;
      r_121__8_ <= r_n_121__8_;
      r_121__7_ <= r_n_121__7_;
      r_121__6_ <= r_n_121__6_;
      r_121__5_ <= r_n_121__5_;
      r_121__4_ <= r_n_121__4_;
      r_121__3_ <= r_n_121__3_;
      r_121__2_ <= r_n_121__2_;
      r_121__1_ <= r_n_121__1_;
      r_121__0_ <= r_n_121__0_;
    end 
    if(N3706) begin
      r_122__63_ <= r_n_122__63_;
      r_122__62_ <= r_n_122__62_;
      r_122__61_ <= r_n_122__61_;
      r_122__60_ <= r_n_122__60_;
      r_122__59_ <= r_n_122__59_;
      r_122__58_ <= r_n_122__58_;
      r_122__57_ <= r_n_122__57_;
      r_122__56_ <= r_n_122__56_;
      r_122__55_ <= r_n_122__55_;
      r_122__54_ <= r_n_122__54_;
      r_122__53_ <= r_n_122__53_;
      r_122__52_ <= r_n_122__52_;
      r_122__51_ <= r_n_122__51_;
      r_122__50_ <= r_n_122__50_;
      r_122__49_ <= r_n_122__49_;
      r_122__48_ <= r_n_122__48_;
      r_122__47_ <= r_n_122__47_;
      r_122__46_ <= r_n_122__46_;
      r_122__45_ <= r_n_122__45_;
      r_122__44_ <= r_n_122__44_;
      r_122__43_ <= r_n_122__43_;
      r_122__42_ <= r_n_122__42_;
      r_122__41_ <= r_n_122__41_;
      r_122__40_ <= r_n_122__40_;
      r_122__39_ <= r_n_122__39_;
      r_122__38_ <= r_n_122__38_;
      r_122__37_ <= r_n_122__37_;
      r_122__36_ <= r_n_122__36_;
      r_122__35_ <= r_n_122__35_;
      r_122__34_ <= r_n_122__34_;
      r_122__33_ <= r_n_122__33_;
      r_122__32_ <= r_n_122__32_;
      r_122__31_ <= r_n_122__31_;
      r_122__30_ <= r_n_122__30_;
      r_122__29_ <= r_n_122__29_;
      r_122__28_ <= r_n_122__28_;
      r_122__27_ <= r_n_122__27_;
      r_122__26_ <= r_n_122__26_;
      r_122__25_ <= r_n_122__25_;
      r_122__24_ <= r_n_122__24_;
      r_122__23_ <= r_n_122__23_;
      r_122__22_ <= r_n_122__22_;
      r_122__21_ <= r_n_122__21_;
      r_122__20_ <= r_n_122__20_;
      r_122__19_ <= r_n_122__19_;
      r_122__18_ <= r_n_122__18_;
      r_122__17_ <= r_n_122__17_;
      r_122__16_ <= r_n_122__16_;
      r_122__15_ <= r_n_122__15_;
      r_122__14_ <= r_n_122__14_;
      r_122__13_ <= r_n_122__13_;
      r_122__12_ <= r_n_122__12_;
      r_122__11_ <= r_n_122__11_;
      r_122__10_ <= r_n_122__10_;
      r_122__9_ <= r_n_122__9_;
      r_122__8_ <= r_n_122__8_;
      r_122__7_ <= r_n_122__7_;
      r_122__6_ <= r_n_122__6_;
      r_122__5_ <= r_n_122__5_;
      r_122__4_ <= r_n_122__4_;
      r_122__3_ <= r_n_122__3_;
      r_122__2_ <= r_n_122__2_;
      r_122__1_ <= r_n_122__1_;
      r_122__0_ <= r_n_122__0_;
    end 
    if(N3707) begin
      r_123__63_ <= r_n_123__63_;
      r_123__62_ <= r_n_123__62_;
      r_123__61_ <= r_n_123__61_;
      r_123__60_ <= r_n_123__60_;
      r_123__59_ <= r_n_123__59_;
      r_123__58_ <= r_n_123__58_;
      r_123__57_ <= r_n_123__57_;
      r_123__56_ <= r_n_123__56_;
      r_123__55_ <= r_n_123__55_;
      r_123__54_ <= r_n_123__54_;
      r_123__53_ <= r_n_123__53_;
      r_123__52_ <= r_n_123__52_;
      r_123__51_ <= r_n_123__51_;
      r_123__50_ <= r_n_123__50_;
      r_123__49_ <= r_n_123__49_;
      r_123__48_ <= r_n_123__48_;
      r_123__47_ <= r_n_123__47_;
      r_123__46_ <= r_n_123__46_;
      r_123__45_ <= r_n_123__45_;
      r_123__44_ <= r_n_123__44_;
      r_123__43_ <= r_n_123__43_;
      r_123__42_ <= r_n_123__42_;
      r_123__41_ <= r_n_123__41_;
      r_123__40_ <= r_n_123__40_;
      r_123__39_ <= r_n_123__39_;
      r_123__38_ <= r_n_123__38_;
      r_123__37_ <= r_n_123__37_;
      r_123__36_ <= r_n_123__36_;
      r_123__35_ <= r_n_123__35_;
      r_123__34_ <= r_n_123__34_;
      r_123__33_ <= r_n_123__33_;
      r_123__32_ <= r_n_123__32_;
      r_123__31_ <= r_n_123__31_;
      r_123__30_ <= r_n_123__30_;
      r_123__29_ <= r_n_123__29_;
      r_123__28_ <= r_n_123__28_;
      r_123__27_ <= r_n_123__27_;
      r_123__26_ <= r_n_123__26_;
      r_123__25_ <= r_n_123__25_;
      r_123__24_ <= r_n_123__24_;
      r_123__23_ <= r_n_123__23_;
      r_123__22_ <= r_n_123__22_;
      r_123__21_ <= r_n_123__21_;
      r_123__20_ <= r_n_123__20_;
      r_123__19_ <= r_n_123__19_;
      r_123__18_ <= r_n_123__18_;
      r_123__17_ <= r_n_123__17_;
      r_123__16_ <= r_n_123__16_;
      r_123__15_ <= r_n_123__15_;
      r_123__14_ <= r_n_123__14_;
      r_123__13_ <= r_n_123__13_;
      r_123__12_ <= r_n_123__12_;
      r_123__11_ <= r_n_123__11_;
      r_123__10_ <= r_n_123__10_;
      r_123__9_ <= r_n_123__9_;
      r_123__8_ <= r_n_123__8_;
      r_123__7_ <= r_n_123__7_;
      r_123__6_ <= r_n_123__6_;
      r_123__5_ <= r_n_123__5_;
      r_123__4_ <= r_n_123__4_;
      r_123__3_ <= r_n_123__3_;
      r_123__2_ <= r_n_123__2_;
      r_123__1_ <= r_n_123__1_;
      r_123__0_ <= r_n_123__0_;
    end 
    if(N3708) begin
      r_124__63_ <= r_n_124__63_;
      r_124__62_ <= r_n_124__62_;
      r_124__61_ <= r_n_124__61_;
      r_124__60_ <= r_n_124__60_;
      r_124__59_ <= r_n_124__59_;
      r_124__58_ <= r_n_124__58_;
      r_124__57_ <= r_n_124__57_;
      r_124__56_ <= r_n_124__56_;
      r_124__55_ <= r_n_124__55_;
      r_124__54_ <= r_n_124__54_;
      r_124__53_ <= r_n_124__53_;
      r_124__52_ <= r_n_124__52_;
      r_124__51_ <= r_n_124__51_;
      r_124__50_ <= r_n_124__50_;
      r_124__49_ <= r_n_124__49_;
      r_124__48_ <= r_n_124__48_;
      r_124__47_ <= r_n_124__47_;
      r_124__46_ <= r_n_124__46_;
      r_124__45_ <= r_n_124__45_;
      r_124__44_ <= r_n_124__44_;
      r_124__43_ <= r_n_124__43_;
      r_124__42_ <= r_n_124__42_;
      r_124__41_ <= r_n_124__41_;
      r_124__40_ <= r_n_124__40_;
      r_124__39_ <= r_n_124__39_;
      r_124__38_ <= r_n_124__38_;
      r_124__37_ <= r_n_124__37_;
      r_124__36_ <= r_n_124__36_;
      r_124__35_ <= r_n_124__35_;
      r_124__34_ <= r_n_124__34_;
      r_124__33_ <= r_n_124__33_;
      r_124__32_ <= r_n_124__32_;
      r_124__31_ <= r_n_124__31_;
      r_124__30_ <= r_n_124__30_;
      r_124__29_ <= r_n_124__29_;
      r_124__28_ <= r_n_124__28_;
      r_124__27_ <= r_n_124__27_;
      r_124__26_ <= r_n_124__26_;
      r_124__25_ <= r_n_124__25_;
      r_124__24_ <= r_n_124__24_;
      r_124__23_ <= r_n_124__23_;
      r_124__22_ <= r_n_124__22_;
      r_124__21_ <= r_n_124__21_;
      r_124__20_ <= r_n_124__20_;
      r_124__19_ <= r_n_124__19_;
      r_124__18_ <= r_n_124__18_;
      r_124__17_ <= r_n_124__17_;
      r_124__16_ <= r_n_124__16_;
      r_124__15_ <= r_n_124__15_;
      r_124__14_ <= r_n_124__14_;
      r_124__13_ <= r_n_124__13_;
      r_124__12_ <= r_n_124__12_;
      r_124__11_ <= r_n_124__11_;
      r_124__10_ <= r_n_124__10_;
      r_124__9_ <= r_n_124__9_;
      r_124__8_ <= r_n_124__8_;
      r_124__7_ <= r_n_124__7_;
      r_124__6_ <= r_n_124__6_;
      r_124__5_ <= r_n_124__5_;
      r_124__4_ <= r_n_124__4_;
      r_124__3_ <= r_n_124__3_;
      r_124__2_ <= r_n_124__2_;
      r_124__1_ <= r_n_124__1_;
      r_124__0_ <= r_n_124__0_;
    end 
    if(N3709) begin
      r_125__63_ <= r_n_125__63_;
      r_125__62_ <= r_n_125__62_;
      r_125__61_ <= r_n_125__61_;
      r_125__60_ <= r_n_125__60_;
      r_125__59_ <= r_n_125__59_;
      r_125__58_ <= r_n_125__58_;
      r_125__57_ <= r_n_125__57_;
      r_125__56_ <= r_n_125__56_;
      r_125__55_ <= r_n_125__55_;
      r_125__54_ <= r_n_125__54_;
      r_125__53_ <= r_n_125__53_;
      r_125__52_ <= r_n_125__52_;
      r_125__51_ <= r_n_125__51_;
      r_125__50_ <= r_n_125__50_;
      r_125__49_ <= r_n_125__49_;
      r_125__48_ <= r_n_125__48_;
      r_125__47_ <= r_n_125__47_;
      r_125__46_ <= r_n_125__46_;
      r_125__45_ <= r_n_125__45_;
      r_125__44_ <= r_n_125__44_;
      r_125__43_ <= r_n_125__43_;
      r_125__42_ <= r_n_125__42_;
      r_125__41_ <= r_n_125__41_;
      r_125__40_ <= r_n_125__40_;
      r_125__39_ <= r_n_125__39_;
      r_125__38_ <= r_n_125__38_;
      r_125__37_ <= r_n_125__37_;
      r_125__36_ <= r_n_125__36_;
      r_125__35_ <= r_n_125__35_;
      r_125__34_ <= r_n_125__34_;
      r_125__33_ <= r_n_125__33_;
      r_125__32_ <= r_n_125__32_;
      r_125__31_ <= r_n_125__31_;
      r_125__30_ <= r_n_125__30_;
      r_125__29_ <= r_n_125__29_;
      r_125__28_ <= r_n_125__28_;
      r_125__27_ <= r_n_125__27_;
      r_125__26_ <= r_n_125__26_;
      r_125__25_ <= r_n_125__25_;
      r_125__24_ <= r_n_125__24_;
      r_125__23_ <= r_n_125__23_;
      r_125__22_ <= r_n_125__22_;
      r_125__21_ <= r_n_125__21_;
      r_125__20_ <= r_n_125__20_;
      r_125__19_ <= r_n_125__19_;
      r_125__18_ <= r_n_125__18_;
      r_125__17_ <= r_n_125__17_;
      r_125__16_ <= r_n_125__16_;
      r_125__15_ <= r_n_125__15_;
      r_125__14_ <= r_n_125__14_;
      r_125__13_ <= r_n_125__13_;
      r_125__12_ <= r_n_125__12_;
      r_125__11_ <= r_n_125__11_;
      r_125__10_ <= r_n_125__10_;
      r_125__9_ <= r_n_125__9_;
      r_125__8_ <= r_n_125__8_;
      r_125__7_ <= r_n_125__7_;
      r_125__6_ <= r_n_125__6_;
      r_125__5_ <= r_n_125__5_;
      r_125__4_ <= r_n_125__4_;
      r_125__3_ <= r_n_125__3_;
      r_125__2_ <= r_n_125__2_;
      r_125__1_ <= r_n_125__1_;
      r_125__0_ <= r_n_125__0_;
    end 
    if(N3710) begin
      r_126__63_ <= r_n_126__63_;
      r_126__62_ <= r_n_126__62_;
      r_126__61_ <= r_n_126__61_;
      r_126__60_ <= r_n_126__60_;
      r_126__59_ <= r_n_126__59_;
      r_126__58_ <= r_n_126__58_;
      r_126__57_ <= r_n_126__57_;
      r_126__56_ <= r_n_126__56_;
      r_126__55_ <= r_n_126__55_;
      r_126__54_ <= r_n_126__54_;
      r_126__53_ <= r_n_126__53_;
      r_126__52_ <= r_n_126__52_;
      r_126__51_ <= r_n_126__51_;
      r_126__50_ <= r_n_126__50_;
      r_126__49_ <= r_n_126__49_;
      r_126__48_ <= r_n_126__48_;
      r_126__47_ <= r_n_126__47_;
      r_126__46_ <= r_n_126__46_;
      r_126__45_ <= r_n_126__45_;
      r_126__44_ <= r_n_126__44_;
      r_126__43_ <= r_n_126__43_;
      r_126__42_ <= r_n_126__42_;
      r_126__41_ <= r_n_126__41_;
      r_126__40_ <= r_n_126__40_;
      r_126__39_ <= r_n_126__39_;
      r_126__38_ <= r_n_126__38_;
      r_126__37_ <= r_n_126__37_;
      r_126__36_ <= r_n_126__36_;
      r_126__35_ <= r_n_126__35_;
      r_126__34_ <= r_n_126__34_;
      r_126__33_ <= r_n_126__33_;
      r_126__32_ <= r_n_126__32_;
      r_126__31_ <= r_n_126__31_;
      r_126__30_ <= r_n_126__30_;
      r_126__29_ <= r_n_126__29_;
      r_126__28_ <= r_n_126__28_;
      r_126__27_ <= r_n_126__27_;
      r_126__26_ <= r_n_126__26_;
      r_126__25_ <= r_n_126__25_;
      r_126__24_ <= r_n_126__24_;
      r_126__23_ <= r_n_126__23_;
      r_126__22_ <= r_n_126__22_;
      r_126__21_ <= r_n_126__21_;
      r_126__20_ <= r_n_126__20_;
      r_126__19_ <= r_n_126__19_;
      r_126__18_ <= r_n_126__18_;
      r_126__17_ <= r_n_126__17_;
      r_126__16_ <= r_n_126__16_;
      r_126__15_ <= r_n_126__15_;
      r_126__14_ <= r_n_126__14_;
      r_126__13_ <= r_n_126__13_;
      r_126__12_ <= r_n_126__12_;
      r_126__11_ <= r_n_126__11_;
      r_126__10_ <= r_n_126__10_;
      r_126__9_ <= r_n_126__9_;
      r_126__8_ <= r_n_126__8_;
      r_126__7_ <= r_n_126__7_;
      r_126__6_ <= r_n_126__6_;
      r_126__5_ <= r_n_126__5_;
      r_126__4_ <= r_n_126__4_;
      r_126__3_ <= r_n_126__3_;
      r_126__2_ <= r_n_126__2_;
      r_126__1_ <= r_n_126__1_;
      r_126__0_ <= r_n_126__0_;
    end 
    if(N3711) begin
      r_127__63_ <= r_n_127__63_;
      r_127__62_ <= r_n_127__62_;
      r_127__61_ <= r_n_127__61_;
      r_127__60_ <= r_n_127__60_;
      r_127__59_ <= r_n_127__59_;
      r_127__58_ <= r_n_127__58_;
      r_127__57_ <= r_n_127__57_;
      r_127__56_ <= r_n_127__56_;
      r_127__55_ <= r_n_127__55_;
      r_127__54_ <= r_n_127__54_;
      r_127__53_ <= r_n_127__53_;
      r_127__52_ <= r_n_127__52_;
      r_127__51_ <= r_n_127__51_;
      r_127__50_ <= r_n_127__50_;
      r_127__49_ <= r_n_127__49_;
      r_127__48_ <= r_n_127__48_;
      r_127__47_ <= r_n_127__47_;
      r_127__46_ <= r_n_127__46_;
      r_127__45_ <= r_n_127__45_;
      r_127__44_ <= r_n_127__44_;
      r_127__43_ <= r_n_127__43_;
      r_127__42_ <= r_n_127__42_;
      r_127__41_ <= r_n_127__41_;
      r_127__40_ <= r_n_127__40_;
      r_127__39_ <= r_n_127__39_;
      r_127__38_ <= r_n_127__38_;
      r_127__37_ <= r_n_127__37_;
      r_127__36_ <= r_n_127__36_;
      r_127__35_ <= r_n_127__35_;
      r_127__34_ <= r_n_127__34_;
      r_127__33_ <= r_n_127__33_;
      r_127__32_ <= r_n_127__32_;
      r_127__31_ <= r_n_127__31_;
      r_127__30_ <= r_n_127__30_;
      r_127__29_ <= r_n_127__29_;
      r_127__28_ <= r_n_127__28_;
      r_127__27_ <= r_n_127__27_;
      r_127__26_ <= r_n_127__26_;
      r_127__25_ <= r_n_127__25_;
      r_127__24_ <= r_n_127__24_;
      r_127__23_ <= r_n_127__23_;
      r_127__22_ <= r_n_127__22_;
      r_127__21_ <= r_n_127__21_;
      r_127__20_ <= r_n_127__20_;
      r_127__19_ <= r_n_127__19_;
      r_127__18_ <= r_n_127__18_;
      r_127__17_ <= r_n_127__17_;
      r_127__16_ <= r_n_127__16_;
      r_127__15_ <= r_n_127__15_;
      r_127__14_ <= r_n_127__14_;
      r_127__13_ <= r_n_127__13_;
      r_127__12_ <= r_n_127__12_;
      r_127__11_ <= r_n_127__11_;
      r_127__10_ <= r_n_127__10_;
      r_127__9_ <= r_n_127__9_;
      r_127__8_ <= r_n_127__8_;
      r_127__7_ <= r_n_127__7_;
      r_127__6_ <= r_n_127__6_;
      r_127__5_ <= r_n_127__5_;
      r_127__4_ <= r_n_127__4_;
      r_127__3_ <= r_n_127__3_;
      r_127__2_ <= r_n_127__2_;
      r_127__1_ <= r_n_127__1_;
      r_127__0_ <= r_n_127__0_;
    end 
    if(N3712) begin
      r_128__63_ <= r_n_128__63_;
      r_128__62_ <= r_n_128__62_;
      r_128__61_ <= r_n_128__61_;
      r_128__60_ <= r_n_128__60_;
      r_128__59_ <= r_n_128__59_;
      r_128__58_ <= r_n_128__58_;
      r_128__57_ <= r_n_128__57_;
      r_128__56_ <= r_n_128__56_;
      r_128__55_ <= r_n_128__55_;
      r_128__54_ <= r_n_128__54_;
      r_128__53_ <= r_n_128__53_;
      r_128__52_ <= r_n_128__52_;
      r_128__51_ <= r_n_128__51_;
      r_128__50_ <= r_n_128__50_;
      r_128__49_ <= r_n_128__49_;
      r_128__48_ <= r_n_128__48_;
      r_128__47_ <= r_n_128__47_;
      r_128__46_ <= r_n_128__46_;
      r_128__45_ <= r_n_128__45_;
      r_128__44_ <= r_n_128__44_;
      r_128__43_ <= r_n_128__43_;
      r_128__42_ <= r_n_128__42_;
      r_128__41_ <= r_n_128__41_;
      r_128__40_ <= r_n_128__40_;
      r_128__39_ <= r_n_128__39_;
      r_128__38_ <= r_n_128__38_;
      r_128__37_ <= r_n_128__37_;
      r_128__36_ <= r_n_128__36_;
      r_128__35_ <= r_n_128__35_;
      r_128__34_ <= r_n_128__34_;
      r_128__33_ <= r_n_128__33_;
      r_128__32_ <= r_n_128__32_;
      r_128__31_ <= r_n_128__31_;
      r_128__30_ <= r_n_128__30_;
      r_128__29_ <= r_n_128__29_;
      r_128__28_ <= r_n_128__28_;
      r_128__27_ <= r_n_128__27_;
      r_128__26_ <= r_n_128__26_;
      r_128__25_ <= r_n_128__25_;
      r_128__24_ <= r_n_128__24_;
      r_128__23_ <= r_n_128__23_;
      r_128__22_ <= r_n_128__22_;
      r_128__21_ <= r_n_128__21_;
      r_128__20_ <= r_n_128__20_;
      r_128__19_ <= r_n_128__19_;
      r_128__18_ <= r_n_128__18_;
      r_128__17_ <= r_n_128__17_;
      r_128__16_ <= r_n_128__16_;
      r_128__15_ <= r_n_128__15_;
      r_128__14_ <= r_n_128__14_;
      r_128__13_ <= r_n_128__13_;
      r_128__12_ <= r_n_128__12_;
      r_128__11_ <= r_n_128__11_;
      r_128__10_ <= r_n_128__10_;
      r_128__9_ <= r_n_128__9_;
      r_128__8_ <= r_n_128__8_;
      r_128__7_ <= r_n_128__7_;
      r_128__6_ <= r_n_128__6_;
      r_128__5_ <= r_n_128__5_;
      r_128__4_ <= r_n_128__4_;
      r_128__3_ <= r_n_128__3_;
      r_128__2_ <= r_n_128__2_;
      r_128__1_ <= r_n_128__1_;
      r_128__0_ <= r_n_128__0_;
    end 
    if(N3713) begin
      r_129__63_ <= r_n_129__63_;
      r_129__62_ <= r_n_129__62_;
      r_129__61_ <= r_n_129__61_;
      r_129__60_ <= r_n_129__60_;
      r_129__59_ <= r_n_129__59_;
      r_129__58_ <= r_n_129__58_;
      r_129__57_ <= r_n_129__57_;
      r_129__56_ <= r_n_129__56_;
      r_129__55_ <= r_n_129__55_;
      r_129__54_ <= r_n_129__54_;
      r_129__53_ <= r_n_129__53_;
      r_129__52_ <= r_n_129__52_;
      r_129__51_ <= r_n_129__51_;
      r_129__50_ <= r_n_129__50_;
      r_129__49_ <= r_n_129__49_;
      r_129__48_ <= r_n_129__48_;
      r_129__47_ <= r_n_129__47_;
      r_129__46_ <= r_n_129__46_;
      r_129__45_ <= r_n_129__45_;
      r_129__44_ <= r_n_129__44_;
      r_129__43_ <= r_n_129__43_;
      r_129__42_ <= r_n_129__42_;
      r_129__41_ <= r_n_129__41_;
      r_129__40_ <= r_n_129__40_;
      r_129__39_ <= r_n_129__39_;
      r_129__38_ <= r_n_129__38_;
      r_129__37_ <= r_n_129__37_;
      r_129__36_ <= r_n_129__36_;
      r_129__35_ <= r_n_129__35_;
      r_129__34_ <= r_n_129__34_;
      r_129__33_ <= r_n_129__33_;
      r_129__32_ <= r_n_129__32_;
      r_129__31_ <= r_n_129__31_;
      r_129__30_ <= r_n_129__30_;
      r_129__29_ <= r_n_129__29_;
      r_129__28_ <= r_n_129__28_;
      r_129__27_ <= r_n_129__27_;
      r_129__26_ <= r_n_129__26_;
      r_129__25_ <= r_n_129__25_;
      r_129__24_ <= r_n_129__24_;
      r_129__23_ <= r_n_129__23_;
      r_129__22_ <= r_n_129__22_;
      r_129__21_ <= r_n_129__21_;
      r_129__20_ <= r_n_129__20_;
      r_129__19_ <= r_n_129__19_;
      r_129__18_ <= r_n_129__18_;
      r_129__17_ <= r_n_129__17_;
      r_129__16_ <= r_n_129__16_;
      r_129__15_ <= r_n_129__15_;
      r_129__14_ <= r_n_129__14_;
      r_129__13_ <= r_n_129__13_;
      r_129__12_ <= r_n_129__12_;
      r_129__11_ <= r_n_129__11_;
      r_129__10_ <= r_n_129__10_;
      r_129__9_ <= r_n_129__9_;
      r_129__8_ <= r_n_129__8_;
      r_129__7_ <= r_n_129__7_;
      r_129__6_ <= r_n_129__6_;
      r_129__5_ <= r_n_129__5_;
      r_129__4_ <= r_n_129__4_;
      r_129__3_ <= r_n_129__3_;
      r_129__2_ <= r_n_129__2_;
      r_129__1_ <= r_n_129__1_;
      r_129__0_ <= r_n_129__0_;
    end 
    if(N3714) begin
      r_130__63_ <= r_n_130__63_;
      r_130__62_ <= r_n_130__62_;
      r_130__61_ <= r_n_130__61_;
      r_130__60_ <= r_n_130__60_;
      r_130__59_ <= r_n_130__59_;
      r_130__58_ <= r_n_130__58_;
      r_130__57_ <= r_n_130__57_;
      r_130__56_ <= r_n_130__56_;
      r_130__55_ <= r_n_130__55_;
      r_130__54_ <= r_n_130__54_;
      r_130__53_ <= r_n_130__53_;
      r_130__52_ <= r_n_130__52_;
      r_130__51_ <= r_n_130__51_;
      r_130__50_ <= r_n_130__50_;
      r_130__49_ <= r_n_130__49_;
      r_130__48_ <= r_n_130__48_;
      r_130__47_ <= r_n_130__47_;
      r_130__46_ <= r_n_130__46_;
      r_130__45_ <= r_n_130__45_;
      r_130__44_ <= r_n_130__44_;
      r_130__43_ <= r_n_130__43_;
      r_130__42_ <= r_n_130__42_;
      r_130__41_ <= r_n_130__41_;
      r_130__40_ <= r_n_130__40_;
      r_130__39_ <= r_n_130__39_;
      r_130__38_ <= r_n_130__38_;
      r_130__37_ <= r_n_130__37_;
      r_130__36_ <= r_n_130__36_;
      r_130__35_ <= r_n_130__35_;
      r_130__34_ <= r_n_130__34_;
      r_130__33_ <= r_n_130__33_;
      r_130__32_ <= r_n_130__32_;
      r_130__31_ <= r_n_130__31_;
      r_130__30_ <= r_n_130__30_;
      r_130__29_ <= r_n_130__29_;
      r_130__28_ <= r_n_130__28_;
      r_130__27_ <= r_n_130__27_;
      r_130__26_ <= r_n_130__26_;
      r_130__25_ <= r_n_130__25_;
      r_130__24_ <= r_n_130__24_;
      r_130__23_ <= r_n_130__23_;
      r_130__22_ <= r_n_130__22_;
      r_130__21_ <= r_n_130__21_;
      r_130__20_ <= r_n_130__20_;
      r_130__19_ <= r_n_130__19_;
      r_130__18_ <= r_n_130__18_;
      r_130__17_ <= r_n_130__17_;
      r_130__16_ <= r_n_130__16_;
      r_130__15_ <= r_n_130__15_;
      r_130__14_ <= r_n_130__14_;
      r_130__13_ <= r_n_130__13_;
      r_130__12_ <= r_n_130__12_;
      r_130__11_ <= r_n_130__11_;
      r_130__10_ <= r_n_130__10_;
      r_130__9_ <= r_n_130__9_;
      r_130__8_ <= r_n_130__8_;
      r_130__7_ <= r_n_130__7_;
      r_130__6_ <= r_n_130__6_;
      r_130__5_ <= r_n_130__5_;
      r_130__4_ <= r_n_130__4_;
      r_130__3_ <= r_n_130__3_;
      r_130__2_ <= r_n_130__2_;
      r_130__1_ <= r_n_130__1_;
      r_130__0_ <= r_n_130__0_;
    end 
    if(N3715) begin
      r_131__63_ <= r_n_131__63_;
      r_131__62_ <= r_n_131__62_;
      r_131__61_ <= r_n_131__61_;
      r_131__60_ <= r_n_131__60_;
      r_131__59_ <= r_n_131__59_;
      r_131__58_ <= r_n_131__58_;
      r_131__57_ <= r_n_131__57_;
      r_131__56_ <= r_n_131__56_;
      r_131__55_ <= r_n_131__55_;
      r_131__54_ <= r_n_131__54_;
      r_131__53_ <= r_n_131__53_;
      r_131__52_ <= r_n_131__52_;
      r_131__51_ <= r_n_131__51_;
      r_131__50_ <= r_n_131__50_;
      r_131__49_ <= r_n_131__49_;
      r_131__48_ <= r_n_131__48_;
      r_131__47_ <= r_n_131__47_;
      r_131__46_ <= r_n_131__46_;
      r_131__45_ <= r_n_131__45_;
      r_131__44_ <= r_n_131__44_;
      r_131__43_ <= r_n_131__43_;
      r_131__42_ <= r_n_131__42_;
      r_131__41_ <= r_n_131__41_;
      r_131__40_ <= r_n_131__40_;
      r_131__39_ <= r_n_131__39_;
      r_131__38_ <= r_n_131__38_;
      r_131__37_ <= r_n_131__37_;
      r_131__36_ <= r_n_131__36_;
      r_131__35_ <= r_n_131__35_;
      r_131__34_ <= r_n_131__34_;
      r_131__33_ <= r_n_131__33_;
      r_131__32_ <= r_n_131__32_;
      r_131__31_ <= r_n_131__31_;
      r_131__30_ <= r_n_131__30_;
      r_131__29_ <= r_n_131__29_;
      r_131__28_ <= r_n_131__28_;
      r_131__27_ <= r_n_131__27_;
      r_131__26_ <= r_n_131__26_;
      r_131__25_ <= r_n_131__25_;
      r_131__24_ <= r_n_131__24_;
      r_131__23_ <= r_n_131__23_;
      r_131__22_ <= r_n_131__22_;
      r_131__21_ <= r_n_131__21_;
      r_131__20_ <= r_n_131__20_;
      r_131__19_ <= r_n_131__19_;
      r_131__18_ <= r_n_131__18_;
      r_131__17_ <= r_n_131__17_;
      r_131__16_ <= r_n_131__16_;
      r_131__15_ <= r_n_131__15_;
      r_131__14_ <= r_n_131__14_;
      r_131__13_ <= r_n_131__13_;
      r_131__12_ <= r_n_131__12_;
      r_131__11_ <= r_n_131__11_;
      r_131__10_ <= r_n_131__10_;
      r_131__9_ <= r_n_131__9_;
      r_131__8_ <= r_n_131__8_;
      r_131__7_ <= r_n_131__7_;
      r_131__6_ <= r_n_131__6_;
      r_131__5_ <= r_n_131__5_;
      r_131__4_ <= r_n_131__4_;
      r_131__3_ <= r_n_131__3_;
      r_131__2_ <= r_n_131__2_;
      r_131__1_ <= r_n_131__1_;
      r_131__0_ <= r_n_131__0_;
    end 
    if(N3716) begin
      r_132__63_ <= r_n_132__63_;
      r_132__62_ <= r_n_132__62_;
      r_132__61_ <= r_n_132__61_;
      r_132__60_ <= r_n_132__60_;
      r_132__59_ <= r_n_132__59_;
      r_132__58_ <= r_n_132__58_;
      r_132__57_ <= r_n_132__57_;
      r_132__56_ <= r_n_132__56_;
      r_132__55_ <= r_n_132__55_;
      r_132__54_ <= r_n_132__54_;
      r_132__53_ <= r_n_132__53_;
      r_132__52_ <= r_n_132__52_;
      r_132__51_ <= r_n_132__51_;
      r_132__50_ <= r_n_132__50_;
      r_132__49_ <= r_n_132__49_;
      r_132__48_ <= r_n_132__48_;
      r_132__47_ <= r_n_132__47_;
      r_132__46_ <= r_n_132__46_;
      r_132__45_ <= r_n_132__45_;
      r_132__44_ <= r_n_132__44_;
      r_132__43_ <= r_n_132__43_;
      r_132__42_ <= r_n_132__42_;
      r_132__41_ <= r_n_132__41_;
      r_132__40_ <= r_n_132__40_;
      r_132__39_ <= r_n_132__39_;
      r_132__38_ <= r_n_132__38_;
      r_132__37_ <= r_n_132__37_;
      r_132__36_ <= r_n_132__36_;
      r_132__35_ <= r_n_132__35_;
      r_132__34_ <= r_n_132__34_;
      r_132__33_ <= r_n_132__33_;
      r_132__32_ <= r_n_132__32_;
      r_132__31_ <= r_n_132__31_;
      r_132__30_ <= r_n_132__30_;
      r_132__29_ <= r_n_132__29_;
      r_132__28_ <= r_n_132__28_;
      r_132__27_ <= r_n_132__27_;
      r_132__26_ <= r_n_132__26_;
      r_132__25_ <= r_n_132__25_;
      r_132__24_ <= r_n_132__24_;
      r_132__23_ <= r_n_132__23_;
      r_132__22_ <= r_n_132__22_;
      r_132__21_ <= r_n_132__21_;
      r_132__20_ <= r_n_132__20_;
      r_132__19_ <= r_n_132__19_;
      r_132__18_ <= r_n_132__18_;
      r_132__17_ <= r_n_132__17_;
      r_132__16_ <= r_n_132__16_;
      r_132__15_ <= r_n_132__15_;
      r_132__14_ <= r_n_132__14_;
      r_132__13_ <= r_n_132__13_;
      r_132__12_ <= r_n_132__12_;
      r_132__11_ <= r_n_132__11_;
      r_132__10_ <= r_n_132__10_;
      r_132__9_ <= r_n_132__9_;
      r_132__8_ <= r_n_132__8_;
      r_132__7_ <= r_n_132__7_;
      r_132__6_ <= r_n_132__6_;
      r_132__5_ <= r_n_132__5_;
      r_132__4_ <= r_n_132__4_;
      r_132__3_ <= r_n_132__3_;
      r_132__2_ <= r_n_132__2_;
      r_132__1_ <= r_n_132__1_;
      r_132__0_ <= r_n_132__0_;
    end 
    if(N3717) begin
      r_133__63_ <= r_n_133__63_;
      r_133__62_ <= r_n_133__62_;
      r_133__61_ <= r_n_133__61_;
      r_133__60_ <= r_n_133__60_;
      r_133__59_ <= r_n_133__59_;
      r_133__58_ <= r_n_133__58_;
      r_133__57_ <= r_n_133__57_;
      r_133__56_ <= r_n_133__56_;
      r_133__55_ <= r_n_133__55_;
      r_133__54_ <= r_n_133__54_;
      r_133__53_ <= r_n_133__53_;
      r_133__52_ <= r_n_133__52_;
      r_133__51_ <= r_n_133__51_;
      r_133__50_ <= r_n_133__50_;
      r_133__49_ <= r_n_133__49_;
      r_133__48_ <= r_n_133__48_;
      r_133__47_ <= r_n_133__47_;
      r_133__46_ <= r_n_133__46_;
      r_133__45_ <= r_n_133__45_;
      r_133__44_ <= r_n_133__44_;
      r_133__43_ <= r_n_133__43_;
      r_133__42_ <= r_n_133__42_;
      r_133__41_ <= r_n_133__41_;
      r_133__40_ <= r_n_133__40_;
      r_133__39_ <= r_n_133__39_;
      r_133__38_ <= r_n_133__38_;
      r_133__37_ <= r_n_133__37_;
      r_133__36_ <= r_n_133__36_;
      r_133__35_ <= r_n_133__35_;
      r_133__34_ <= r_n_133__34_;
      r_133__33_ <= r_n_133__33_;
      r_133__32_ <= r_n_133__32_;
      r_133__31_ <= r_n_133__31_;
      r_133__30_ <= r_n_133__30_;
      r_133__29_ <= r_n_133__29_;
      r_133__28_ <= r_n_133__28_;
      r_133__27_ <= r_n_133__27_;
      r_133__26_ <= r_n_133__26_;
      r_133__25_ <= r_n_133__25_;
      r_133__24_ <= r_n_133__24_;
      r_133__23_ <= r_n_133__23_;
      r_133__22_ <= r_n_133__22_;
      r_133__21_ <= r_n_133__21_;
      r_133__20_ <= r_n_133__20_;
      r_133__19_ <= r_n_133__19_;
      r_133__18_ <= r_n_133__18_;
      r_133__17_ <= r_n_133__17_;
      r_133__16_ <= r_n_133__16_;
      r_133__15_ <= r_n_133__15_;
      r_133__14_ <= r_n_133__14_;
      r_133__13_ <= r_n_133__13_;
      r_133__12_ <= r_n_133__12_;
      r_133__11_ <= r_n_133__11_;
      r_133__10_ <= r_n_133__10_;
      r_133__9_ <= r_n_133__9_;
      r_133__8_ <= r_n_133__8_;
      r_133__7_ <= r_n_133__7_;
      r_133__6_ <= r_n_133__6_;
      r_133__5_ <= r_n_133__5_;
      r_133__4_ <= r_n_133__4_;
      r_133__3_ <= r_n_133__3_;
      r_133__2_ <= r_n_133__2_;
      r_133__1_ <= r_n_133__1_;
      r_133__0_ <= r_n_133__0_;
    end 
    if(N3718) begin
      r_134__63_ <= r_n_134__63_;
      r_134__62_ <= r_n_134__62_;
      r_134__61_ <= r_n_134__61_;
      r_134__60_ <= r_n_134__60_;
      r_134__59_ <= r_n_134__59_;
      r_134__58_ <= r_n_134__58_;
      r_134__57_ <= r_n_134__57_;
      r_134__56_ <= r_n_134__56_;
      r_134__55_ <= r_n_134__55_;
      r_134__54_ <= r_n_134__54_;
      r_134__53_ <= r_n_134__53_;
      r_134__52_ <= r_n_134__52_;
      r_134__51_ <= r_n_134__51_;
      r_134__50_ <= r_n_134__50_;
      r_134__49_ <= r_n_134__49_;
      r_134__48_ <= r_n_134__48_;
      r_134__47_ <= r_n_134__47_;
      r_134__46_ <= r_n_134__46_;
      r_134__45_ <= r_n_134__45_;
      r_134__44_ <= r_n_134__44_;
      r_134__43_ <= r_n_134__43_;
      r_134__42_ <= r_n_134__42_;
      r_134__41_ <= r_n_134__41_;
      r_134__40_ <= r_n_134__40_;
      r_134__39_ <= r_n_134__39_;
      r_134__38_ <= r_n_134__38_;
      r_134__37_ <= r_n_134__37_;
      r_134__36_ <= r_n_134__36_;
      r_134__35_ <= r_n_134__35_;
      r_134__34_ <= r_n_134__34_;
      r_134__33_ <= r_n_134__33_;
      r_134__32_ <= r_n_134__32_;
      r_134__31_ <= r_n_134__31_;
      r_134__30_ <= r_n_134__30_;
      r_134__29_ <= r_n_134__29_;
      r_134__28_ <= r_n_134__28_;
      r_134__27_ <= r_n_134__27_;
      r_134__26_ <= r_n_134__26_;
      r_134__25_ <= r_n_134__25_;
      r_134__24_ <= r_n_134__24_;
      r_134__23_ <= r_n_134__23_;
      r_134__22_ <= r_n_134__22_;
      r_134__21_ <= r_n_134__21_;
      r_134__20_ <= r_n_134__20_;
      r_134__19_ <= r_n_134__19_;
      r_134__18_ <= r_n_134__18_;
      r_134__17_ <= r_n_134__17_;
      r_134__16_ <= r_n_134__16_;
      r_134__15_ <= r_n_134__15_;
      r_134__14_ <= r_n_134__14_;
      r_134__13_ <= r_n_134__13_;
      r_134__12_ <= r_n_134__12_;
      r_134__11_ <= r_n_134__11_;
      r_134__10_ <= r_n_134__10_;
      r_134__9_ <= r_n_134__9_;
      r_134__8_ <= r_n_134__8_;
      r_134__7_ <= r_n_134__7_;
      r_134__6_ <= r_n_134__6_;
      r_134__5_ <= r_n_134__5_;
      r_134__4_ <= r_n_134__4_;
      r_134__3_ <= r_n_134__3_;
      r_134__2_ <= r_n_134__2_;
      r_134__1_ <= r_n_134__1_;
      r_134__0_ <= r_n_134__0_;
    end 
    if(N3719) begin
      r_135__63_ <= r_n_135__63_;
      r_135__62_ <= r_n_135__62_;
      r_135__61_ <= r_n_135__61_;
      r_135__60_ <= r_n_135__60_;
      r_135__59_ <= r_n_135__59_;
      r_135__58_ <= r_n_135__58_;
      r_135__57_ <= r_n_135__57_;
      r_135__56_ <= r_n_135__56_;
      r_135__55_ <= r_n_135__55_;
      r_135__54_ <= r_n_135__54_;
      r_135__53_ <= r_n_135__53_;
      r_135__52_ <= r_n_135__52_;
      r_135__51_ <= r_n_135__51_;
      r_135__50_ <= r_n_135__50_;
      r_135__49_ <= r_n_135__49_;
      r_135__48_ <= r_n_135__48_;
      r_135__47_ <= r_n_135__47_;
      r_135__46_ <= r_n_135__46_;
      r_135__45_ <= r_n_135__45_;
      r_135__44_ <= r_n_135__44_;
      r_135__43_ <= r_n_135__43_;
      r_135__42_ <= r_n_135__42_;
      r_135__41_ <= r_n_135__41_;
      r_135__40_ <= r_n_135__40_;
      r_135__39_ <= r_n_135__39_;
      r_135__38_ <= r_n_135__38_;
      r_135__37_ <= r_n_135__37_;
      r_135__36_ <= r_n_135__36_;
      r_135__35_ <= r_n_135__35_;
      r_135__34_ <= r_n_135__34_;
      r_135__33_ <= r_n_135__33_;
      r_135__32_ <= r_n_135__32_;
      r_135__31_ <= r_n_135__31_;
      r_135__30_ <= r_n_135__30_;
      r_135__29_ <= r_n_135__29_;
      r_135__28_ <= r_n_135__28_;
      r_135__27_ <= r_n_135__27_;
      r_135__26_ <= r_n_135__26_;
      r_135__25_ <= r_n_135__25_;
      r_135__24_ <= r_n_135__24_;
      r_135__23_ <= r_n_135__23_;
      r_135__22_ <= r_n_135__22_;
      r_135__21_ <= r_n_135__21_;
      r_135__20_ <= r_n_135__20_;
      r_135__19_ <= r_n_135__19_;
      r_135__18_ <= r_n_135__18_;
      r_135__17_ <= r_n_135__17_;
      r_135__16_ <= r_n_135__16_;
      r_135__15_ <= r_n_135__15_;
      r_135__14_ <= r_n_135__14_;
      r_135__13_ <= r_n_135__13_;
      r_135__12_ <= r_n_135__12_;
      r_135__11_ <= r_n_135__11_;
      r_135__10_ <= r_n_135__10_;
      r_135__9_ <= r_n_135__9_;
      r_135__8_ <= r_n_135__8_;
      r_135__7_ <= r_n_135__7_;
      r_135__6_ <= r_n_135__6_;
      r_135__5_ <= r_n_135__5_;
      r_135__4_ <= r_n_135__4_;
      r_135__3_ <= r_n_135__3_;
      r_135__2_ <= r_n_135__2_;
      r_135__1_ <= r_n_135__1_;
      r_135__0_ <= r_n_135__0_;
    end 
    if(N3720) begin
      r_136__63_ <= r_n_136__63_;
      r_136__62_ <= r_n_136__62_;
      r_136__61_ <= r_n_136__61_;
      r_136__60_ <= r_n_136__60_;
      r_136__59_ <= r_n_136__59_;
      r_136__58_ <= r_n_136__58_;
      r_136__57_ <= r_n_136__57_;
      r_136__56_ <= r_n_136__56_;
      r_136__55_ <= r_n_136__55_;
      r_136__54_ <= r_n_136__54_;
      r_136__53_ <= r_n_136__53_;
      r_136__52_ <= r_n_136__52_;
      r_136__51_ <= r_n_136__51_;
      r_136__50_ <= r_n_136__50_;
      r_136__49_ <= r_n_136__49_;
      r_136__48_ <= r_n_136__48_;
      r_136__47_ <= r_n_136__47_;
      r_136__46_ <= r_n_136__46_;
      r_136__45_ <= r_n_136__45_;
      r_136__44_ <= r_n_136__44_;
      r_136__43_ <= r_n_136__43_;
      r_136__42_ <= r_n_136__42_;
      r_136__41_ <= r_n_136__41_;
      r_136__40_ <= r_n_136__40_;
      r_136__39_ <= r_n_136__39_;
      r_136__38_ <= r_n_136__38_;
      r_136__37_ <= r_n_136__37_;
      r_136__36_ <= r_n_136__36_;
      r_136__35_ <= r_n_136__35_;
      r_136__34_ <= r_n_136__34_;
      r_136__33_ <= r_n_136__33_;
      r_136__32_ <= r_n_136__32_;
      r_136__31_ <= r_n_136__31_;
      r_136__30_ <= r_n_136__30_;
      r_136__29_ <= r_n_136__29_;
      r_136__28_ <= r_n_136__28_;
      r_136__27_ <= r_n_136__27_;
      r_136__26_ <= r_n_136__26_;
      r_136__25_ <= r_n_136__25_;
      r_136__24_ <= r_n_136__24_;
      r_136__23_ <= r_n_136__23_;
      r_136__22_ <= r_n_136__22_;
      r_136__21_ <= r_n_136__21_;
      r_136__20_ <= r_n_136__20_;
      r_136__19_ <= r_n_136__19_;
      r_136__18_ <= r_n_136__18_;
      r_136__17_ <= r_n_136__17_;
      r_136__16_ <= r_n_136__16_;
      r_136__15_ <= r_n_136__15_;
      r_136__14_ <= r_n_136__14_;
      r_136__13_ <= r_n_136__13_;
      r_136__12_ <= r_n_136__12_;
      r_136__11_ <= r_n_136__11_;
      r_136__10_ <= r_n_136__10_;
      r_136__9_ <= r_n_136__9_;
      r_136__8_ <= r_n_136__8_;
      r_136__7_ <= r_n_136__7_;
      r_136__6_ <= r_n_136__6_;
      r_136__5_ <= r_n_136__5_;
      r_136__4_ <= r_n_136__4_;
      r_136__3_ <= r_n_136__3_;
      r_136__2_ <= r_n_136__2_;
      r_136__1_ <= r_n_136__1_;
      r_136__0_ <= r_n_136__0_;
    end 
    if(N3721) begin
      r_137__63_ <= r_n_137__63_;
      r_137__62_ <= r_n_137__62_;
      r_137__61_ <= r_n_137__61_;
      r_137__60_ <= r_n_137__60_;
      r_137__59_ <= r_n_137__59_;
      r_137__58_ <= r_n_137__58_;
      r_137__57_ <= r_n_137__57_;
      r_137__56_ <= r_n_137__56_;
      r_137__55_ <= r_n_137__55_;
      r_137__54_ <= r_n_137__54_;
      r_137__53_ <= r_n_137__53_;
      r_137__52_ <= r_n_137__52_;
      r_137__51_ <= r_n_137__51_;
      r_137__50_ <= r_n_137__50_;
      r_137__49_ <= r_n_137__49_;
      r_137__48_ <= r_n_137__48_;
      r_137__47_ <= r_n_137__47_;
      r_137__46_ <= r_n_137__46_;
      r_137__45_ <= r_n_137__45_;
      r_137__44_ <= r_n_137__44_;
      r_137__43_ <= r_n_137__43_;
      r_137__42_ <= r_n_137__42_;
      r_137__41_ <= r_n_137__41_;
      r_137__40_ <= r_n_137__40_;
      r_137__39_ <= r_n_137__39_;
      r_137__38_ <= r_n_137__38_;
      r_137__37_ <= r_n_137__37_;
      r_137__36_ <= r_n_137__36_;
      r_137__35_ <= r_n_137__35_;
      r_137__34_ <= r_n_137__34_;
      r_137__33_ <= r_n_137__33_;
      r_137__32_ <= r_n_137__32_;
      r_137__31_ <= r_n_137__31_;
      r_137__30_ <= r_n_137__30_;
      r_137__29_ <= r_n_137__29_;
      r_137__28_ <= r_n_137__28_;
      r_137__27_ <= r_n_137__27_;
      r_137__26_ <= r_n_137__26_;
      r_137__25_ <= r_n_137__25_;
      r_137__24_ <= r_n_137__24_;
      r_137__23_ <= r_n_137__23_;
      r_137__22_ <= r_n_137__22_;
      r_137__21_ <= r_n_137__21_;
      r_137__20_ <= r_n_137__20_;
      r_137__19_ <= r_n_137__19_;
      r_137__18_ <= r_n_137__18_;
      r_137__17_ <= r_n_137__17_;
      r_137__16_ <= r_n_137__16_;
      r_137__15_ <= r_n_137__15_;
      r_137__14_ <= r_n_137__14_;
      r_137__13_ <= r_n_137__13_;
      r_137__12_ <= r_n_137__12_;
      r_137__11_ <= r_n_137__11_;
      r_137__10_ <= r_n_137__10_;
      r_137__9_ <= r_n_137__9_;
      r_137__8_ <= r_n_137__8_;
      r_137__7_ <= r_n_137__7_;
      r_137__6_ <= r_n_137__6_;
      r_137__5_ <= r_n_137__5_;
      r_137__4_ <= r_n_137__4_;
      r_137__3_ <= r_n_137__3_;
      r_137__2_ <= r_n_137__2_;
      r_137__1_ <= r_n_137__1_;
      r_137__0_ <= r_n_137__0_;
    end 
    if(N3722) begin
      r_138__63_ <= r_n_138__63_;
      r_138__62_ <= r_n_138__62_;
      r_138__61_ <= r_n_138__61_;
      r_138__60_ <= r_n_138__60_;
      r_138__59_ <= r_n_138__59_;
      r_138__58_ <= r_n_138__58_;
      r_138__57_ <= r_n_138__57_;
      r_138__56_ <= r_n_138__56_;
      r_138__55_ <= r_n_138__55_;
      r_138__54_ <= r_n_138__54_;
      r_138__53_ <= r_n_138__53_;
      r_138__52_ <= r_n_138__52_;
      r_138__51_ <= r_n_138__51_;
      r_138__50_ <= r_n_138__50_;
      r_138__49_ <= r_n_138__49_;
      r_138__48_ <= r_n_138__48_;
      r_138__47_ <= r_n_138__47_;
      r_138__46_ <= r_n_138__46_;
      r_138__45_ <= r_n_138__45_;
      r_138__44_ <= r_n_138__44_;
      r_138__43_ <= r_n_138__43_;
      r_138__42_ <= r_n_138__42_;
      r_138__41_ <= r_n_138__41_;
      r_138__40_ <= r_n_138__40_;
      r_138__39_ <= r_n_138__39_;
      r_138__38_ <= r_n_138__38_;
      r_138__37_ <= r_n_138__37_;
      r_138__36_ <= r_n_138__36_;
      r_138__35_ <= r_n_138__35_;
      r_138__34_ <= r_n_138__34_;
      r_138__33_ <= r_n_138__33_;
      r_138__32_ <= r_n_138__32_;
      r_138__31_ <= r_n_138__31_;
      r_138__30_ <= r_n_138__30_;
      r_138__29_ <= r_n_138__29_;
      r_138__28_ <= r_n_138__28_;
      r_138__27_ <= r_n_138__27_;
      r_138__26_ <= r_n_138__26_;
      r_138__25_ <= r_n_138__25_;
      r_138__24_ <= r_n_138__24_;
      r_138__23_ <= r_n_138__23_;
      r_138__22_ <= r_n_138__22_;
      r_138__21_ <= r_n_138__21_;
      r_138__20_ <= r_n_138__20_;
      r_138__19_ <= r_n_138__19_;
      r_138__18_ <= r_n_138__18_;
      r_138__17_ <= r_n_138__17_;
      r_138__16_ <= r_n_138__16_;
      r_138__15_ <= r_n_138__15_;
      r_138__14_ <= r_n_138__14_;
      r_138__13_ <= r_n_138__13_;
      r_138__12_ <= r_n_138__12_;
      r_138__11_ <= r_n_138__11_;
      r_138__10_ <= r_n_138__10_;
      r_138__9_ <= r_n_138__9_;
      r_138__8_ <= r_n_138__8_;
      r_138__7_ <= r_n_138__7_;
      r_138__6_ <= r_n_138__6_;
      r_138__5_ <= r_n_138__5_;
      r_138__4_ <= r_n_138__4_;
      r_138__3_ <= r_n_138__3_;
      r_138__2_ <= r_n_138__2_;
      r_138__1_ <= r_n_138__1_;
      r_138__0_ <= r_n_138__0_;
    end 
    if(N3723) begin
      r_139__63_ <= r_n_139__63_;
      r_139__62_ <= r_n_139__62_;
      r_139__61_ <= r_n_139__61_;
      r_139__60_ <= r_n_139__60_;
      r_139__59_ <= r_n_139__59_;
      r_139__58_ <= r_n_139__58_;
      r_139__57_ <= r_n_139__57_;
      r_139__56_ <= r_n_139__56_;
      r_139__55_ <= r_n_139__55_;
      r_139__54_ <= r_n_139__54_;
      r_139__53_ <= r_n_139__53_;
      r_139__52_ <= r_n_139__52_;
      r_139__51_ <= r_n_139__51_;
      r_139__50_ <= r_n_139__50_;
      r_139__49_ <= r_n_139__49_;
      r_139__48_ <= r_n_139__48_;
      r_139__47_ <= r_n_139__47_;
      r_139__46_ <= r_n_139__46_;
      r_139__45_ <= r_n_139__45_;
      r_139__44_ <= r_n_139__44_;
      r_139__43_ <= r_n_139__43_;
      r_139__42_ <= r_n_139__42_;
      r_139__41_ <= r_n_139__41_;
      r_139__40_ <= r_n_139__40_;
      r_139__39_ <= r_n_139__39_;
      r_139__38_ <= r_n_139__38_;
      r_139__37_ <= r_n_139__37_;
      r_139__36_ <= r_n_139__36_;
      r_139__35_ <= r_n_139__35_;
      r_139__34_ <= r_n_139__34_;
      r_139__33_ <= r_n_139__33_;
      r_139__32_ <= r_n_139__32_;
      r_139__31_ <= r_n_139__31_;
      r_139__30_ <= r_n_139__30_;
      r_139__29_ <= r_n_139__29_;
      r_139__28_ <= r_n_139__28_;
      r_139__27_ <= r_n_139__27_;
      r_139__26_ <= r_n_139__26_;
      r_139__25_ <= r_n_139__25_;
      r_139__24_ <= r_n_139__24_;
      r_139__23_ <= r_n_139__23_;
      r_139__22_ <= r_n_139__22_;
      r_139__21_ <= r_n_139__21_;
      r_139__20_ <= r_n_139__20_;
      r_139__19_ <= r_n_139__19_;
      r_139__18_ <= r_n_139__18_;
      r_139__17_ <= r_n_139__17_;
      r_139__16_ <= r_n_139__16_;
      r_139__15_ <= r_n_139__15_;
      r_139__14_ <= r_n_139__14_;
      r_139__13_ <= r_n_139__13_;
      r_139__12_ <= r_n_139__12_;
      r_139__11_ <= r_n_139__11_;
      r_139__10_ <= r_n_139__10_;
      r_139__9_ <= r_n_139__9_;
      r_139__8_ <= r_n_139__8_;
      r_139__7_ <= r_n_139__7_;
      r_139__6_ <= r_n_139__6_;
      r_139__5_ <= r_n_139__5_;
      r_139__4_ <= r_n_139__4_;
      r_139__3_ <= r_n_139__3_;
      r_139__2_ <= r_n_139__2_;
      r_139__1_ <= r_n_139__1_;
      r_139__0_ <= r_n_139__0_;
    end 
    if(N3724) begin
      r_140__63_ <= r_n_140__63_;
      r_140__62_ <= r_n_140__62_;
      r_140__61_ <= r_n_140__61_;
      r_140__60_ <= r_n_140__60_;
      r_140__59_ <= r_n_140__59_;
      r_140__58_ <= r_n_140__58_;
      r_140__57_ <= r_n_140__57_;
      r_140__56_ <= r_n_140__56_;
      r_140__55_ <= r_n_140__55_;
      r_140__54_ <= r_n_140__54_;
      r_140__53_ <= r_n_140__53_;
      r_140__52_ <= r_n_140__52_;
      r_140__51_ <= r_n_140__51_;
      r_140__50_ <= r_n_140__50_;
      r_140__49_ <= r_n_140__49_;
      r_140__48_ <= r_n_140__48_;
      r_140__47_ <= r_n_140__47_;
      r_140__46_ <= r_n_140__46_;
      r_140__45_ <= r_n_140__45_;
      r_140__44_ <= r_n_140__44_;
      r_140__43_ <= r_n_140__43_;
      r_140__42_ <= r_n_140__42_;
      r_140__41_ <= r_n_140__41_;
      r_140__40_ <= r_n_140__40_;
      r_140__39_ <= r_n_140__39_;
      r_140__38_ <= r_n_140__38_;
      r_140__37_ <= r_n_140__37_;
      r_140__36_ <= r_n_140__36_;
      r_140__35_ <= r_n_140__35_;
      r_140__34_ <= r_n_140__34_;
      r_140__33_ <= r_n_140__33_;
      r_140__32_ <= r_n_140__32_;
      r_140__31_ <= r_n_140__31_;
      r_140__30_ <= r_n_140__30_;
      r_140__29_ <= r_n_140__29_;
      r_140__28_ <= r_n_140__28_;
      r_140__27_ <= r_n_140__27_;
      r_140__26_ <= r_n_140__26_;
      r_140__25_ <= r_n_140__25_;
      r_140__24_ <= r_n_140__24_;
      r_140__23_ <= r_n_140__23_;
      r_140__22_ <= r_n_140__22_;
      r_140__21_ <= r_n_140__21_;
      r_140__20_ <= r_n_140__20_;
      r_140__19_ <= r_n_140__19_;
      r_140__18_ <= r_n_140__18_;
      r_140__17_ <= r_n_140__17_;
      r_140__16_ <= r_n_140__16_;
      r_140__15_ <= r_n_140__15_;
      r_140__14_ <= r_n_140__14_;
      r_140__13_ <= r_n_140__13_;
      r_140__12_ <= r_n_140__12_;
      r_140__11_ <= r_n_140__11_;
      r_140__10_ <= r_n_140__10_;
      r_140__9_ <= r_n_140__9_;
      r_140__8_ <= r_n_140__8_;
      r_140__7_ <= r_n_140__7_;
      r_140__6_ <= r_n_140__6_;
      r_140__5_ <= r_n_140__5_;
      r_140__4_ <= r_n_140__4_;
      r_140__3_ <= r_n_140__3_;
      r_140__2_ <= r_n_140__2_;
      r_140__1_ <= r_n_140__1_;
      r_140__0_ <= r_n_140__0_;
    end 
    if(N3725) begin
      r_141__63_ <= r_n_141__63_;
      r_141__62_ <= r_n_141__62_;
      r_141__61_ <= r_n_141__61_;
      r_141__60_ <= r_n_141__60_;
      r_141__59_ <= r_n_141__59_;
      r_141__58_ <= r_n_141__58_;
      r_141__57_ <= r_n_141__57_;
      r_141__56_ <= r_n_141__56_;
      r_141__55_ <= r_n_141__55_;
      r_141__54_ <= r_n_141__54_;
      r_141__53_ <= r_n_141__53_;
      r_141__52_ <= r_n_141__52_;
      r_141__51_ <= r_n_141__51_;
      r_141__50_ <= r_n_141__50_;
      r_141__49_ <= r_n_141__49_;
      r_141__48_ <= r_n_141__48_;
      r_141__47_ <= r_n_141__47_;
      r_141__46_ <= r_n_141__46_;
      r_141__45_ <= r_n_141__45_;
      r_141__44_ <= r_n_141__44_;
      r_141__43_ <= r_n_141__43_;
      r_141__42_ <= r_n_141__42_;
      r_141__41_ <= r_n_141__41_;
      r_141__40_ <= r_n_141__40_;
      r_141__39_ <= r_n_141__39_;
      r_141__38_ <= r_n_141__38_;
      r_141__37_ <= r_n_141__37_;
      r_141__36_ <= r_n_141__36_;
      r_141__35_ <= r_n_141__35_;
      r_141__34_ <= r_n_141__34_;
      r_141__33_ <= r_n_141__33_;
      r_141__32_ <= r_n_141__32_;
      r_141__31_ <= r_n_141__31_;
      r_141__30_ <= r_n_141__30_;
      r_141__29_ <= r_n_141__29_;
      r_141__28_ <= r_n_141__28_;
      r_141__27_ <= r_n_141__27_;
      r_141__26_ <= r_n_141__26_;
      r_141__25_ <= r_n_141__25_;
      r_141__24_ <= r_n_141__24_;
      r_141__23_ <= r_n_141__23_;
      r_141__22_ <= r_n_141__22_;
      r_141__21_ <= r_n_141__21_;
      r_141__20_ <= r_n_141__20_;
      r_141__19_ <= r_n_141__19_;
      r_141__18_ <= r_n_141__18_;
      r_141__17_ <= r_n_141__17_;
      r_141__16_ <= r_n_141__16_;
      r_141__15_ <= r_n_141__15_;
      r_141__14_ <= r_n_141__14_;
      r_141__13_ <= r_n_141__13_;
      r_141__12_ <= r_n_141__12_;
      r_141__11_ <= r_n_141__11_;
      r_141__10_ <= r_n_141__10_;
      r_141__9_ <= r_n_141__9_;
      r_141__8_ <= r_n_141__8_;
      r_141__7_ <= r_n_141__7_;
      r_141__6_ <= r_n_141__6_;
      r_141__5_ <= r_n_141__5_;
      r_141__4_ <= r_n_141__4_;
      r_141__3_ <= r_n_141__3_;
      r_141__2_ <= r_n_141__2_;
      r_141__1_ <= r_n_141__1_;
      r_141__0_ <= r_n_141__0_;
    end 
    if(N3726) begin
      r_142__63_ <= r_n_142__63_;
      r_142__62_ <= r_n_142__62_;
      r_142__61_ <= r_n_142__61_;
      r_142__60_ <= r_n_142__60_;
      r_142__59_ <= r_n_142__59_;
      r_142__58_ <= r_n_142__58_;
      r_142__57_ <= r_n_142__57_;
      r_142__56_ <= r_n_142__56_;
      r_142__55_ <= r_n_142__55_;
      r_142__54_ <= r_n_142__54_;
      r_142__53_ <= r_n_142__53_;
      r_142__52_ <= r_n_142__52_;
      r_142__51_ <= r_n_142__51_;
      r_142__50_ <= r_n_142__50_;
      r_142__49_ <= r_n_142__49_;
      r_142__48_ <= r_n_142__48_;
      r_142__47_ <= r_n_142__47_;
      r_142__46_ <= r_n_142__46_;
      r_142__45_ <= r_n_142__45_;
      r_142__44_ <= r_n_142__44_;
      r_142__43_ <= r_n_142__43_;
      r_142__42_ <= r_n_142__42_;
      r_142__41_ <= r_n_142__41_;
      r_142__40_ <= r_n_142__40_;
      r_142__39_ <= r_n_142__39_;
      r_142__38_ <= r_n_142__38_;
      r_142__37_ <= r_n_142__37_;
      r_142__36_ <= r_n_142__36_;
      r_142__35_ <= r_n_142__35_;
      r_142__34_ <= r_n_142__34_;
      r_142__33_ <= r_n_142__33_;
      r_142__32_ <= r_n_142__32_;
      r_142__31_ <= r_n_142__31_;
      r_142__30_ <= r_n_142__30_;
      r_142__29_ <= r_n_142__29_;
      r_142__28_ <= r_n_142__28_;
      r_142__27_ <= r_n_142__27_;
      r_142__26_ <= r_n_142__26_;
      r_142__25_ <= r_n_142__25_;
      r_142__24_ <= r_n_142__24_;
      r_142__23_ <= r_n_142__23_;
      r_142__22_ <= r_n_142__22_;
      r_142__21_ <= r_n_142__21_;
      r_142__20_ <= r_n_142__20_;
      r_142__19_ <= r_n_142__19_;
      r_142__18_ <= r_n_142__18_;
      r_142__17_ <= r_n_142__17_;
      r_142__16_ <= r_n_142__16_;
      r_142__15_ <= r_n_142__15_;
      r_142__14_ <= r_n_142__14_;
      r_142__13_ <= r_n_142__13_;
      r_142__12_ <= r_n_142__12_;
      r_142__11_ <= r_n_142__11_;
      r_142__10_ <= r_n_142__10_;
      r_142__9_ <= r_n_142__9_;
      r_142__8_ <= r_n_142__8_;
      r_142__7_ <= r_n_142__7_;
      r_142__6_ <= r_n_142__6_;
      r_142__5_ <= r_n_142__5_;
      r_142__4_ <= r_n_142__4_;
      r_142__3_ <= r_n_142__3_;
      r_142__2_ <= r_n_142__2_;
      r_142__1_ <= r_n_142__1_;
      r_142__0_ <= r_n_142__0_;
    end 
    if(N3727) begin
      r_143__63_ <= r_n_143__63_;
      r_143__62_ <= r_n_143__62_;
      r_143__61_ <= r_n_143__61_;
      r_143__60_ <= r_n_143__60_;
      r_143__59_ <= r_n_143__59_;
      r_143__58_ <= r_n_143__58_;
      r_143__57_ <= r_n_143__57_;
      r_143__56_ <= r_n_143__56_;
      r_143__55_ <= r_n_143__55_;
      r_143__54_ <= r_n_143__54_;
      r_143__53_ <= r_n_143__53_;
      r_143__52_ <= r_n_143__52_;
      r_143__51_ <= r_n_143__51_;
      r_143__50_ <= r_n_143__50_;
      r_143__49_ <= r_n_143__49_;
      r_143__48_ <= r_n_143__48_;
      r_143__47_ <= r_n_143__47_;
      r_143__46_ <= r_n_143__46_;
      r_143__45_ <= r_n_143__45_;
      r_143__44_ <= r_n_143__44_;
      r_143__43_ <= r_n_143__43_;
      r_143__42_ <= r_n_143__42_;
      r_143__41_ <= r_n_143__41_;
      r_143__40_ <= r_n_143__40_;
      r_143__39_ <= r_n_143__39_;
      r_143__38_ <= r_n_143__38_;
      r_143__37_ <= r_n_143__37_;
      r_143__36_ <= r_n_143__36_;
      r_143__35_ <= r_n_143__35_;
      r_143__34_ <= r_n_143__34_;
      r_143__33_ <= r_n_143__33_;
      r_143__32_ <= r_n_143__32_;
      r_143__31_ <= r_n_143__31_;
      r_143__30_ <= r_n_143__30_;
      r_143__29_ <= r_n_143__29_;
      r_143__28_ <= r_n_143__28_;
      r_143__27_ <= r_n_143__27_;
      r_143__26_ <= r_n_143__26_;
      r_143__25_ <= r_n_143__25_;
      r_143__24_ <= r_n_143__24_;
      r_143__23_ <= r_n_143__23_;
      r_143__22_ <= r_n_143__22_;
      r_143__21_ <= r_n_143__21_;
      r_143__20_ <= r_n_143__20_;
      r_143__19_ <= r_n_143__19_;
      r_143__18_ <= r_n_143__18_;
      r_143__17_ <= r_n_143__17_;
      r_143__16_ <= r_n_143__16_;
      r_143__15_ <= r_n_143__15_;
      r_143__14_ <= r_n_143__14_;
      r_143__13_ <= r_n_143__13_;
      r_143__12_ <= r_n_143__12_;
      r_143__11_ <= r_n_143__11_;
      r_143__10_ <= r_n_143__10_;
      r_143__9_ <= r_n_143__9_;
      r_143__8_ <= r_n_143__8_;
      r_143__7_ <= r_n_143__7_;
      r_143__6_ <= r_n_143__6_;
      r_143__5_ <= r_n_143__5_;
      r_143__4_ <= r_n_143__4_;
      r_143__3_ <= r_n_143__3_;
      r_143__2_ <= r_n_143__2_;
      r_143__1_ <= r_n_143__1_;
      r_143__0_ <= r_n_143__0_;
    end 
    if(N3728) begin
      r_144__63_ <= r_n_144__63_;
      r_144__62_ <= r_n_144__62_;
      r_144__61_ <= r_n_144__61_;
      r_144__60_ <= r_n_144__60_;
      r_144__59_ <= r_n_144__59_;
      r_144__58_ <= r_n_144__58_;
      r_144__57_ <= r_n_144__57_;
      r_144__56_ <= r_n_144__56_;
      r_144__55_ <= r_n_144__55_;
      r_144__54_ <= r_n_144__54_;
      r_144__53_ <= r_n_144__53_;
      r_144__52_ <= r_n_144__52_;
      r_144__51_ <= r_n_144__51_;
      r_144__50_ <= r_n_144__50_;
      r_144__49_ <= r_n_144__49_;
      r_144__48_ <= r_n_144__48_;
      r_144__47_ <= r_n_144__47_;
      r_144__46_ <= r_n_144__46_;
      r_144__45_ <= r_n_144__45_;
      r_144__44_ <= r_n_144__44_;
      r_144__43_ <= r_n_144__43_;
      r_144__42_ <= r_n_144__42_;
      r_144__41_ <= r_n_144__41_;
      r_144__40_ <= r_n_144__40_;
      r_144__39_ <= r_n_144__39_;
      r_144__38_ <= r_n_144__38_;
      r_144__37_ <= r_n_144__37_;
      r_144__36_ <= r_n_144__36_;
      r_144__35_ <= r_n_144__35_;
      r_144__34_ <= r_n_144__34_;
      r_144__33_ <= r_n_144__33_;
      r_144__32_ <= r_n_144__32_;
      r_144__31_ <= r_n_144__31_;
      r_144__30_ <= r_n_144__30_;
      r_144__29_ <= r_n_144__29_;
      r_144__28_ <= r_n_144__28_;
      r_144__27_ <= r_n_144__27_;
      r_144__26_ <= r_n_144__26_;
      r_144__25_ <= r_n_144__25_;
      r_144__24_ <= r_n_144__24_;
      r_144__23_ <= r_n_144__23_;
      r_144__22_ <= r_n_144__22_;
      r_144__21_ <= r_n_144__21_;
      r_144__20_ <= r_n_144__20_;
      r_144__19_ <= r_n_144__19_;
      r_144__18_ <= r_n_144__18_;
      r_144__17_ <= r_n_144__17_;
      r_144__16_ <= r_n_144__16_;
      r_144__15_ <= r_n_144__15_;
      r_144__14_ <= r_n_144__14_;
      r_144__13_ <= r_n_144__13_;
      r_144__12_ <= r_n_144__12_;
      r_144__11_ <= r_n_144__11_;
      r_144__10_ <= r_n_144__10_;
      r_144__9_ <= r_n_144__9_;
      r_144__8_ <= r_n_144__8_;
      r_144__7_ <= r_n_144__7_;
      r_144__6_ <= r_n_144__6_;
      r_144__5_ <= r_n_144__5_;
      r_144__4_ <= r_n_144__4_;
      r_144__3_ <= r_n_144__3_;
      r_144__2_ <= r_n_144__2_;
      r_144__1_ <= r_n_144__1_;
      r_144__0_ <= r_n_144__0_;
    end 
    if(N3729) begin
      r_145__63_ <= r_n_145__63_;
      r_145__62_ <= r_n_145__62_;
      r_145__61_ <= r_n_145__61_;
      r_145__60_ <= r_n_145__60_;
      r_145__59_ <= r_n_145__59_;
      r_145__58_ <= r_n_145__58_;
      r_145__57_ <= r_n_145__57_;
      r_145__56_ <= r_n_145__56_;
      r_145__55_ <= r_n_145__55_;
      r_145__54_ <= r_n_145__54_;
      r_145__53_ <= r_n_145__53_;
      r_145__52_ <= r_n_145__52_;
      r_145__51_ <= r_n_145__51_;
      r_145__50_ <= r_n_145__50_;
      r_145__49_ <= r_n_145__49_;
      r_145__48_ <= r_n_145__48_;
      r_145__47_ <= r_n_145__47_;
      r_145__46_ <= r_n_145__46_;
      r_145__45_ <= r_n_145__45_;
      r_145__44_ <= r_n_145__44_;
      r_145__43_ <= r_n_145__43_;
      r_145__42_ <= r_n_145__42_;
      r_145__41_ <= r_n_145__41_;
      r_145__40_ <= r_n_145__40_;
      r_145__39_ <= r_n_145__39_;
      r_145__38_ <= r_n_145__38_;
      r_145__37_ <= r_n_145__37_;
      r_145__36_ <= r_n_145__36_;
      r_145__35_ <= r_n_145__35_;
      r_145__34_ <= r_n_145__34_;
      r_145__33_ <= r_n_145__33_;
      r_145__32_ <= r_n_145__32_;
      r_145__31_ <= r_n_145__31_;
      r_145__30_ <= r_n_145__30_;
      r_145__29_ <= r_n_145__29_;
      r_145__28_ <= r_n_145__28_;
      r_145__27_ <= r_n_145__27_;
      r_145__26_ <= r_n_145__26_;
      r_145__25_ <= r_n_145__25_;
      r_145__24_ <= r_n_145__24_;
      r_145__23_ <= r_n_145__23_;
      r_145__22_ <= r_n_145__22_;
      r_145__21_ <= r_n_145__21_;
      r_145__20_ <= r_n_145__20_;
      r_145__19_ <= r_n_145__19_;
      r_145__18_ <= r_n_145__18_;
      r_145__17_ <= r_n_145__17_;
      r_145__16_ <= r_n_145__16_;
      r_145__15_ <= r_n_145__15_;
      r_145__14_ <= r_n_145__14_;
      r_145__13_ <= r_n_145__13_;
      r_145__12_ <= r_n_145__12_;
      r_145__11_ <= r_n_145__11_;
      r_145__10_ <= r_n_145__10_;
      r_145__9_ <= r_n_145__9_;
      r_145__8_ <= r_n_145__8_;
      r_145__7_ <= r_n_145__7_;
      r_145__6_ <= r_n_145__6_;
      r_145__5_ <= r_n_145__5_;
      r_145__4_ <= r_n_145__4_;
      r_145__3_ <= r_n_145__3_;
      r_145__2_ <= r_n_145__2_;
      r_145__1_ <= r_n_145__1_;
      r_145__0_ <= r_n_145__0_;
    end 
    if(N3730) begin
      r_146__63_ <= r_n_146__63_;
      r_146__62_ <= r_n_146__62_;
      r_146__61_ <= r_n_146__61_;
      r_146__60_ <= r_n_146__60_;
      r_146__59_ <= r_n_146__59_;
      r_146__58_ <= r_n_146__58_;
      r_146__57_ <= r_n_146__57_;
      r_146__56_ <= r_n_146__56_;
      r_146__55_ <= r_n_146__55_;
      r_146__54_ <= r_n_146__54_;
      r_146__53_ <= r_n_146__53_;
      r_146__52_ <= r_n_146__52_;
      r_146__51_ <= r_n_146__51_;
      r_146__50_ <= r_n_146__50_;
      r_146__49_ <= r_n_146__49_;
      r_146__48_ <= r_n_146__48_;
      r_146__47_ <= r_n_146__47_;
      r_146__46_ <= r_n_146__46_;
      r_146__45_ <= r_n_146__45_;
      r_146__44_ <= r_n_146__44_;
      r_146__43_ <= r_n_146__43_;
      r_146__42_ <= r_n_146__42_;
      r_146__41_ <= r_n_146__41_;
      r_146__40_ <= r_n_146__40_;
      r_146__39_ <= r_n_146__39_;
      r_146__38_ <= r_n_146__38_;
      r_146__37_ <= r_n_146__37_;
      r_146__36_ <= r_n_146__36_;
      r_146__35_ <= r_n_146__35_;
      r_146__34_ <= r_n_146__34_;
      r_146__33_ <= r_n_146__33_;
      r_146__32_ <= r_n_146__32_;
      r_146__31_ <= r_n_146__31_;
      r_146__30_ <= r_n_146__30_;
      r_146__29_ <= r_n_146__29_;
      r_146__28_ <= r_n_146__28_;
      r_146__27_ <= r_n_146__27_;
      r_146__26_ <= r_n_146__26_;
      r_146__25_ <= r_n_146__25_;
      r_146__24_ <= r_n_146__24_;
      r_146__23_ <= r_n_146__23_;
      r_146__22_ <= r_n_146__22_;
      r_146__21_ <= r_n_146__21_;
      r_146__20_ <= r_n_146__20_;
      r_146__19_ <= r_n_146__19_;
      r_146__18_ <= r_n_146__18_;
      r_146__17_ <= r_n_146__17_;
      r_146__16_ <= r_n_146__16_;
      r_146__15_ <= r_n_146__15_;
      r_146__14_ <= r_n_146__14_;
      r_146__13_ <= r_n_146__13_;
      r_146__12_ <= r_n_146__12_;
      r_146__11_ <= r_n_146__11_;
      r_146__10_ <= r_n_146__10_;
      r_146__9_ <= r_n_146__9_;
      r_146__8_ <= r_n_146__8_;
      r_146__7_ <= r_n_146__7_;
      r_146__6_ <= r_n_146__6_;
      r_146__5_ <= r_n_146__5_;
      r_146__4_ <= r_n_146__4_;
      r_146__3_ <= r_n_146__3_;
      r_146__2_ <= r_n_146__2_;
      r_146__1_ <= r_n_146__1_;
      r_146__0_ <= r_n_146__0_;
    end 
    if(N3731) begin
      r_147__63_ <= r_n_147__63_;
      r_147__62_ <= r_n_147__62_;
      r_147__61_ <= r_n_147__61_;
      r_147__60_ <= r_n_147__60_;
      r_147__59_ <= r_n_147__59_;
      r_147__58_ <= r_n_147__58_;
      r_147__57_ <= r_n_147__57_;
      r_147__56_ <= r_n_147__56_;
      r_147__55_ <= r_n_147__55_;
      r_147__54_ <= r_n_147__54_;
      r_147__53_ <= r_n_147__53_;
      r_147__52_ <= r_n_147__52_;
      r_147__51_ <= r_n_147__51_;
      r_147__50_ <= r_n_147__50_;
      r_147__49_ <= r_n_147__49_;
      r_147__48_ <= r_n_147__48_;
      r_147__47_ <= r_n_147__47_;
      r_147__46_ <= r_n_147__46_;
      r_147__45_ <= r_n_147__45_;
      r_147__44_ <= r_n_147__44_;
      r_147__43_ <= r_n_147__43_;
      r_147__42_ <= r_n_147__42_;
      r_147__41_ <= r_n_147__41_;
      r_147__40_ <= r_n_147__40_;
      r_147__39_ <= r_n_147__39_;
      r_147__38_ <= r_n_147__38_;
      r_147__37_ <= r_n_147__37_;
      r_147__36_ <= r_n_147__36_;
      r_147__35_ <= r_n_147__35_;
      r_147__34_ <= r_n_147__34_;
      r_147__33_ <= r_n_147__33_;
      r_147__32_ <= r_n_147__32_;
      r_147__31_ <= r_n_147__31_;
      r_147__30_ <= r_n_147__30_;
      r_147__29_ <= r_n_147__29_;
      r_147__28_ <= r_n_147__28_;
      r_147__27_ <= r_n_147__27_;
      r_147__26_ <= r_n_147__26_;
      r_147__25_ <= r_n_147__25_;
      r_147__24_ <= r_n_147__24_;
      r_147__23_ <= r_n_147__23_;
      r_147__22_ <= r_n_147__22_;
      r_147__21_ <= r_n_147__21_;
      r_147__20_ <= r_n_147__20_;
      r_147__19_ <= r_n_147__19_;
      r_147__18_ <= r_n_147__18_;
      r_147__17_ <= r_n_147__17_;
      r_147__16_ <= r_n_147__16_;
      r_147__15_ <= r_n_147__15_;
      r_147__14_ <= r_n_147__14_;
      r_147__13_ <= r_n_147__13_;
      r_147__12_ <= r_n_147__12_;
      r_147__11_ <= r_n_147__11_;
      r_147__10_ <= r_n_147__10_;
      r_147__9_ <= r_n_147__9_;
      r_147__8_ <= r_n_147__8_;
      r_147__7_ <= r_n_147__7_;
      r_147__6_ <= r_n_147__6_;
      r_147__5_ <= r_n_147__5_;
      r_147__4_ <= r_n_147__4_;
      r_147__3_ <= r_n_147__3_;
      r_147__2_ <= r_n_147__2_;
      r_147__1_ <= r_n_147__1_;
      r_147__0_ <= r_n_147__0_;
    end 
    if(N3732) begin
      r_148__63_ <= r_n_148__63_;
      r_148__62_ <= r_n_148__62_;
      r_148__61_ <= r_n_148__61_;
      r_148__60_ <= r_n_148__60_;
      r_148__59_ <= r_n_148__59_;
      r_148__58_ <= r_n_148__58_;
      r_148__57_ <= r_n_148__57_;
      r_148__56_ <= r_n_148__56_;
      r_148__55_ <= r_n_148__55_;
      r_148__54_ <= r_n_148__54_;
      r_148__53_ <= r_n_148__53_;
      r_148__52_ <= r_n_148__52_;
      r_148__51_ <= r_n_148__51_;
      r_148__50_ <= r_n_148__50_;
      r_148__49_ <= r_n_148__49_;
      r_148__48_ <= r_n_148__48_;
      r_148__47_ <= r_n_148__47_;
      r_148__46_ <= r_n_148__46_;
      r_148__45_ <= r_n_148__45_;
      r_148__44_ <= r_n_148__44_;
      r_148__43_ <= r_n_148__43_;
      r_148__42_ <= r_n_148__42_;
      r_148__41_ <= r_n_148__41_;
      r_148__40_ <= r_n_148__40_;
      r_148__39_ <= r_n_148__39_;
      r_148__38_ <= r_n_148__38_;
      r_148__37_ <= r_n_148__37_;
      r_148__36_ <= r_n_148__36_;
      r_148__35_ <= r_n_148__35_;
      r_148__34_ <= r_n_148__34_;
      r_148__33_ <= r_n_148__33_;
      r_148__32_ <= r_n_148__32_;
      r_148__31_ <= r_n_148__31_;
      r_148__30_ <= r_n_148__30_;
      r_148__29_ <= r_n_148__29_;
      r_148__28_ <= r_n_148__28_;
      r_148__27_ <= r_n_148__27_;
      r_148__26_ <= r_n_148__26_;
      r_148__25_ <= r_n_148__25_;
      r_148__24_ <= r_n_148__24_;
      r_148__23_ <= r_n_148__23_;
      r_148__22_ <= r_n_148__22_;
      r_148__21_ <= r_n_148__21_;
      r_148__20_ <= r_n_148__20_;
      r_148__19_ <= r_n_148__19_;
      r_148__18_ <= r_n_148__18_;
      r_148__17_ <= r_n_148__17_;
      r_148__16_ <= r_n_148__16_;
      r_148__15_ <= r_n_148__15_;
      r_148__14_ <= r_n_148__14_;
      r_148__13_ <= r_n_148__13_;
      r_148__12_ <= r_n_148__12_;
      r_148__11_ <= r_n_148__11_;
      r_148__10_ <= r_n_148__10_;
      r_148__9_ <= r_n_148__9_;
      r_148__8_ <= r_n_148__8_;
      r_148__7_ <= r_n_148__7_;
      r_148__6_ <= r_n_148__6_;
      r_148__5_ <= r_n_148__5_;
      r_148__4_ <= r_n_148__4_;
      r_148__3_ <= r_n_148__3_;
      r_148__2_ <= r_n_148__2_;
      r_148__1_ <= r_n_148__1_;
      r_148__0_ <= r_n_148__0_;
    end 
    if(N3733) begin
      r_149__63_ <= r_n_149__63_;
      r_149__62_ <= r_n_149__62_;
      r_149__61_ <= r_n_149__61_;
      r_149__60_ <= r_n_149__60_;
      r_149__59_ <= r_n_149__59_;
      r_149__58_ <= r_n_149__58_;
      r_149__57_ <= r_n_149__57_;
      r_149__56_ <= r_n_149__56_;
      r_149__55_ <= r_n_149__55_;
      r_149__54_ <= r_n_149__54_;
      r_149__53_ <= r_n_149__53_;
      r_149__52_ <= r_n_149__52_;
      r_149__51_ <= r_n_149__51_;
      r_149__50_ <= r_n_149__50_;
      r_149__49_ <= r_n_149__49_;
      r_149__48_ <= r_n_149__48_;
      r_149__47_ <= r_n_149__47_;
      r_149__46_ <= r_n_149__46_;
      r_149__45_ <= r_n_149__45_;
      r_149__44_ <= r_n_149__44_;
      r_149__43_ <= r_n_149__43_;
      r_149__42_ <= r_n_149__42_;
      r_149__41_ <= r_n_149__41_;
      r_149__40_ <= r_n_149__40_;
      r_149__39_ <= r_n_149__39_;
      r_149__38_ <= r_n_149__38_;
      r_149__37_ <= r_n_149__37_;
      r_149__36_ <= r_n_149__36_;
      r_149__35_ <= r_n_149__35_;
      r_149__34_ <= r_n_149__34_;
      r_149__33_ <= r_n_149__33_;
      r_149__32_ <= r_n_149__32_;
      r_149__31_ <= r_n_149__31_;
      r_149__30_ <= r_n_149__30_;
      r_149__29_ <= r_n_149__29_;
      r_149__28_ <= r_n_149__28_;
      r_149__27_ <= r_n_149__27_;
      r_149__26_ <= r_n_149__26_;
      r_149__25_ <= r_n_149__25_;
      r_149__24_ <= r_n_149__24_;
      r_149__23_ <= r_n_149__23_;
      r_149__22_ <= r_n_149__22_;
      r_149__21_ <= r_n_149__21_;
      r_149__20_ <= r_n_149__20_;
      r_149__19_ <= r_n_149__19_;
      r_149__18_ <= r_n_149__18_;
      r_149__17_ <= r_n_149__17_;
      r_149__16_ <= r_n_149__16_;
      r_149__15_ <= r_n_149__15_;
      r_149__14_ <= r_n_149__14_;
      r_149__13_ <= r_n_149__13_;
      r_149__12_ <= r_n_149__12_;
      r_149__11_ <= r_n_149__11_;
      r_149__10_ <= r_n_149__10_;
      r_149__9_ <= r_n_149__9_;
      r_149__8_ <= r_n_149__8_;
      r_149__7_ <= r_n_149__7_;
      r_149__6_ <= r_n_149__6_;
      r_149__5_ <= r_n_149__5_;
      r_149__4_ <= r_n_149__4_;
      r_149__3_ <= r_n_149__3_;
      r_149__2_ <= r_n_149__2_;
      r_149__1_ <= r_n_149__1_;
      r_149__0_ <= r_n_149__0_;
    end 
    if(N3734) begin
      r_150__63_ <= r_n_150__63_;
      r_150__62_ <= r_n_150__62_;
      r_150__61_ <= r_n_150__61_;
      r_150__60_ <= r_n_150__60_;
      r_150__59_ <= r_n_150__59_;
      r_150__58_ <= r_n_150__58_;
      r_150__57_ <= r_n_150__57_;
      r_150__56_ <= r_n_150__56_;
      r_150__55_ <= r_n_150__55_;
      r_150__54_ <= r_n_150__54_;
      r_150__53_ <= r_n_150__53_;
      r_150__52_ <= r_n_150__52_;
      r_150__51_ <= r_n_150__51_;
      r_150__50_ <= r_n_150__50_;
      r_150__49_ <= r_n_150__49_;
      r_150__48_ <= r_n_150__48_;
      r_150__47_ <= r_n_150__47_;
      r_150__46_ <= r_n_150__46_;
      r_150__45_ <= r_n_150__45_;
      r_150__44_ <= r_n_150__44_;
      r_150__43_ <= r_n_150__43_;
      r_150__42_ <= r_n_150__42_;
      r_150__41_ <= r_n_150__41_;
      r_150__40_ <= r_n_150__40_;
      r_150__39_ <= r_n_150__39_;
      r_150__38_ <= r_n_150__38_;
      r_150__37_ <= r_n_150__37_;
      r_150__36_ <= r_n_150__36_;
      r_150__35_ <= r_n_150__35_;
      r_150__34_ <= r_n_150__34_;
      r_150__33_ <= r_n_150__33_;
      r_150__32_ <= r_n_150__32_;
      r_150__31_ <= r_n_150__31_;
      r_150__30_ <= r_n_150__30_;
      r_150__29_ <= r_n_150__29_;
      r_150__28_ <= r_n_150__28_;
      r_150__27_ <= r_n_150__27_;
      r_150__26_ <= r_n_150__26_;
      r_150__25_ <= r_n_150__25_;
      r_150__24_ <= r_n_150__24_;
      r_150__23_ <= r_n_150__23_;
      r_150__22_ <= r_n_150__22_;
      r_150__21_ <= r_n_150__21_;
      r_150__20_ <= r_n_150__20_;
      r_150__19_ <= r_n_150__19_;
      r_150__18_ <= r_n_150__18_;
      r_150__17_ <= r_n_150__17_;
      r_150__16_ <= r_n_150__16_;
      r_150__15_ <= r_n_150__15_;
      r_150__14_ <= r_n_150__14_;
      r_150__13_ <= r_n_150__13_;
      r_150__12_ <= r_n_150__12_;
      r_150__11_ <= r_n_150__11_;
      r_150__10_ <= r_n_150__10_;
      r_150__9_ <= r_n_150__9_;
      r_150__8_ <= r_n_150__8_;
      r_150__7_ <= r_n_150__7_;
      r_150__6_ <= r_n_150__6_;
      r_150__5_ <= r_n_150__5_;
      r_150__4_ <= r_n_150__4_;
      r_150__3_ <= r_n_150__3_;
      r_150__2_ <= r_n_150__2_;
      r_150__1_ <= r_n_150__1_;
      r_150__0_ <= r_n_150__0_;
    end 
    if(N3735) begin
      r_151__63_ <= r_n_151__63_;
      r_151__62_ <= r_n_151__62_;
      r_151__61_ <= r_n_151__61_;
      r_151__60_ <= r_n_151__60_;
      r_151__59_ <= r_n_151__59_;
      r_151__58_ <= r_n_151__58_;
      r_151__57_ <= r_n_151__57_;
      r_151__56_ <= r_n_151__56_;
      r_151__55_ <= r_n_151__55_;
      r_151__54_ <= r_n_151__54_;
      r_151__53_ <= r_n_151__53_;
      r_151__52_ <= r_n_151__52_;
      r_151__51_ <= r_n_151__51_;
      r_151__50_ <= r_n_151__50_;
      r_151__49_ <= r_n_151__49_;
      r_151__48_ <= r_n_151__48_;
      r_151__47_ <= r_n_151__47_;
      r_151__46_ <= r_n_151__46_;
      r_151__45_ <= r_n_151__45_;
      r_151__44_ <= r_n_151__44_;
      r_151__43_ <= r_n_151__43_;
      r_151__42_ <= r_n_151__42_;
      r_151__41_ <= r_n_151__41_;
      r_151__40_ <= r_n_151__40_;
      r_151__39_ <= r_n_151__39_;
      r_151__38_ <= r_n_151__38_;
      r_151__37_ <= r_n_151__37_;
      r_151__36_ <= r_n_151__36_;
      r_151__35_ <= r_n_151__35_;
      r_151__34_ <= r_n_151__34_;
      r_151__33_ <= r_n_151__33_;
      r_151__32_ <= r_n_151__32_;
      r_151__31_ <= r_n_151__31_;
      r_151__30_ <= r_n_151__30_;
      r_151__29_ <= r_n_151__29_;
      r_151__28_ <= r_n_151__28_;
      r_151__27_ <= r_n_151__27_;
      r_151__26_ <= r_n_151__26_;
      r_151__25_ <= r_n_151__25_;
      r_151__24_ <= r_n_151__24_;
      r_151__23_ <= r_n_151__23_;
      r_151__22_ <= r_n_151__22_;
      r_151__21_ <= r_n_151__21_;
      r_151__20_ <= r_n_151__20_;
      r_151__19_ <= r_n_151__19_;
      r_151__18_ <= r_n_151__18_;
      r_151__17_ <= r_n_151__17_;
      r_151__16_ <= r_n_151__16_;
      r_151__15_ <= r_n_151__15_;
      r_151__14_ <= r_n_151__14_;
      r_151__13_ <= r_n_151__13_;
      r_151__12_ <= r_n_151__12_;
      r_151__11_ <= r_n_151__11_;
      r_151__10_ <= r_n_151__10_;
      r_151__9_ <= r_n_151__9_;
      r_151__8_ <= r_n_151__8_;
      r_151__7_ <= r_n_151__7_;
      r_151__6_ <= r_n_151__6_;
      r_151__5_ <= r_n_151__5_;
      r_151__4_ <= r_n_151__4_;
      r_151__3_ <= r_n_151__3_;
      r_151__2_ <= r_n_151__2_;
      r_151__1_ <= r_n_151__1_;
      r_151__0_ <= r_n_151__0_;
    end 
    if(N3736) begin
      r_152__63_ <= r_n_152__63_;
      r_152__62_ <= r_n_152__62_;
      r_152__61_ <= r_n_152__61_;
      r_152__60_ <= r_n_152__60_;
      r_152__59_ <= r_n_152__59_;
      r_152__58_ <= r_n_152__58_;
      r_152__57_ <= r_n_152__57_;
      r_152__56_ <= r_n_152__56_;
      r_152__55_ <= r_n_152__55_;
      r_152__54_ <= r_n_152__54_;
      r_152__53_ <= r_n_152__53_;
      r_152__52_ <= r_n_152__52_;
      r_152__51_ <= r_n_152__51_;
      r_152__50_ <= r_n_152__50_;
      r_152__49_ <= r_n_152__49_;
      r_152__48_ <= r_n_152__48_;
      r_152__47_ <= r_n_152__47_;
      r_152__46_ <= r_n_152__46_;
      r_152__45_ <= r_n_152__45_;
      r_152__44_ <= r_n_152__44_;
      r_152__43_ <= r_n_152__43_;
      r_152__42_ <= r_n_152__42_;
      r_152__41_ <= r_n_152__41_;
      r_152__40_ <= r_n_152__40_;
      r_152__39_ <= r_n_152__39_;
      r_152__38_ <= r_n_152__38_;
      r_152__37_ <= r_n_152__37_;
      r_152__36_ <= r_n_152__36_;
      r_152__35_ <= r_n_152__35_;
      r_152__34_ <= r_n_152__34_;
      r_152__33_ <= r_n_152__33_;
      r_152__32_ <= r_n_152__32_;
      r_152__31_ <= r_n_152__31_;
      r_152__30_ <= r_n_152__30_;
      r_152__29_ <= r_n_152__29_;
      r_152__28_ <= r_n_152__28_;
      r_152__27_ <= r_n_152__27_;
      r_152__26_ <= r_n_152__26_;
      r_152__25_ <= r_n_152__25_;
      r_152__24_ <= r_n_152__24_;
      r_152__23_ <= r_n_152__23_;
      r_152__22_ <= r_n_152__22_;
      r_152__21_ <= r_n_152__21_;
      r_152__20_ <= r_n_152__20_;
      r_152__19_ <= r_n_152__19_;
      r_152__18_ <= r_n_152__18_;
      r_152__17_ <= r_n_152__17_;
      r_152__16_ <= r_n_152__16_;
      r_152__15_ <= r_n_152__15_;
      r_152__14_ <= r_n_152__14_;
      r_152__13_ <= r_n_152__13_;
      r_152__12_ <= r_n_152__12_;
      r_152__11_ <= r_n_152__11_;
      r_152__10_ <= r_n_152__10_;
      r_152__9_ <= r_n_152__9_;
      r_152__8_ <= r_n_152__8_;
      r_152__7_ <= r_n_152__7_;
      r_152__6_ <= r_n_152__6_;
      r_152__5_ <= r_n_152__5_;
      r_152__4_ <= r_n_152__4_;
      r_152__3_ <= r_n_152__3_;
      r_152__2_ <= r_n_152__2_;
      r_152__1_ <= r_n_152__1_;
      r_152__0_ <= r_n_152__0_;
    end 
    if(N3737) begin
      r_153__63_ <= r_n_153__63_;
      r_153__62_ <= r_n_153__62_;
      r_153__61_ <= r_n_153__61_;
      r_153__60_ <= r_n_153__60_;
      r_153__59_ <= r_n_153__59_;
      r_153__58_ <= r_n_153__58_;
      r_153__57_ <= r_n_153__57_;
      r_153__56_ <= r_n_153__56_;
      r_153__55_ <= r_n_153__55_;
      r_153__54_ <= r_n_153__54_;
      r_153__53_ <= r_n_153__53_;
      r_153__52_ <= r_n_153__52_;
      r_153__51_ <= r_n_153__51_;
      r_153__50_ <= r_n_153__50_;
      r_153__49_ <= r_n_153__49_;
      r_153__48_ <= r_n_153__48_;
      r_153__47_ <= r_n_153__47_;
      r_153__46_ <= r_n_153__46_;
      r_153__45_ <= r_n_153__45_;
      r_153__44_ <= r_n_153__44_;
      r_153__43_ <= r_n_153__43_;
      r_153__42_ <= r_n_153__42_;
      r_153__41_ <= r_n_153__41_;
      r_153__40_ <= r_n_153__40_;
      r_153__39_ <= r_n_153__39_;
      r_153__38_ <= r_n_153__38_;
      r_153__37_ <= r_n_153__37_;
      r_153__36_ <= r_n_153__36_;
      r_153__35_ <= r_n_153__35_;
      r_153__34_ <= r_n_153__34_;
      r_153__33_ <= r_n_153__33_;
      r_153__32_ <= r_n_153__32_;
      r_153__31_ <= r_n_153__31_;
      r_153__30_ <= r_n_153__30_;
      r_153__29_ <= r_n_153__29_;
      r_153__28_ <= r_n_153__28_;
      r_153__27_ <= r_n_153__27_;
      r_153__26_ <= r_n_153__26_;
      r_153__25_ <= r_n_153__25_;
      r_153__24_ <= r_n_153__24_;
      r_153__23_ <= r_n_153__23_;
      r_153__22_ <= r_n_153__22_;
      r_153__21_ <= r_n_153__21_;
      r_153__20_ <= r_n_153__20_;
      r_153__19_ <= r_n_153__19_;
      r_153__18_ <= r_n_153__18_;
      r_153__17_ <= r_n_153__17_;
      r_153__16_ <= r_n_153__16_;
      r_153__15_ <= r_n_153__15_;
      r_153__14_ <= r_n_153__14_;
      r_153__13_ <= r_n_153__13_;
      r_153__12_ <= r_n_153__12_;
      r_153__11_ <= r_n_153__11_;
      r_153__10_ <= r_n_153__10_;
      r_153__9_ <= r_n_153__9_;
      r_153__8_ <= r_n_153__8_;
      r_153__7_ <= r_n_153__7_;
      r_153__6_ <= r_n_153__6_;
      r_153__5_ <= r_n_153__5_;
      r_153__4_ <= r_n_153__4_;
      r_153__3_ <= r_n_153__3_;
      r_153__2_ <= r_n_153__2_;
      r_153__1_ <= r_n_153__1_;
      r_153__0_ <= r_n_153__0_;
    end 
    if(N3738) begin
      r_154__63_ <= r_n_154__63_;
      r_154__62_ <= r_n_154__62_;
      r_154__61_ <= r_n_154__61_;
      r_154__60_ <= r_n_154__60_;
      r_154__59_ <= r_n_154__59_;
      r_154__58_ <= r_n_154__58_;
      r_154__57_ <= r_n_154__57_;
      r_154__56_ <= r_n_154__56_;
      r_154__55_ <= r_n_154__55_;
      r_154__54_ <= r_n_154__54_;
      r_154__53_ <= r_n_154__53_;
      r_154__52_ <= r_n_154__52_;
      r_154__51_ <= r_n_154__51_;
      r_154__50_ <= r_n_154__50_;
      r_154__49_ <= r_n_154__49_;
      r_154__48_ <= r_n_154__48_;
      r_154__47_ <= r_n_154__47_;
      r_154__46_ <= r_n_154__46_;
      r_154__45_ <= r_n_154__45_;
      r_154__44_ <= r_n_154__44_;
      r_154__43_ <= r_n_154__43_;
      r_154__42_ <= r_n_154__42_;
      r_154__41_ <= r_n_154__41_;
      r_154__40_ <= r_n_154__40_;
      r_154__39_ <= r_n_154__39_;
      r_154__38_ <= r_n_154__38_;
      r_154__37_ <= r_n_154__37_;
      r_154__36_ <= r_n_154__36_;
      r_154__35_ <= r_n_154__35_;
      r_154__34_ <= r_n_154__34_;
      r_154__33_ <= r_n_154__33_;
      r_154__32_ <= r_n_154__32_;
      r_154__31_ <= r_n_154__31_;
      r_154__30_ <= r_n_154__30_;
      r_154__29_ <= r_n_154__29_;
      r_154__28_ <= r_n_154__28_;
      r_154__27_ <= r_n_154__27_;
      r_154__26_ <= r_n_154__26_;
      r_154__25_ <= r_n_154__25_;
      r_154__24_ <= r_n_154__24_;
      r_154__23_ <= r_n_154__23_;
      r_154__22_ <= r_n_154__22_;
      r_154__21_ <= r_n_154__21_;
      r_154__20_ <= r_n_154__20_;
      r_154__19_ <= r_n_154__19_;
      r_154__18_ <= r_n_154__18_;
      r_154__17_ <= r_n_154__17_;
      r_154__16_ <= r_n_154__16_;
      r_154__15_ <= r_n_154__15_;
      r_154__14_ <= r_n_154__14_;
      r_154__13_ <= r_n_154__13_;
      r_154__12_ <= r_n_154__12_;
      r_154__11_ <= r_n_154__11_;
      r_154__10_ <= r_n_154__10_;
      r_154__9_ <= r_n_154__9_;
      r_154__8_ <= r_n_154__8_;
      r_154__7_ <= r_n_154__7_;
      r_154__6_ <= r_n_154__6_;
      r_154__5_ <= r_n_154__5_;
      r_154__4_ <= r_n_154__4_;
      r_154__3_ <= r_n_154__3_;
      r_154__2_ <= r_n_154__2_;
      r_154__1_ <= r_n_154__1_;
      r_154__0_ <= r_n_154__0_;
    end 
    if(N3739) begin
      r_155__63_ <= r_n_155__63_;
      r_155__62_ <= r_n_155__62_;
      r_155__61_ <= r_n_155__61_;
      r_155__60_ <= r_n_155__60_;
      r_155__59_ <= r_n_155__59_;
      r_155__58_ <= r_n_155__58_;
      r_155__57_ <= r_n_155__57_;
      r_155__56_ <= r_n_155__56_;
      r_155__55_ <= r_n_155__55_;
      r_155__54_ <= r_n_155__54_;
      r_155__53_ <= r_n_155__53_;
      r_155__52_ <= r_n_155__52_;
      r_155__51_ <= r_n_155__51_;
      r_155__50_ <= r_n_155__50_;
      r_155__49_ <= r_n_155__49_;
      r_155__48_ <= r_n_155__48_;
      r_155__47_ <= r_n_155__47_;
      r_155__46_ <= r_n_155__46_;
      r_155__45_ <= r_n_155__45_;
      r_155__44_ <= r_n_155__44_;
      r_155__43_ <= r_n_155__43_;
      r_155__42_ <= r_n_155__42_;
      r_155__41_ <= r_n_155__41_;
      r_155__40_ <= r_n_155__40_;
      r_155__39_ <= r_n_155__39_;
      r_155__38_ <= r_n_155__38_;
      r_155__37_ <= r_n_155__37_;
      r_155__36_ <= r_n_155__36_;
      r_155__35_ <= r_n_155__35_;
      r_155__34_ <= r_n_155__34_;
      r_155__33_ <= r_n_155__33_;
      r_155__32_ <= r_n_155__32_;
      r_155__31_ <= r_n_155__31_;
      r_155__30_ <= r_n_155__30_;
      r_155__29_ <= r_n_155__29_;
      r_155__28_ <= r_n_155__28_;
      r_155__27_ <= r_n_155__27_;
      r_155__26_ <= r_n_155__26_;
      r_155__25_ <= r_n_155__25_;
      r_155__24_ <= r_n_155__24_;
      r_155__23_ <= r_n_155__23_;
      r_155__22_ <= r_n_155__22_;
      r_155__21_ <= r_n_155__21_;
      r_155__20_ <= r_n_155__20_;
      r_155__19_ <= r_n_155__19_;
      r_155__18_ <= r_n_155__18_;
      r_155__17_ <= r_n_155__17_;
      r_155__16_ <= r_n_155__16_;
      r_155__15_ <= r_n_155__15_;
      r_155__14_ <= r_n_155__14_;
      r_155__13_ <= r_n_155__13_;
      r_155__12_ <= r_n_155__12_;
      r_155__11_ <= r_n_155__11_;
      r_155__10_ <= r_n_155__10_;
      r_155__9_ <= r_n_155__9_;
      r_155__8_ <= r_n_155__8_;
      r_155__7_ <= r_n_155__7_;
      r_155__6_ <= r_n_155__6_;
      r_155__5_ <= r_n_155__5_;
      r_155__4_ <= r_n_155__4_;
      r_155__3_ <= r_n_155__3_;
      r_155__2_ <= r_n_155__2_;
      r_155__1_ <= r_n_155__1_;
      r_155__0_ <= r_n_155__0_;
    end 
    if(N3740) begin
      r_156__63_ <= r_n_156__63_;
      r_156__62_ <= r_n_156__62_;
      r_156__61_ <= r_n_156__61_;
      r_156__60_ <= r_n_156__60_;
      r_156__59_ <= r_n_156__59_;
      r_156__58_ <= r_n_156__58_;
      r_156__57_ <= r_n_156__57_;
      r_156__56_ <= r_n_156__56_;
      r_156__55_ <= r_n_156__55_;
      r_156__54_ <= r_n_156__54_;
      r_156__53_ <= r_n_156__53_;
      r_156__52_ <= r_n_156__52_;
      r_156__51_ <= r_n_156__51_;
      r_156__50_ <= r_n_156__50_;
      r_156__49_ <= r_n_156__49_;
      r_156__48_ <= r_n_156__48_;
      r_156__47_ <= r_n_156__47_;
      r_156__46_ <= r_n_156__46_;
      r_156__45_ <= r_n_156__45_;
      r_156__44_ <= r_n_156__44_;
      r_156__43_ <= r_n_156__43_;
      r_156__42_ <= r_n_156__42_;
      r_156__41_ <= r_n_156__41_;
      r_156__40_ <= r_n_156__40_;
      r_156__39_ <= r_n_156__39_;
      r_156__38_ <= r_n_156__38_;
      r_156__37_ <= r_n_156__37_;
      r_156__36_ <= r_n_156__36_;
      r_156__35_ <= r_n_156__35_;
      r_156__34_ <= r_n_156__34_;
      r_156__33_ <= r_n_156__33_;
      r_156__32_ <= r_n_156__32_;
      r_156__31_ <= r_n_156__31_;
      r_156__30_ <= r_n_156__30_;
      r_156__29_ <= r_n_156__29_;
      r_156__28_ <= r_n_156__28_;
      r_156__27_ <= r_n_156__27_;
      r_156__26_ <= r_n_156__26_;
      r_156__25_ <= r_n_156__25_;
      r_156__24_ <= r_n_156__24_;
      r_156__23_ <= r_n_156__23_;
      r_156__22_ <= r_n_156__22_;
      r_156__21_ <= r_n_156__21_;
      r_156__20_ <= r_n_156__20_;
      r_156__19_ <= r_n_156__19_;
      r_156__18_ <= r_n_156__18_;
      r_156__17_ <= r_n_156__17_;
      r_156__16_ <= r_n_156__16_;
      r_156__15_ <= r_n_156__15_;
      r_156__14_ <= r_n_156__14_;
      r_156__13_ <= r_n_156__13_;
      r_156__12_ <= r_n_156__12_;
      r_156__11_ <= r_n_156__11_;
      r_156__10_ <= r_n_156__10_;
      r_156__9_ <= r_n_156__9_;
      r_156__8_ <= r_n_156__8_;
      r_156__7_ <= r_n_156__7_;
      r_156__6_ <= r_n_156__6_;
      r_156__5_ <= r_n_156__5_;
      r_156__4_ <= r_n_156__4_;
      r_156__3_ <= r_n_156__3_;
      r_156__2_ <= r_n_156__2_;
      r_156__1_ <= r_n_156__1_;
      r_156__0_ <= r_n_156__0_;
    end 
    if(N3741) begin
      r_157__63_ <= r_n_157__63_;
      r_157__62_ <= r_n_157__62_;
      r_157__61_ <= r_n_157__61_;
      r_157__60_ <= r_n_157__60_;
      r_157__59_ <= r_n_157__59_;
      r_157__58_ <= r_n_157__58_;
      r_157__57_ <= r_n_157__57_;
      r_157__56_ <= r_n_157__56_;
      r_157__55_ <= r_n_157__55_;
      r_157__54_ <= r_n_157__54_;
      r_157__53_ <= r_n_157__53_;
      r_157__52_ <= r_n_157__52_;
      r_157__51_ <= r_n_157__51_;
      r_157__50_ <= r_n_157__50_;
      r_157__49_ <= r_n_157__49_;
      r_157__48_ <= r_n_157__48_;
      r_157__47_ <= r_n_157__47_;
      r_157__46_ <= r_n_157__46_;
      r_157__45_ <= r_n_157__45_;
      r_157__44_ <= r_n_157__44_;
      r_157__43_ <= r_n_157__43_;
      r_157__42_ <= r_n_157__42_;
      r_157__41_ <= r_n_157__41_;
      r_157__40_ <= r_n_157__40_;
      r_157__39_ <= r_n_157__39_;
      r_157__38_ <= r_n_157__38_;
      r_157__37_ <= r_n_157__37_;
      r_157__36_ <= r_n_157__36_;
      r_157__35_ <= r_n_157__35_;
      r_157__34_ <= r_n_157__34_;
      r_157__33_ <= r_n_157__33_;
      r_157__32_ <= r_n_157__32_;
      r_157__31_ <= r_n_157__31_;
      r_157__30_ <= r_n_157__30_;
      r_157__29_ <= r_n_157__29_;
      r_157__28_ <= r_n_157__28_;
      r_157__27_ <= r_n_157__27_;
      r_157__26_ <= r_n_157__26_;
      r_157__25_ <= r_n_157__25_;
      r_157__24_ <= r_n_157__24_;
      r_157__23_ <= r_n_157__23_;
      r_157__22_ <= r_n_157__22_;
      r_157__21_ <= r_n_157__21_;
      r_157__20_ <= r_n_157__20_;
      r_157__19_ <= r_n_157__19_;
      r_157__18_ <= r_n_157__18_;
      r_157__17_ <= r_n_157__17_;
      r_157__16_ <= r_n_157__16_;
      r_157__15_ <= r_n_157__15_;
      r_157__14_ <= r_n_157__14_;
      r_157__13_ <= r_n_157__13_;
      r_157__12_ <= r_n_157__12_;
      r_157__11_ <= r_n_157__11_;
      r_157__10_ <= r_n_157__10_;
      r_157__9_ <= r_n_157__9_;
      r_157__8_ <= r_n_157__8_;
      r_157__7_ <= r_n_157__7_;
      r_157__6_ <= r_n_157__6_;
      r_157__5_ <= r_n_157__5_;
      r_157__4_ <= r_n_157__4_;
      r_157__3_ <= r_n_157__3_;
      r_157__2_ <= r_n_157__2_;
      r_157__1_ <= r_n_157__1_;
      r_157__0_ <= r_n_157__0_;
    end 
    if(N3742) begin
      r_158__63_ <= r_n_158__63_;
      r_158__62_ <= r_n_158__62_;
      r_158__61_ <= r_n_158__61_;
      r_158__60_ <= r_n_158__60_;
      r_158__59_ <= r_n_158__59_;
      r_158__58_ <= r_n_158__58_;
      r_158__57_ <= r_n_158__57_;
      r_158__56_ <= r_n_158__56_;
      r_158__55_ <= r_n_158__55_;
      r_158__54_ <= r_n_158__54_;
      r_158__53_ <= r_n_158__53_;
      r_158__52_ <= r_n_158__52_;
      r_158__51_ <= r_n_158__51_;
      r_158__50_ <= r_n_158__50_;
      r_158__49_ <= r_n_158__49_;
      r_158__48_ <= r_n_158__48_;
      r_158__47_ <= r_n_158__47_;
      r_158__46_ <= r_n_158__46_;
      r_158__45_ <= r_n_158__45_;
      r_158__44_ <= r_n_158__44_;
      r_158__43_ <= r_n_158__43_;
      r_158__42_ <= r_n_158__42_;
      r_158__41_ <= r_n_158__41_;
      r_158__40_ <= r_n_158__40_;
      r_158__39_ <= r_n_158__39_;
      r_158__38_ <= r_n_158__38_;
      r_158__37_ <= r_n_158__37_;
      r_158__36_ <= r_n_158__36_;
      r_158__35_ <= r_n_158__35_;
      r_158__34_ <= r_n_158__34_;
      r_158__33_ <= r_n_158__33_;
      r_158__32_ <= r_n_158__32_;
      r_158__31_ <= r_n_158__31_;
      r_158__30_ <= r_n_158__30_;
      r_158__29_ <= r_n_158__29_;
      r_158__28_ <= r_n_158__28_;
      r_158__27_ <= r_n_158__27_;
      r_158__26_ <= r_n_158__26_;
      r_158__25_ <= r_n_158__25_;
      r_158__24_ <= r_n_158__24_;
      r_158__23_ <= r_n_158__23_;
      r_158__22_ <= r_n_158__22_;
      r_158__21_ <= r_n_158__21_;
      r_158__20_ <= r_n_158__20_;
      r_158__19_ <= r_n_158__19_;
      r_158__18_ <= r_n_158__18_;
      r_158__17_ <= r_n_158__17_;
      r_158__16_ <= r_n_158__16_;
      r_158__15_ <= r_n_158__15_;
      r_158__14_ <= r_n_158__14_;
      r_158__13_ <= r_n_158__13_;
      r_158__12_ <= r_n_158__12_;
      r_158__11_ <= r_n_158__11_;
      r_158__10_ <= r_n_158__10_;
      r_158__9_ <= r_n_158__9_;
      r_158__8_ <= r_n_158__8_;
      r_158__7_ <= r_n_158__7_;
      r_158__6_ <= r_n_158__6_;
      r_158__5_ <= r_n_158__5_;
      r_158__4_ <= r_n_158__4_;
      r_158__3_ <= r_n_158__3_;
      r_158__2_ <= r_n_158__2_;
      r_158__1_ <= r_n_158__1_;
      r_158__0_ <= r_n_158__0_;
    end 
    if(N3743) begin
      r_159__63_ <= r_n_159__63_;
      r_159__62_ <= r_n_159__62_;
      r_159__61_ <= r_n_159__61_;
      r_159__60_ <= r_n_159__60_;
      r_159__59_ <= r_n_159__59_;
      r_159__58_ <= r_n_159__58_;
      r_159__57_ <= r_n_159__57_;
      r_159__56_ <= r_n_159__56_;
      r_159__55_ <= r_n_159__55_;
      r_159__54_ <= r_n_159__54_;
      r_159__53_ <= r_n_159__53_;
      r_159__52_ <= r_n_159__52_;
      r_159__51_ <= r_n_159__51_;
      r_159__50_ <= r_n_159__50_;
      r_159__49_ <= r_n_159__49_;
      r_159__48_ <= r_n_159__48_;
      r_159__47_ <= r_n_159__47_;
      r_159__46_ <= r_n_159__46_;
      r_159__45_ <= r_n_159__45_;
      r_159__44_ <= r_n_159__44_;
      r_159__43_ <= r_n_159__43_;
      r_159__42_ <= r_n_159__42_;
      r_159__41_ <= r_n_159__41_;
      r_159__40_ <= r_n_159__40_;
      r_159__39_ <= r_n_159__39_;
      r_159__38_ <= r_n_159__38_;
      r_159__37_ <= r_n_159__37_;
      r_159__36_ <= r_n_159__36_;
      r_159__35_ <= r_n_159__35_;
      r_159__34_ <= r_n_159__34_;
      r_159__33_ <= r_n_159__33_;
      r_159__32_ <= r_n_159__32_;
      r_159__31_ <= r_n_159__31_;
      r_159__30_ <= r_n_159__30_;
      r_159__29_ <= r_n_159__29_;
      r_159__28_ <= r_n_159__28_;
      r_159__27_ <= r_n_159__27_;
      r_159__26_ <= r_n_159__26_;
      r_159__25_ <= r_n_159__25_;
      r_159__24_ <= r_n_159__24_;
      r_159__23_ <= r_n_159__23_;
      r_159__22_ <= r_n_159__22_;
      r_159__21_ <= r_n_159__21_;
      r_159__20_ <= r_n_159__20_;
      r_159__19_ <= r_n_159__19_;
      r_159__18_ <= r_n_159__18_;
      r_159__17_ <= r_n_159__17_;
      r_159__16_ <= r_n_159__16_;
      r_159__15_ <= r_n_159__15_;
      r_159__14_ <= r_n_159__14_;
      r_159__13_ <= r_n_159__13_;
      r_159__12_ <= r_n_159__12_;
      r_159__11_ <= r_n_159__11_;
      r_159__10_ <= r_n_159__10_;
      r_159__9_ <= r_n_159__9_;
      r_159__8_ <= r_n_159__8_;
      r_159__7_ <= r_n_159__7_;
      r_159__6_ <= r_n_159__6_;
      r_159__5_ <= r_n_159__5_;
      r_159__4_ <= r_n_159__4_;
      r_159__3_ <= r_n_159__3_;
      r_159__2_ <= r_n_159__2_;
      r_159__1_ <= r_n_159__1_;
      r_159__0_ <= r_n_159__0_;
    end 
    if(N3744) begin
      r_160__63_ <= r_n_160__63_;
      r_160__62_ <= r_n_160__62_;
      r_160__61_ <= r_n_160__61_;
      r_160__60_ <= r_n_160__60_;
      r_160__59_ <= r_n_160__59_;
      r_160__58_ <= r_n_160__58_;
      r_160__57_ <= r_n_160__57_;
      r_160__56_ <= r_n_160__56_;
      r_160__55_ <= r_n_160__55_;
      r_160__54_ <= r_n_160__54_;
      r_160__53_ <= r_n_160__53_;
      r_160__52_ <= r_n_160__52_;
      r_160__51_ <= r_n_160__51_;
      r_160__50_ <= r_n_160__50_;
      r_160__49_ <= r_n_160__49_;
      r_160__48_ <= r_n_160__48_;
      r_160__47_ <= r_n_160__47_;
      r_160__46_ <= r_n_160__46_;
      r_160__45_ <= r_n_160__45_;
      r_160__44_ <= r_n_160__44_;
      r_160__43_ <= r_n_160__43_;
      r_160__42_ <= r_n_160__42_;
      r_160__41_ <= r_n_160__41_;
      r_160__40_ <= r_n_160__40_;
      r_160__39_ <= r_n_160__39_;
      r_160__38_ <= r_n_160__38_;
      r_160__37_ <= r_n_160__37_;
      r_160__36_ <= r_n_160__36_;
      r_160__35_ <= r_n_160__35_;
      r_160__34_ <= r_n_160__34_;
      r_160__33_ <= r_n_160__33_;
      r_160__32_ <= r_n_160__32_;
      r_160__31_ <= r_n_160__31_;
      r_160__30_ <= r_n_160__30_;
      r_160__29_ <= r_n_160__29_;
      r_160__28_ <= r_n_160__28_;
      r_160__27_ <= r_n_160__27_;
      r_160__26_ <= r_n_160__26_;
      r_160__25_ <= r_n_160__25_;
      r_160__24_ <= r_n_160__24_;
      r_160__23_ <= r_n_160__23_;
      r_160__22_ <= r_n_160__22_;
      r_160__21_ <= r_n_160__21_;
      r_160__20_ <= r_n_160__20_;
      r_160__19_ <= r_n_160__19_;
      r_160__18_ <= r_n_160__18_;
      r_160__17_ <= r_n_160__17_;
      r_160__16_ <= r_n_160__16_;
      r_160__15_ <= r_n_160__15_;
      r_160__14_ <= r_n_160__14_;
      r_160__13_ <= r_n_160__13_;
      r_160__12_ <= r_n_160__12_;
      r_160__11_ <= r_n_160__11_;
      r_160__10_ <= r_n_160__10_;
      r_160__9_ <= r_n_160__9_;
      r_160__8_ <= r_n_160__8_;
      r_160__7_ <= r_n_160__7_;
      r_160__6_ <= r_n_160__6_;
      r_160__5_ <= r_n_160__5_;
      r_160__4_ <= r_n_160__4_;
      r_160__3_ <= r_n_160__3_;
      r_160__2_ <= r_n_160__2_;
      r_160__1_ <= r_n_160__1_;
      r_160__0_ <= r_n_160__0_;
    end 
    if(N3745) begin
      r_161__63_ <= r_n_161__63_;
      r_161__62_ <= r_n_161__62_;
      r_161__61_ <= r_n_161__61_;
      r_161__60_ <= r_n_161__60_;
      r_161__59_ <= r_n_161__59_;
      r_161__58_ <= r_n_161__58_;
      r_161__57_ <= r_n_161__57_;
      r_161__56_ <= r_n_161__56_;
      r_161__55_ <= r_n_161__55_;
      r_161__54_ <= r_n_161__54_;
      r_161__53_ <= r_n_161__53_;
      r_161__52_ <= r_n_161__52_;
      r_161__51_ <= r_n_161__51_;
      r_161__50_ <= r_n_161__50_;
      r_161__49_ <= r_n_161__49_;
      r_161__48_ <= r_n_161__48_;
      r_161__47_ <= r_n_161__47_;
      r_161__46_ <= r_n_161__46_;
      r_161__45_ <= r_n_161__45_;
      r_161__44_ <= r_n_161__44_;
      r_161__43_ <= r_n_161__43_;
      r_161__42_ <= r_n_161__42_;
      r_161__41_ <= r_n_161__41_;
      r_161__40_ <= r_n_161__40_;
      r_161__39_ <= r_n_161__39_;
      r_161__38_ <= r_n_161__38_;
      r_161__37_ <= r_n_161__37_;
      r_161__36_ <= r_n_161__36_;
      r_161__35_ <= r_n_161__35_;
      r_161__34_ <= r_n_161__34_;
      r_161__33_ <= r_n_161__33_;
      r_161__32_ <= r_n_161__32_;
      r_161__31_ <= r_n_161__31_;
      r_161__30_ <= r_n_161__30_;
      r_161__29_ <= r_n_161__29_;
      r_161__28_ <= r_n_161__28_;
      r_161__27_ <= r_n_161__27_;
      r_161__26_ <= r_n_161__26_;
      r_161__25_ <= r_n_161__25_;
      r_161__24_ <= r_n_161__24_;
      r_161__23_ <= r_n_161__23_;
      r_161__22_ <= r_n_161__22_;
      r_161__21_ <= r_n_161__21_;
      r_161__20_ <= r_n_161__20_;
      r_161__19_ <= r_n_161__19_;
      r_161__18_ <= r_n_161__18_;
      r_161__17_ <= r_n_161__17_;
      r_161__16_ <= r_n_161__16_;
      r_161__15_ <= r_n_161__15_;
      r_161__14_ <= r_n_161__14_;
      r_161__13_ <= r_n_161__13_;
      r_161__12_ <= r_n_161__12_;
      r_161__11_ <= r_n_161__11_;
      r_161__10_ <= r_n_161__10_;
      r_161__9_ <= r_n_161__9_;
      r_161__8_ <= r_n_161__8_;
      r_161__7_ <= r_n_161__7_;
      r_161__6_ <= r_n_161__6_;
      r_161__5_ <= r_n_161__5_;
      r_161__4_ <= r_n_161__4_;
      r_161__3_ <= r_n_161__3_;
      r_161__2_ <= r_n_161__2_;
      r_161__1_ <= r_n_161__1_;
      r_161__0_ <= r_n_161__0_;
    end 
    if(N3746) begin
      r_162__63_ <= r_n_162__63_;
      r_162__62_ <= r_n_162__62_;
      r_162__61_ <= r_n_162__61_;
      r_162__60_ <= r_n_162__60_;
      r_162__59_ <= r_n_162__59_;
      r_162__58_ <= r_n_162__58_;
      r_162__57_ <= r_n_162__57_;
      r_162__56_ <= r_n_162__56_;
      r_162__55_ <= r_n_162__55_;
      r_162__54_ <= r_n_162__54_;
      r_162__53_ <= r_n_162__53_;
      r_162__52_ <= r_n_162__52_;
      r_162__51_ <= r_n_162__51_;
      r_162__50_ <= r_n_162__50_;
      r_162__49_ <= r_n_162__49_;
      r_162__48_ <= r_n_162__48_;
      r_162__47_ <= r_n_162__47_;
      r_162__46_ <= r_n_162__46_;
      r_162__45_ <= r_n_162__45_;
      r_162__44_ <= r_n_162__44_;
      r_162__43_ <= r_n_162__43_;
      r_162__42_ <= r_n_162__42_;
      r_162__41_ <= r_n_162__41_;
      r_162__40_ <= r_n_162__40_;
      r_162__39_ <= r_n_162__39_;
      r_162__38_ <= r_n_162__38_;
      r_162__37_ <= r_n_162__37_;
      r_162__36_ <= r_n_162__36_;
      r_162__35_ <= r_n_162__35_;
      r_162__34_ <= r_n_162__34_;
      r_162__33_ <= r_n_162__33_;
      r_162__32_ <= r_n_162__32_;
      r_162__31_ <= r_n_162__31_;
      r_162__30_ <= r_n_162__30_;
      r_162__29_ <= r_n_162__29_;
      r_162__28_ <= r_n_162__28_;
      r_162__27_ <= r_n_162__27_;
      r_162__26_ <= r_n_162__26_;
      r_162__25_ <= r_n_162__25_;
      r_162__24_ <= r_n_162__24_;
      r_162__23_ <= r_n_162__23_;
      r_162__22_ <= r_n_162__22_;
      r_162__21_ <= r_n_162__21_;
      r_162__20_ <= r_n_162__20_;
      r_162__19_ <= r_n_162__19_;
      r_162__18_ <= r_n_162__18_;
      r_162__17_ <= r_n_162__17_;
      r_162__16_ <= r_n_162__16_;
      r_162__15_ <= r_n_162__15_;
      r_162__14_ <= r_n_162__14_;
      r_162__13_ <= r_n_162__13_;
      r_162__12_ <= r_n_162__12_;
      r_162__11_ <= r_n_162__11_;
      r_162__10_ <= r_n_162__10_;
      r_162__9_ <= r_n_162__9_;
      r_162__8_ <= r_n_162__8_;
      r_162__7_ <= r_n_162__7_;
      r_162__6_ <= r_n_162__6_;
      r_162__5_ <= r_n_162__5_;
      r_162__4_ <= r_n_162__4_;
      r_162__3_ <= r_n_162__3_;
      r_162__2_ <= r_n_162__2_;
      r_162__1_ <= r_n_162__1_;
      r_162__0_ <= r_n_162__0_;
    end 
    if(N3747) begin
      r_163__63_ <= r_n_163__63_;
      r_163__62_ <= r_n_163__62_;
      r_163__61_ <= r_n_163__61_;
      r_163__60_ <= r_n_163__60_;
      r_163__59_ <= r_n_163__59_;
      r_163__58_ <= r_n_163__58_;
      r_163__57_ <= r_n_163__57_;
      r_163__56_ <= r_n_163__56_;
      r_163__55_ <= r_n_163__55_;
      r_163__54_ <= r_n_163__54_;
      r_163__53_ <= r_n_163__53_;
      r_163__52_ <= r_n_163__52_;
      r_163__51_ <= r_n_163__51_;
      r_163__50_ <= r_n_163__50_;
      r_163__49_ <= r_n_163__49_;
      r_163__48_ <= r_n_163__48_;
      r_163__47_ <= r_n_163__47_;
      r_163__46_ <= r_n_163__46_;
      r_163__45_ <= r_n_163__45_;
      r_163__44_ <= r_n_163__44_;
      r_163__43_ <= r_n_163__43_;
      r_163__42_ <= r_n_163__42_;
      r_163__41_ <= r_n_163__41_;
      r_163__40_ <= r_n_163__40_;
      r_163__39_ <= r_n_163__39_;
      r_163__38_ <= r_n_163__38_;
      r_163__37_ <= r_n_163__37_;
      r_163__36_ <= r_n_163__36_;
      r_163__35_ <= r_n_163__35_;
      r_163__34_ <= r_n_163__34_;
      r_163__33_ <= r_n_163__33_;
      r_163__32_ <= r_n_163__32_;
      r_163__31_ <= r_n_163__31_;
      r_163__30_ <= r_n_163__30_;
      r_163__29_ <= r_n_163__29_;
      r_163__28_ <= r_n_163__28_;
      r_163__27_ <= r_n_163__27_;
      r_163__26_ <= r_n_163__26_;
      r_163__25_ <= r_n_163__25_;
      r_163__24_ <= r_n_163__24_;
      r_163__23_ <= r_n_163__23_;
      r_163__22_ <= r_n_163__22_;
      r_163__21_ <= r_n_163__21_;
      r_163__20_ <= r_n_163__20_;
      r_163__19_ <= r_n_163__19_;
      r_163__18_ <= r_n_163__18_;
      r_163__17_ <= r_n_163__17_;
      r_163__16_ <= r_n_163__16_;
      r_163__15_ <= r_n_163__15_;
      r_163__14_ <= r_n_163__14_;
      r_163__13_ <= r_n_163__13_;
      r_163__12_ <= r_n_163__12_;
      r_163__11_ <= r_n_163__11_;
      r_163__10_ <= r_n_163__10_;
      r_163__9_ <= r_n_163__9_;
      r_163__8_ <= r_n_163__8_;
      r_163__7_ <= r_n_163__7_;
      r_163__6_ <= r_n_163__6_;
      r_163__5_ <= r_n_163__5_;
      r_163__4_ <= r_n_163__4_;
      r_163__3_ <= r_n_163__3_;
      r_163__2_ <= r_n_163__2_;
      r_163__1_ <= r_n_163__1_;
      r_163__0_ <= r_n_163__0_;
    end 
    if(N3748) begin
      r_164__63_ <= r_n_164__63_;
      r_164__62_ <= r_n_164__62_;
      r_164__61_ <= r_n_164__61_;
      r_164__60_ <= r_n_164__60_;
      r_164__59_ <= r_n_164__59_;
      r_164__58_ <= r_n_164__58_;
      r_164__57_ <= r_n_164__57_;
      r_164__56_ <= r_n_164__56_;
      r_164__55_ <= r_n_164__55_;
      r_164__54_ <= r_n_164__54_;
      r_164__53_ <= r_n_164__53_;
      r_164__52_ <= r_n_164__52_;
      r_164__51_ <= r_n_164__51_;
      r_164__50_ <= r_n_164__50_;
      r_164__49_ <= r_n_164__49_;
      r_164__48_ <= r_n_164__48_;
      r_164__47_ <= r_n_164__47_;
      r_164__46_ <= r_n_164__46_;
      r_164__45_ <= r_n_164__45_;
      r_164__44_ <= r_n_164__44_;
      r_164__43_ <= r_n_164__43_;
      r_164__42_ <= r_n_164__42_;
      r_164__41_ <= r_n_164__41_;
      r_164__40_ <= r_n_164__40_;
      r_164__39_ <= r_n_164__39_;
      r_164__38_ <= r_n_164__38_;
      r_164__37_ <= r_n_164__37_;
      r_164__36_ <= r_n_164__36_;
      r_164__35_ <= r_n_164__35_;
      r_164__34_ <= r_n_164__34_;
      r_164__33_ <= r_n_164__33_;
      r_164__32_ <= r_n_164__32_;
      r_164__31_ <= r_n_164__31_;
      r_164__30_ <= r_n_164__30_;
      r_164__29_ <= r_n_164__29_;
      r_164__28_ <= r_n_164__28_;
      r_164__27_ <= r_n_164__27_;
      r_164__26_ <= r_n_164__26_;
      r_164__25_ <= r_n_164__25_;
      r_164__24_ <= r_n_164__24_;
      r_164__23_ <= r_n_164__23_;
      r_164__22_ <= r_n_164__22_;
      r_164__21_ <= r_n_164__21_;
      r_164__20_ <= r_n_164__20_;
      r_164__19_ <= r_n_164__19_;
      r_164__18_ <= r_n_164__18_;
      r_164__17_ <= r_n_164__17_;
      r_164__16_ <= r_n_164__16_;
      r_164__15_ <= r_n_164__15_;
      r_164__14_ <= r_n_164__14_;
      r_164__13_ <= r_n_164__13_;
      r_164__12_ <= r_n_164__12_;
      r_164__11_ <= r_n_164__11_;
      r_164__10_ <= r_n_164__10_;
      r_164__9_ <= r_n_164__9_;
      r_164__8_ <= r_n_164__8_;
      r_164__7_ <= r_n_164__7_;
      r_164__6_ <= r_n_164__6_;
      r_164__5_ <= r_n_164__5_;
      r_164__4_ <= r_n_164__4_;
      r_164__3_ <= r_n_164__3_;
      r_164__2_ <= r_n_164__2_;
      r_164__1_ <= r_n_164__1_;
      r_164__0_ <= r_n_164__0_;
    end 
    if(N3749) begin
      r_165__63_ <= r_n_165__63_;
      r_165__62_ <= r_n_165__62_;
      r_165__61_ <= r_n_165__61_;
      r_165__60_ <= r_n_165__60_;
      r_165__59_ <= r_n_165__59_;
      r_165__58_ <= r_n_165__58_;
      r_165__57_ <= r_n_165__57_;
      r_165__56_ <= r_n_165__56_;
      r_165__55_ <= r_n_165__55_;
      r_165__54_ <= r_n_165__54_;
      r_165__53_ <= r_n_165__53_;
      r_165__52_ <= r_n_165__52_;
      r_165__51_ <= r_n_165__51_;
      r_165__50_ <= r_n_165__50_;
      r_165__49_ <= r_n_165__49_;
      r_165__48_ <= r_n_165__48_;
      r_165__47_ <= r_n_165__47_;
      r_165__46_ <= r_n_165__46_;
      r_165__45_ <= r_n_165__45_;
      r_165__44_ <= r_n_165__44_;
      r_165__43_ <= r_n_165__43_;
      r_165__42_ <= r_n_165__42_;
      r_165__41_ <= r_n_165__41_;
      r_165__40_ <= r_n_165__40_;
      r_165__39_ <= r_n_165__39_;
      r_165__38_ <= r_n_165__38_;
      r_165__37_ <= r_n_165__37_;
      r_165__36_ <= r_n_165__36_;
      r_165__35_ <= r_n_165__35_;
      r_165__34_ <= r_n_165__34_;
      r_165__33_ <= r_n_165__33_;
      r_165__32_ <= r_n_165__32_;
      r_165__31_ <= r_n_165__31_;
      r_165__30_ <= r_n_165__30_;
      r_165__29_ <= r_n_165__29_;
      r_165__28_ <= r_n_165__28_;
      r_165__27_ <= r_n_165__27_;
      r_165__26_ <= r_n_165__26_;
      r_165__25_ <= r_n_165__25_;
      r_165__24_ <= r_n_165__24_;
      r_165__23_ <= r_n_165__23_;
      r_165__22_ <= r_n_165__22_;
      r_165__21_ <= r_n_165__21_;
      r_165__20_ <= r_n_165__20_;
      r_165__19_ <= r_n_165__19_;
      r_165__18_ <= r_n_165__18_;
      r_165__17_ <= r_n_165__17_;
      r_165__16_ <= r_n_165__16_;
      r_165__15_ <= r_n_165__15_;
      r_165__14_ <= r_n_165__14_;
      r_165__13_ <= r_n_165__13_;
      r_165__12_ <= r_n_165__12_;
      r_165__11_ <= r_n_165__11_;
      r_165__10_ <= r_n_165__10_;
      r_165__9_ <= r_n_165__9_;
      r_165__8_ <= r_n_165__8_;
      r_165__7_ <= r_n_165__7_;
      r_165__6_ <= r_n_165__6_;
      r_165__5_ <= r_n_165__5_;
      r_165__4_ <= r_n_165__4_;
      r_165__3_ <= r_n_165__3_;
      r_165__2_ <= r_n_165__2_;
      r_165__1_ <= r_n_165__1_;
      r_165__0_ <= r_n_165__0_;
    end 
    if(N3750) begin
      r_166__63_ <= r_n_166__63_;
      r_166__62_ <= r_n_166__62_;
      r_166__61_ <= r_n_166__61_;
      r_166__60_ <= r_n_166__60_;
      r_166__59_ <= r_n_166__59_;
      r_166__58_ <= r_n_166__58_;
      r_166__57_ <= r_n_166__57_;
      r_166__56_ <= r_n_166__56_;
      r_166__55_ <= r_n_166__55_;
      r_166__54_ <= r_n_166__54_;
      r_166__53_ <= r_n_166__53_;
      r_166__52_ <= r_n_166__52_;
      r_166__51_ <= r_n_166__51_;
      r_166__50_ <= r_n_166__50_;
      r_166__49_ <= r_n_166__49_;
      r_166__48_ <= r_n_166__48_;
      r_166__47_ <= r_n_166__47_;
      r_166__46_ <= r_n_166__46_;
      r_166__45_ <= r_n_166__45_;
      r_166__44_ <= r_n_166__44_;
      r_166__43_ <= r_n_166__43_;
      r_166__42_ <= r_n_166__42_;
      r_166__41_ <= r_n_166__41_;
      r_166__40_ <= r_n_166__40_;
      r_166__39_ <= r_n_166__39_;
      r_166__38_ <= r_n_166__38_;
      r_166__37_ <= r_n_166__37_;
      r_166__36_ <= r_n_166__36_;
      r_166__35_ <= r_n_166__35_;
      r_166__34_ <= r_n_166__34_;
      r_166__33_ <= r_n_166__33_;
      r_166__32_ <= r_n_166__32_;
      r_166__31_ <= r_n_166__31_;
      r_166__30_ <= r_n_166__30_;
      r_166__29_ <= r_n_166__29_;
      r_166__28_ <= r_n_166__28_;
      r_166__27_ <= r_n_166__27_;
      r_166__26_ <= r_n_166__26_;
      r_166__25_ <= r_n_166__25_;
      r_166__24_ <= r_n_166__24_;
      r_166__23_ <= r_n_166__23_;
      r_166__22_ <= r_n_166__22_;
      r_166__21_ <= r_n_166__21_;
      r_166__20_ <= r_n_166__20_;
      r_166__19_ <= r_n_166__19_;
      r_166__18_ <= r_n_166__18_;
      r_166__17_ <= r_n_166__17_;
      r_166__16_ <= r_n_166__16_;
      r_166__15_ <= r_n_166__15_;
      r_166__14_ <= r_n_166__14_;
      r_166__13_ <= r_n_166__13_;
      r_166__12_ <= r_n_166__12_;
      r_166__11_ <= r_n_166__11_;
      r_166__10_ <= r_n_166__10_;
      r_166__9_ <= r_n_166__9_;
      r_166__8_ <= r_n_166__8_;
      r_166__7_ <= r_n_166__7_;
      r_166__6_ <= r_n_166__6_;
      r_166__5_ <= r_n_166__5_;
      r_166__4_ <= r_n_166__4_;
      r_166__3_ <= r_n_166__3_;
      r_166__2_ <= r_n_166__2_;
      r_166__1_ <= r_n_166__1_;
      r_166__0_ <= r_n_166__0_;
    end 
    if(N3751) begin
      r_167__63_ <= r_n_167__63_;
      r_167__62_ <= r_n_167__62_;
      r_167__61_ <= r_n_167__61_;
      r_167__60_ <= r_n_167__60_;
      r_167__59_ <= r_n_167__59_;
      r_167__58_ <= r_n_167__58_;
      r_167__57_ <= r_n_167__57_;
      r_167__56_ <= r_n_167__56_;
      r_167__55_ <= r_n_167__55_;
      r_167__54_ <= r_n_167__54_;
      r_167__53_ <= r_n_167__53_;
      r_167__52_ <= r_n_167__52_;
      r_167__51_ <= r_n_167__51_;
      r_167__50_ <= r_n_167__50_;
      r_167__49_ <= r_n_167__49_;
      r_167__48_ <= r_n_167__48_;
      r_167__47_ <= r_n_167__47_;
      r_167__46_ <= r_n_167__46_;
      r_167__45_ <= r_n_167__45_;
      r_167__44_ <= r_n_167__44_;
      r_167__43_ <= r_n_167__43_;
      r_167__42_ <= r_n_167__42_;
      r_167__41_ <= r_n_167__41_;
      r_167__40_ <= r_n_167__40_;
      r_167__39_ <= r_n_167__39_;
      r_167__38_ <= r_n_167__38_;
      r_167__37_ <= r_n_167__37_;
      r_167__36_ <= r_n_167__36_;
      r_167__35_ <= r_n_167__35_;
      r_167__34_ <= r_n_167__34_;
      r_167__33_ <= r_n_167__33_;
      r_167__32_ <= r_n_167__32_;
      r_167__31_ <= r_n_167__31_;
      r_167__30_ <= r_n_167__30_;
      r_167__29_ <= r_n_167__29_;
      r_167__28_ <= r_n_167__28_;
      r_167__27_ <= r_n_167__27_;
      r_167__26_ <= r_n_167__26_;
      r_167__25_ <= r_n_167__25_;
      r_167__24_ <= r_n_167__24_;
      r_167__23_ <= r_n_167__23_;
      r_167__22_ <= r_n_167__22_;
      r_167__21_ <= r_n_167__21_;
      r_167__20_ <= r_n_167__20_;
      r_167__19_ <= r_n_167__19_;
      r_167__18_ <= r_n_167__18_;
      r_167__17_ <= r_n_167__17_;
      r_167__16_ <= r_n_167__16_;
      r_167__15_ <= r_n_167__15_;
      r_167__14_ <= r_n_167__14_;
      r_167__13_ <= r_n_167__13_;
      r_167__12_ <= r_n_167__12_;
      r_167__11_ <= r_n_167__11_;
      r_167__10_ <= r_n_167__10_;
      r_167__9_ <= r_n_167__9_;
      r_167__8_ <= r_n_167__8_;
      r_167__7_ <= r_n_167__7_;
      r_167__6_ <= r_n_167__6_;
      r_167__5_ <= r_n_167__5_;
      r_167__4_ <= r_n_167__4_;
      r_167__3_ <= r_n_167__3_;
      r_167__2_ <= r_n_167__2_;
      r_167__1_ <= r_n_167__1_;
      r_167__0_ <= r_n_167__0_;
    end 
    if(N3752) begin
      r_168__63_ <= r_n_168__63_;
      r_168__62_ <= r_n_168__62_;
      r_168__61_ <= r_n_168__61_;
      r_168__60_ <= r_n_168__60_;
      r_168__59_ <= r_n_168__59_;
      r_168__58_ <= r_n_168__58_;
      r_168__57_ <= r_n_168__57_;
      r_168__56_ <= r_n_168__56_;
      r_168__55_ <= r_n_168__55_;
      r_168__54_ <= r_n_168__54_;
      r_168__53_ <= r_n_168__53_;
      r_168__52_ <= r_n_168__52_;
      r_168__51_ <= r_n_168__51_;
      r_168__50_ <= r_n_168__50_;
      r_168__49_ <= r_n_168__49_;
      r_168__48_ <= r_n_168__48_;
      r_168__47_ <= r_n_168__47_;
      r_168__46_ <= r_n_168__46_;
      r_168__45_ <= r_n_168__45_;
      r_168__44_ <= r_n_168__44_;
      r_168__43_ <= r_n_168__43_;
      r_168__42_ <= r_n_168__42_;
      r_168__41_ <= r_n_168__41_;
      r_168__40_ <= r_n_168__40_;
      r_168__39_ <= r_n_168__39_;
      r_168__38_ <= r_n_168__38_;
      r_168__37_ <= r_n_168__37_;
      r_168__36_ <= r_n_168__36_;
      r_168__35_ <= r_n_168__35_;
      r_168__34_ <= r_n_168__34_;
      r_168__33_ <= r_n_168__33_;
      r_168__32_ <= r_n_168__32_;
      r_168__31_ <= r_n_168__31_;
      r_168__30_ <= r_n_168__30_;
      r_168__29_ <= r_n_168__29_;
      r_168__28_ <= r_n_168__28_;
      r_168__27_ <= r_n_168__27_;
      r_168__26_ <= r_n_168__26_;
      r_168__25_ <= r_n_168__25_;
      r_168__24_ <= r_n_168__24_;
      r_168__23_ <= r_n_168__23_;
      r_168__22_ <= r_n_168__22_;
      r_168__21_ <= r_n_168__21_;
      r_168__20_ <= r_n_168__20_;
      r_168__19_ <= r_n_168__19_;
      r_168__18_ <= r_n_168__18_;
      r_168__17_ <= r_n_168__17_;
      r_168__16_ <= r_n_168__16_;
      r_168__15_ <= r_n_168__15_;
      r_168__14_ <= r_n_168__14_;
      r_168__13_ <= r_n_168__13_;
      r_168__12_ <= r_n_168__12_;
      r_168__11_ <= r_n_168__11_;
      r_168__10_ <= r_n_168__10_;
      r_168__9_ <= r_n_168__9_;
      r_168__8_ <= r_n_168__8_;
      r_168__7_ <= r_n_168__7_;
      r_168__6_ <= r_n_168__6_;
      r_168__5_ <= r_n_168__5_;
      r_168__4_ <= r_n_168__4_;
      r_168__3_ <= r_n_168__3_;
      r_168__2_ <= r_n_168__2_;
      r_168__1_ <= r_n_168__1_;
      r_168__0_ <= r_n_168__0_;
    end 
    if(N3753) begin
      r_169__63_ <= r_n_169__63_;
      r_169__62_ <= r_n_169__62_;
      r_169__61_ <= r_n_169__61_;
      r_169__60_ <= r_n_169__60_;
      r_169__59_ <= r_n_169__59_;
      r_169__58_ <= r_n_169__58_;
      r_169__57_ <= r_n_169__57_;
      r_169__56_ <= r_n_169__56_;
      r_169__55_ <= r_n_169__55_;
      r_169__54_ <= r_n_169__54_;
      r_169__53_ <= r_n_169__53_;
      r_169__52_ <= r_n_169__52_;
      r_169__51_ <= r_n_169__51_;
      r_169__50_ <= r_n_169__50_;
      r_169__49_ <= r_n_169__49_;
      r_169__48_ <= r_n_169__48_;
      r_169__47_ <= r_n_169__47_;
      r_169__46_ <= r_n_169__46_;
      r_169__45_ <= r_n_169__45_;
      r_169__44_ <= r_n_169__44_;
      r_169__43_ <= r_n_169__43_;
      r_169__42_ <= r_n_169__42_;
      r_169__41_ <= r_n_169__41_;
      r_169__40_ <= r_n_169__40_;
      r_169__39_ <= r_n_169__39_;
      r_169__38_ <= r_n_169__38_;
      r_169__37_ <= r_n_169__37_;
      r_169__36_ <= r_n_169__36_;
      r_169__35_ <= r_n_169__35_;
      r_169__34_ <= r_n_169__34_;
      r_169__33_ <= r_n_169__33_;
      r_169__32_ <= r_n_169__32_;
      r_169__31_ <= r_n_169__31_;
      r_169__30_ <= r_n_169__30_;
      r_169__29_ <= r_n_169__29_;
      r_169__28_ <= r_n_169__28_;
      r_169__27_ <= r_n_169__27_;
      r_169__26_ <= r_n_169__26_;
      r_169__25_ <= r_n_169__25_;
      r_169__24_ <= r_n_169__24_;
      r_169__23_ <= r_n_169__23_;
      r_169__22_ <= r_n_169__22_;
      r_169__21_ <= r_n_169__21_;
      r_169__20_ <= r_n_169__20_;
      r_169__19_ <= r_n_169__19_;
      r_169__18_ <= r_n_169__18_;
      r_169__17_ <= r_n_169__17_;
      r_169__16_ <= r_n_169__16_;
      r_169__15_ <= r_n_169__15_;
      r_169__14_ <= r_n_169__14_;
      r_169__13_ <= r_n_169__13_;
      r_169__12_ <= r_n_169__12_;
      r_169__11_ <= r_n_169__11_;
      r_169__10_ <= r_n_169__10_;
      r_169__9_ <= r_n_169__9_;
      r_169__8_ <= r_n_169__8_;
      r_169__7_ <= r_n_169__7_;
      r_169__6_ <= r_n_169__6_;
      r_169__5_ <= r_n_169__5_;
      r_169__4_ <= r_n_169__4_;
      r_169__3_ <= r_n_169__3_;
      r_169__2_ <= r_n_169__2_;
      r_169__1_ <= r_n_169__1_;
      r_169__0_ <= r_n_169__0_;
    end 
    if(N3754) begin
      r_170__63_ <= r_n_170__63_;
      r_170__62_ <= r_n_170__62_;
      r_170__61_ <= r_n_170__61_;
      r_170__60_ <= r_n_170__60_;
      r_170__59_ <= r_n_170__59_;
      r_170__58_ <= r_n_170__58_;
      r_170__57_ <= r_n_170__57_;
      r_170__56_ <= r_n_170__56_;
      r_170__55_ <= r_n_170__55_;
      r_170__54_ <= r_n_170__54_;
      r_170__53_ <= r_n_170__53_;
      r_170__52_ <= r_n_170__52_;
      r_170__51_ <= r_n_170__51_;
      r_170__50_ <= r_n_170__50_;
      r_170__49_ <= r_n_170__49_;
      r_170__48_ <= r_n_170__48_;
      r_170__47_ <= r_n_170__47_;
      r_170__46_ <= r_n_170__46_;
      r_170__45_ <= r_n_170__45_;
      r_170__44_ <= r_n_170__44_;
      r_170__43_ <= r_n_170__43_;
      r_170__42_ <= r_n_170__42_;
      r_170__41_ <= r_n_170__41_;
      r_170__40_ <= r_n_170__40_;
      r_170__39_ <= r_n_170__39_;
      r_170__38_ <= r_n_170__38_;
      r_170__37_ <= r_n_170__37_;
      r_170__36_ <= r_n_170__36_;
      r_170__35_ <= r_n_170__35_;
      r_170__34_ <= r_n_170__34_;
      r_170__33_ <= r_n_170__33_;
      r_170__32_ <= r_n_170__32_;
      r_170__31_ <= r_n_170__31_;
      r_170__30_ <= r_n_170__30_;
      r_170__29_ <= r_n_170__29_;
      r_170__28_ <= r_n_170__28_;
      r_170__27_ <= r_n_170__27_;
      r_170__26_ <= r_n_170__26_;
      r_170__25_ <= r_n_170__25_;
      r_170__24_ <= r_n_170__24_;
      r_170__23_ <= r_n_170__23_;
      r_170__22_ <= r_n_170__22_;
      r_170__21_ <= r_n_170__21_;
      r_170__20_ <= r_n_170__20_;
      r_170__19_ <= r_n_170__19_;
      r_170__18_ <= r_n_170__18_;
      r_170__17_ <= r_n_170__17_;
      r_170__16_ <= r_n_170__16_;
      r_170__15_ <= r_n_170__15_;
      r_170__14_ <= r_n_170__14_;
      r_170__13_ <= r_n_170__13_;
      r_170__12_ <= r_n_170__12_;
      r_170__11_ <= r_n_170__11_;
      r_170__10_ <= r_n_170__10_;
      r_170__9_ <= r_n_170__9_;
      r_170__8_ <= r_n_170__8_;
      r_170__7_ <= r_n_170__7_;
      r_170__6_ <= r_n_170__6_;
      r_170__5_ <= r_n_170__5_;
      r_170__4_ <= r_n_170__4_;
      r_170__3_ <= r_n_170__3_;
      r_170__2_ <= r_n_170__2_;
      r_170__1_ <= r_n_170__1_;
      r_170__0_ <= r_n_170__0_;
    end 
    if(N3755) begin
      r_171__63_ <= r_n_171__63_;
      r_171__62_ <= r_n_171__62_;
      r_171__61_ <= r_n_171__61_;
      r_171__60_ <= r_n_171__60_;
      r_171__59_ <= r_n_171__59_;
      r_171__58_ <= r_n_171__58_;
      r_171__57_ <= r_n_171__57_;
      r_171__56_ <= r_n_171__56_;
      r_171__55_ <= r_n_171__55_;
      r_171__54_ <= r_n_171__54_;
      r_171__53_ <= r_n_171__53_;
      r_171__52_ <= r_n_171__52_;
      r_171__51_ <= r_n_171__51_;
      r_171__50_ <= r_n_171__50_;
      r_171__49_ <= r_n_171__49_;
      r_171__48_ <= r_n_171__48_;
      r_171__47_ <= r_n_171__47_;
      r_171__46_ <= r_n_171__46_;
      r_171__45_ <= r_n_171__45_;
      r_171__44_ <= r_n_171__44_;
      r_171__43_ <= r_n_171__43_;
      r_171__42_ <= r_n_171__42_;
      r_171__41_ <= r_n_171__41_;
      r_171__40_ <= r_n_171__40_;
      r_171__39_ <= r_n_171__39_;
      r_171__38_ <= r_n_171__38_;
      r_171__37_ <= r_n_171__37_;
      r_171__36_ <= r_n_171__36_;
      r_171__35_ <= r_n_171__35_;
      r_171__34_ <= r_n_171__34_;
      r_171__33_ <= r_n_171__33_;
      r_171__32_ <= r_n_171__32_;
      r_171__31_ <= r_n_171__31_;
      r_171__30_ <= r_n_171__30_;
      r_171__29_ <= r_n_171__29_;
      r_171__28_ <= r_n_171__28_;
      r_171__27_ <= r_n_171__27_;
      r_171__26_ <= r_n_171__26_;
      r_171__25_ <= r_n_171__25_;
      r_171__24_ <= r_n_171__24_;
      r_171__23_ <= r_n_171__23_;
      r_171__22_ <= r_n_171__22_;
      r_171__21_ <= r_n_171__21_;
      r_171__20_ <= r_n_171__20_;
      r_171__19_ <= r_n_171__19_;
      r_171__18_ <= r_n_171__18_;
      r_171__17_ <= r_n_171__17_;
      r_171__16_ <= r_n_171__16_;
      r_171__15_ <= r_n_171__15_;
      r_171__14_ <= r_n_171__14_;
      r_171__13_ <= r_n_171__13_;
      r_171__12_ <= r_n_171__12_;
      r_171__11_ <= r_n_171__11_;
      r_171__10_ <= r_n_171__10_;
      r_171__9_ <= r_n_171__9_;
      r_171__8_ <= r_n_171__8_;
      r_171__7_ <= r_n_171__7_;
      r_171__6_ <= r_n_171__6_;
      r_171__5_ <= r_n_171__5_;
      r_171__4_ <= r_n_171__4_;
      r_171__3_ <= r_n_171__3_;
      r_171__2_ <= r_n_171__2_;
      r_171__1_ <= r_n_171__1_;
      r_171__0_ <= r_n_171__0_;
    end 
    if(N3756) begin
      r_172__63_ <= r_n_172__63_;
      r_172__62_ <= r_n_172__62_;
      r_172__61_ <= r_n_172__61_;
      r_172__60_ <= r_n_172__60_;
      r_172__59_ <= r_n_172__59_;
      r_172__58_ <= r_n_172__58_;
      r_172__57_ <= r_n_172__57_;
      r_172__56_ <= r_n_172__56_;
      r_172__55_ <= r_n_172__55_;
      r_172__54_ <= r_n_172__54_;
      r_172__53_ <= r_n_172__53_;
      r_172__52_ <= r_n_172__52_;
      r_172__51_ <= r_n_172__51_;
      r_172__50_ <= r_n_172__50_;
      r_172__49_ <= r_n_172__49_;
      r_172__48_ <= r_n_172__48_;
      r_172__47_ <= r_n_172__47_;
      r_172__46_ <= r_n_172__46_;
      r_172__45_ <= r_n_172__45_;
      r_172__44_ <= r_n_172__44_;
      r_172__43_ <= r_n_172__43_;
      r_172__42_ <= r_n_172__42_;
      r_172__41_ <= r_n_172__41_;
      r_172__40_ <= r_n_172__40_;
      r_172__39_ <= r_n_172__39_;
      r_172__38_ <= r_n_172__38_;
      r_172__37_ <= r_n_172__37_;
      r_172__36_ <= r_n_172__36_;
      r_172__35_ <= r_n_172__35_;
      r_172__34_ <= r_n_172__34_;
      r_172__33_ <= r_n_172__33_;
      r_172__32_ <= r_n_172__32_;
      r_172__31_ <= r_n_172__31_;
      r_172__30_ <= r_n_172__30_;
      r_172__29_ <= r_n_172__29_;
      r_172__28_ <= r_n_172__28_;
      r_172__27_ <= r_n_172__27_;
      r_172__26_ <= r_n_172__26_;
      r_172__25_ <= r_n_172__25_;
      r_172__24_ <= r_n_172__24_;
      r_172__23_ <= r_n_172__23_;
      r_172__22_ <= r_n_172__22_;
      r_172__21_ <= r_n_172__21_;
      r_172__20_ <= r_n_172__20_;
      r_172__19_ <= r_n_172__19_;
      r_172__18_ <= r_n_172__18_;
      r_172__17_ <= r_n_172__17_;
      r_172__16_ <= r_n_172__16_;
      r_172__15_ <= r_n_172__15_;
      r_172__14_ <= r_n_172__14_;
      r_172__13_ <= r_n_172__13_;
      r_172__12_ <= r_n_172__12_;
      r_172__11_ <= r_n_172__11_;
      r_172__10_ <= r_n_172__10_;
      r_172__9_ <= r_n_172__9_;
      r_172__8_ <= r_n_172__8_;
      r_172__7_ <= r_n_172__7_;
      r_172__6_ <= r_n_172__6_;
      r_172__5_ <= r_n_172__5_;
      r_172__4_ <= r_n_172__4_;
      r_172__3_ <= r_n_172__3_;
      r_172__2_ <= r_n_172__2_;
      r_172__1_ <= r_n_172__1_;
      r_172__0_ <= r_n_172__0_;
    end 
    if(N3757) begin
      r_173__63_ <= r_n_173__63_;
      r_173__62_ <= r_n_173__62_;
      r_173__61_ <= r_n_173__61_;
      r_173__60_ <= r_n_173__60_;
      r_173__59_ <= r_n_173__59_;
      r_173__58_ <= r_n_173__58_;
      r_173__57_ <= r_n_173__57_;
      r_173__56_ <= r_n_173__56_;
      r_173__55_ <= r_n_173__55_;
      r_173__54_ <= r_n_173__54_;
      r_173__53_ <= r_n_173__53_;
      r_173__52_ <= r_n_173__52_;
      r_173__51_ <= r_n_173__51_;
      r_173__50_ <= r_n_173__50_;
      r_173__49_ <= r_n_173__49_;
      r_173__48_ <= r_n_173__48_;
      r_173__47_ <= r_n_173__47_;
      r_173__46_ <= r_n_173__46_;
      r_173__45_ <= r_n_173__45_;
      r_173__44_ <= r_n_173__44_;
      r_173__43_ <= r_n_173__43_;
      r_173__42_ <= r_n_173__42_;
      r_173__41_ <= r_n_173__41_;
      r_173__40_ <= r_n_173__40_;
      r_173__39_ <= r_n_173__39_;
      r_173__38_ <= r_n_173__38_;
      r_173__37_ <= r_n_173__37_;
      r_173__36_ <= r_n_173__36_;
      r_173__35_ <= r_n_173__35_;
      r_173__34_ <= r_n_173__34_;
      r_173__33_ <= r_n_173__33_;
      r_173__32_ <= r_n_173__32_;
      r_173__31_ <= r_n_173__31_;
      r_173__30_ <= r_n_173__30_;
      r_173__29_ <= r_n_173__29_;
      r_173__28_ <= r_n_173__28_;
      r_173__27_ <= r_n_173__27_;
      r_173__26_ <= r_n_173__26_;
      r_173__25_ <= r_n_173__25_;
      r_173__24_ <= r_n_173__24_;
      r_173__23_ <= r_n_173__23_;
      r_173__22_ <= r_n_173__22_;
      r_173__21_ <= r_n_173__21_;
      r_173__20_ <= r_n_173__20_;
      r_173__19_ <= r_n_173__19_;
      r_173__18_ <= r_n_173__18_;
      r_173__17_ <= r_n_173__17_;
      r_173__16_ <= r_n_173__16_;
      r_173__15_ <= r_n_173__15_;
      r_173__14_ <= r_n_173__14_;
      r_173__13_ <= r_n_173__13_;
      r_173__12_ <= r_n_173__12_;
      r_173__11_ <= r_n_173__11_;
      r_173__10_ <= r_n_173__10_;
      r_173__9_ <= r_n_173__9_;
      r_173__8_ <= r_n_173__8_;
      r_173__7_ <= r_n_173__7_;
      r_173__6_ <= r_n_173__6_;
      r_173__5_ <= r_n_173__5_;
      r_173__4_ <= r_n_173__4_;
      r_173__3_ <= r_n_173__3_;
      r_173__2_ <= r_n_173__2_;
      r_173__1_ <= r_n_173__1_;
      r_173__0_ <= r_n_173__0_;
    end 
    if(N3758) begin
      r_174__63_ <= r_n_174__63_;
      r_174__62_ <= r_n_174__62_;
      r_174__61_ <= r_n_174__61_;
      r_174__60_ <= r_n_174__60_;
      r_174__59_ <= r_n_174__59_;
      r_174__58_ <= r_n_174__58_;
      r_174__57_ <= r_n_174__57_;
      r_174__56_ <= r_n_174__56_;
      r_174__55_ <= r_n_174__55_;
      r_174__54_ <= r_n_174__54_;
      r_174__53_ <= r_n_174__53_;
      r_174__52_ <= r_n_174__52_;
      r_174__51_ <= r_n_174__51_;
      r_174__50_ <= r_n_174__50_;
      r_174__49_ <= r_n_174__49_;
      r_174__48_ <= r_n_174__48_;
      r_174__47_ <= r_n_174__47_;
      r_174__46_ <= r_n_174__46_;
      r_174__45_ <= r_n_174__45_;
      r_174__44_ <= r_n_174__44_;
      r_174__43_ <= r_n_174__43_;
      r_174__42_ <= r_n_174__42_;
      r_174__41_ <= r_n_174__41_;
      r_174__40_ <= r_n_174__40_;
      r_174__39_ <= r_n_174__39_;
      r_174__38_ <= r_n_174__38_;
      r_174__37_ <= r_n_174__37_;
      r_174__36_ <= r_n_174__36_;
      r_174__35_ <= r_n_174__35_;
      r_174__34_ <= r_n_174__34_;
      r_174__33_ <= r_n_174__33_;
      r_174__32_ <= r_n_174__32_;
      r_174__31_ <= r_n_174__31_;
      r_174__30_ <= r_n_174__30_;
      r_174__29_ <= r_n_174__29_;
      r_174__28_ <= r_n_174__28_;
      r_174__27_ <= r_n_174__27_;
      r_174__26_ <= r_n_174__26_;
      r_174__25_ <= r_n_174__25_;
      r_174__24_ <= r_n_174__24_;
      r_174__23_ <= r_n_174__23_;
      r_174__22_ <= r_n_174__22_;
      r_174__21_ <= r_n_174__21_;
      r_174__20_ <= r_n_174__20_;
      r_174__19_ <= r_n_174__19_;
      r_174__18_ <= r_n_174__18_;
      r_174__17_ <= r_n_174__17_;
      r_174__16_ <= r_n_174__16_;
      r_174__15_ <= r_n_174__15_;
      r_174__14_ <= r_n_174__14_;
      r_174__13_ <= r_n_174__13_;
      r_174__12_ <= r_n_174__12_;
      r_174__11_ <= r_n_174__11_;
      r_174__10_ <= r_n_174__10_;
      r_174__9_ <= r_n_174__9_;
      r_174__8_ <= r_n_174__8_;
      r_174__7_ <= r_n_174__7_;
      r_174__6_ <= r_n_174__6_;
      r_174__5_ <= r_n_174__5_;
      r_174__4_ <= r_n_174__4_;
      r_174__3_ <= r_n_174__3_;
      r_174__2_ <= r_n_174__2_;
      r_174__1_ <= r_n_174__1_;
      r_174__0_ <= r_n_174__0_;
    end 
    if(N3759) begin
      r_175__63_ <= r_n_175__63_;
      r_175__62_ <= r_n_175__62_;
      r_175__61_ <= r_n_175__61_;
      r_175__60_ <= r_n_175__60_;
      r_175__59_ <= r_n_175__59_;
      r_175__58_ <= r_n_175__58_;
      r_175__57_ <= r_n_175__57_;
      r_175__56_ <= r_n_175__56_;
      r_175__55_ <= r_n_175__55_;
      r_175__54_ <= r_n_175__54_;
      r_175__53_ <= r_n_175__53_;
      r_175__52_ <= r_n_175__52_;
      r_175__51_ <= r_n_175__51_;
      r_175__50_ <= r_n_175__50_;
      r_175__49_ <= r_n_175__49_;
      r_175__48_ <= r_n_175__48_;
      r_175__47_ <= r_n_175__47_;
      r_175__46_ <= r_n_175__46_;
      r_175__45_ <= r_n_175__45_;
      r_175__44_ <= r_n_175__44_;
      r_175__43_ <= r_n_175__43_;
      r_175__42_ <= r_n_175__42_;
      r_175__41_ <= r_n_175__41_;
      r_175__40_ <= r_n_175__40_;
      r_175__39_ <= r_n_175__39_;
      r_175__38_ <= r_n_175__38_;
      r_175__37_ <= r_n_175__37_;
      r_175__36_ <= r_n_175__36_;
      r_175__35_ <= r_n_175__35_;
      r_175__34_ <= r_n_175__34_;
      r_175__33_ <= r_n_175__33_;
      r_175__32_ <= r_n_175__32_;
      r_175__31_ <= r_n_175__31_;
      r_175__30_ <= r_n_175__30_;
      r_175__29_ <= r_n_175__29_;
      r_175__28_ <= r_n_175__28_;
      r_175__27_ <= r_n_175__27_;
      r_175__26_ <= r_n_175__26_;
      r_175__25_ <= r_n_175__25_;
      r_175__24_ <= r_n_175__24_;
      r_175__23_ <= r_n_175__23_;
      r_175__22_ <= r_n_175__22_;
      r_175__21_ <= r_n_175__21_;
      r_175__20_ <= r_n_175__20_;
      r_175__19_ <= r_n_175__19_;
      r_175__18_ <= r_n_175__18_;
      r_175__17_ <= r_n_175__17_;
      r_175__16_ <= r_n_175__16_;
      r_175__15_ <= r_n_175__15_;
      r_175__14_ <= r_n_175__14_;
      r_175__13_ <= r_n_175__13_;
      r_175__12_ <= r_n_175__12_;
      r_175__11_ <= r_n_175__11_;
      r_175__10_ <= r_n_175__10_;
      r_175__9_ <= r_n_175__9_;
      r_175__8_ <= r_n_175__8_;
      r_175__7_ <= r_n_175__7_;
      r_175__6_ <= r_n_175__6_;
      r_175__5_ <= r_n_175__5_;
      r_175__4_ <= r_n_175__4_;
      r_175__3_ <= r_n_175__3_;
      r_175__2_ <= r_n_175__2_;
      r_175__1_ <= r_n_175__1_;
      r_175__0_ <= r_n_175__0_;
    end 
    if(N3760) begin
      r_176__63_ <= r_n_176__63_;
      r_176__62_ <= r_n_176__62_;
      r_176__61_ <= r_n_176__61_;
      r_176__60_ <= r_n_176__60_;
      r_176__59_ <= r_n_176__59_;
      r_176__58_ <= r_n_176__58_;
      r_176__57_ <= r_n_176__57_;
      r_176__56_ <= r_n_176__56_;
      r_176__55_ <= r_n_176__55_;
      r_176__54_ <= r_n_176__54_;
      r_176__53_ <= r_n_176__53_;
      r_176__52_ <= r_n_176__52_;
      r_176__51_ <= r_n_176__51_;
      r_176__50_ <= r_n_176__50_;
      r_176__49_ <= r_n_176__49_;
      r_176__48_ <= r_n_176__48_;
      r_176__47_ <= r_n_176__47_;
      r_176__46_ <= r_n_176__46_;
      r_176__45_ <= r_n_176__45_;
      r_176__44_ <= r_n_176__44_;
      r_176__43_ <= r_n_176__43_;
      r_176__42_ <= r_n_176__42_;
      r_176__41_ <= r_n_176__41_;
      r_176__40_ <= r_n_176__40_;
      r_176__39_ <= r_n_176__39_;
      r_176__38_ <= r_n_176__38_;
      r_176__37_ <= r_n_176__37_;
      r_176__36_ <= r_n_176__36_;
      r_176__35_ <= r_n_176__35_;
      r_176__34_ <= r_n_176__34_;
      r_176__33_ <= r_n_176__33_;
      r_176__32_ <= r_n_176__32_;
      r_176__31_ <= r_n_176__31_;
      r_176__30_ <= r_n_176__30_;
      r_176__29_ <= r_n_176__29_;
      r_176__28_ <= r_n_176__28_;
      r_176__27_ <= r_n_176__27_;
      r_176__26_ <= r_n_176__26_;
      r_176__25_ <= r_n_176__25_;
      r_176__24_ <= r_n_176__24_;
      r_176__23_ <= r_n_176__23_;
      r_176__22_ <= r_n_176__22_;
      r_176__21_ <= r_n_176__21_;
      r_176__20_ <= r_n_176__20_;
      r_176__19_ <= r_n_176__19_;
      r_176__18_ <= r_n_176__18_;
      r_176__17_ <= r_n_176__17_;
      r_176__16_ <= r_n_176__16_;
      r_176__15_ <= r_n_176__15_;
      r_176__14_ <= r_n_176__14_;
      r_176__13_ <= r_n_176__13_;
      r_176__12_ <= r_n_176__12_;
      r_176__11_ <= r_n_176__11_;
      r_176__10_ <= r_n_176__10_;
      r_176__9_ <= r_n_176__9_;
      r_176__8_ <= r_n_176__8_;
      r_176__7_ <= r_n_176__7_;
      r_176__6_ <= r_n_176__6_;
      r_176__5_ <= r_n_176__5_;
      r_176__4_ <= r_n_176__4_;
      r_176__3_ <= r_n_176__3_;
      r_176__2_ <= r_n_176__2_;
      r_176__1_ <= r_n_176__1_;
      r_176__0_ <= r_n_176__0_;
    end 
    if(N3761) begin
      r_177__63_ <= r_n_177__63_;
      r_177__62_ <= r_n_177__62_;
      r_177__61_ <= r_n_177__61_;
      r_177__60_ <= r_n_177__60_;
      r_177__59_ <= r_n_177__59_;
      r_177__58_ <= r_n_177__58_;
      r_177__57_ <= r_n_177__57_;
      r_177__56_ <= r_n_177__56_;
      r_177__55_ <= r_n_177__55_;
      r_177__54_ <= r_n_177__54_;
      r_177__53_ <= r_n_177__53_;
      r_177__52_ <= r_n_177__52_;
      r_177__51_ <= r_n_177__51_;
      r_177__50_ <= r_n_177__50_;
      r_177__49_ <= r_n_177__49_;
      r_177__48_ <= r_n_177__48_;
      r_177__47_ <= r_n_177__47_;
      r_177__46_ <= r_n_177__46_;
      r_177__45_ <= r_n_177__45_;
      r_177__44_ <= r_n_177__44_;
      r_177__43_ <= r_n_177__43_;
      r_177__42_ <= r_n_177__42_;
      r_177__41_ <= r_n_177__41_;
      r_177__40_ <= r_n_177__40_;
      r_177__39_ <= r_n_177__39_;
      r_177__38_ <= r_n_177__38_;
      r_177__37_ <= r_n_177__37_;
      r_177__36_ <= r_n_177__36_;
      r_177__35_ <= r_n_177__35_;
      r_177__34_ <= r_n_177__34_;
      r_177__33_ <= r_n_177__33_;
      r_177__32_ <= r_n_177__32_;
      r_177__31_ <= r_n_177__31_;
      r_177__30_ <= r_n_177__30_;
      r_177__29_ <= r_n_177__29_;
      r_177__28_ <= r_n_177__28_;
      r_177__27_ <= r_n_177__27_;
      r_177__26_ <= r_n_177__26_;
      r_177__25_ <= r_n_177__25_;
      r_177__24_ <= r_n_177__24_;
      r_177__23_ <= r_n_177__23_;
      r_177__22_ <= r_n_177__22_;
      r_177__21_ <= r_n_177__21_;
      r_177__20_ <= r_n_177__20_;
      r_177__19_ <= r_n_177__19_;
      r_177__18_ <= r_n_177__18_;
      r_177__17_ <= r_n_177__17_;
      r_177__16_ <= r_n_177__16_;
      r_177__15_ <= r_n_177__15_;
      r_177__14_ <= r_n_177__14_;
      r_177__13_ <= r_n_177__13_;
      r_177__12_ <= r_n_177__12_;
      r_177__11_ <= r_n_177__11_;
      r_177__10_ <= r_n_177__10_;
      r_177__9_ <= r_n_177__9_;
      r_177__8_ <= r_n_177__8_;
      r_177__7_ <= r_n_177__7_;
      r_177__6_ <= r_n_177__6_;
      r_177__5_ <= r_n_177__5_;
      r_177__4_ <= r_n_177__4_;
      r_177__3_ <= r_n_177__3_;
      r_177__2_ <= r_n_177__2_;
      r_177__1_ <= r_n_177__1_;
      r_177__0_ <= r_n_177__0_;
    end 
    if(N3762) begin
      r_178__63_ <= r_n_178__63_;
      r_178__62_ <= r_n_178__62_;
      r_178__61_ <= r_n_178__61_;
      r_178__60_ <= r_n_178__60_;
      r_178__59_ <= r_n_178__59_;
      r_178__58_ <= r_n_178__58_;
      r_178__57_ <= r_n_178__57_;
      r_178__56_ <= r_n_178__56_;
      r_178__55_ <= r_n_178__55_;
      r_178__54_ <= r_n_178__54_;
      r_178__53_ <= r_n_178__53_;
      r_178__52_ <= r_n_178__52_;
      r_178__51_ <= r_n_178__51_;
      r_178__50_ <= r_n_178__50_;
      r_178__49_ <= r_n_178__49_;
      r_178__48_ <= r_n_178__48_;
      r_178__47_ <= r_n_178__47_;
      r_178__46_ <= r_n_178__46_;
      r_178__45_ <= r_n_178__45_;
      r_178__44_ <= r_n_178__44_;
      r_178__43_ <= r_n_178__43_;
      r_178__42_ <= r_n_178__42_;
      r_178__41_ <= r_n_178__41_;
      r_178__40_ <= r_n_178__40_;
      r_178__39_ <= r_n_178__39_;
      r_178__38_ <= r_n_178__38_;
      r_178__37_ <= r_n_178__37_;
      r_178__36_ <= r_n_178__36_;
      r_178__35_ <= r_n_178__35_;
      r_178__34_ <= r_n_178__34_;
      r_178__33_ <= r_n_178__33_;
      r_178__32_ <= r_n_178__32_;
      r_178__31_ <= r_n_178__31_;
      r_178__30_ <= r_n_178__30_;
      r_178__29_ <= r_n_178__29_;
      r_178__28_ <= r_n_178__28_;
      r_178__27_ <= r_n_178__27_;
      r_178__26_ <= r_n_178__26_;
      r_178__25_ <= r_n_178__25_;
      r_178__24_ <= r_n_178__24_;
      r_178__23_ <= r_n_178__23_;
      r_178__22_ <= r_n_178__22_;
      r_178__21_ <= r_n_178__21_;
      r_178__20_ <= r_n_178__20_;
      r_178__19_ <= r_n_178__19_;
      r_178__18_ <= r_n_178__18_;
      r_178__17_ <= r_n_178__17_;
      r_178__16_ <= r_n_178__16_;
      r_178__15_ <= r_n_178__15_;
      r_178__14_ <= r_n_178__14_;
      r_178__13_ <= r_n_178__13_;
      r_178__12_ <= r_n_178__12_;
      r_178__11_ <= r_n_178__11_;
      r_178__10_ <= r_n_178__10_;
      r_178__9_ <= r_n_178__9_;
      r_178__8_ <= r_n_178__8_;
      r_178__7_ <= r_n_178__7_;
      r_178__6_ <= r_n_178__6_;
      r_178__5_ <= r_n_178__5_;
      r_178__4_ <= r_n_178__4_;
      r_178__3_ <= r_n_178__3_;
      r_178__2_ <= r_n_178__2_;
      r_178__1_ <= r_n_178__1_;
      r_178__0_ <= r_n_178__0_;
    end 
    if(N3763) begin
      r_179__63_ <= r_n_179__63_;
      r_179__62_ <= r_n_179__62_;
      r_179__61_ <= r_n_179__61_;
      r_179__60_ <= r_n_179__60_;
      r_179__59_ <= r_n_179__59_;
      r_179__58_ <= r_n_179__58_;
      r_179__57_ <= r_n_179__57_;
      r_179__56_ <= r_n_179__56_;
      r_179__55_ <= r_n_179__55_;
      r_179__54_ <= r_n_179__54_;
      r_179__53_ <= r_n_179__53_;
      r_179__52_ <= r_n_179__52_;
      r_179__51_ <= r_n_179__51_;
      r_179__50_ <= r_n_179__50_;
      r_179__49_ <= r_n_179__49_;
      r_179__48_ <= r_n_179__48_;
      r_179__47_ <= r_n_179__47_;
      r_179__46_ <= r_n_179__46_;
      r_179__45_ <= r_n_179__45_;
      r_179__44_ <= r_n_179__44_;
      r_179__43_ <= r_n_179__43_;
      r_179__42_ <= r_n_179__42_;
      r_179__41_ <= r_n_179__41_;
      r_179__40_ <= r_n_179__40_;
      r_179__39_ <= r_n_179__39_;
      r_179__38_ <= r_n_179__38_;
      r_179__37_ <= r_n_179__37_;
      r_179__36_ <= r_n_179__36_;
      r_179__35_ <= r_n_179__35_;
      r_179__34_ <= r_n_179__34_;
      r_179__33_ <= r_n_179__33_;
      r_179__32_ <= r_n_179__32_;
      r_179__31_ <= r_n_179__31_;
      r_179__30_ <= r_n_179__30_;
      r_179__29_ <= r_n_179__29_;
      r_179__28_ <= r_n_179__28_;
      r_179__27_ <= r_n_179__27_;
      r_179__26_ <= r_n_179__26_;
      r_179__25_ <= r_n_179__25_;
      r_179__24_ <= r_n_179__24_;
      r_179__23_ <= r_n_179__23_;
      r_179__22_ <= r_n_179__22_;
      r_179__21_ <= r_n_179__21_;
      r_179__20_ <= r_n_179__20_;
      r_179__19_ <= r_n_179__19_;
      r_179__18_ <= r_n_179__18_;
      r_179__17_ <= r_n_179__17_;
      r_179__16_ <= r_n_179__16_;
      r_179__15_ <= r_n_179__15_;
      r_179__14_ <= r_n_179__14_;
      r_179__13_ <= r_n_179__13_;
      r_179__12_ <= r_n_179__12_;
      r_179__11_ <= r_n_179__11_;
      r_179__10_ <= r_n_179__10_;
      r_179__9_ <= r_n_179__9_;
      r_179__8_ <= r_n_179__8_;
      r_179__7_ <= r_n_179__7_;
      r_179__6_ <= r_n_179__6_;
      r_179__5_ <= r_n_179__5_;
      r_179__4_ <= r_n_179__4_;
      r_179__3_ <= r_n_179__3_;
      r_179__2_ <= r_n_179__2_;
      r_179__1_ <= r_n_179__1_;
      r_179__0_ <= r_n_179__0_;
    end 
    if(N3764) begin
      r_180__63_ <= r_n_180__63_;
      r_180__62_ <= r_n_180__62_;
      r_180__61_ <= r_n_180__61_;
      r_180__60_ <= r_n_180__60_;
      r_180__59_ <= r_n_180__59_;
      r_180__58_ <= r_n_180__58_;
      r_180__57_ <= r_n_180__57_;
      r_180__56_ <= r_n_180__56_;
      r_180__55_ <= r_n_180__55_;
      r_180__54_ <= r_n_180__54_;
      r_180__53_ <= r_n_180__53_;
      r_180__52_ <= r_n_180__52_;
      r_180__51_ <= r_n_180__51_;
      r_180__50_ <= r_n_180__50_;
      r_180__49_ <= r_n_180__49_;
      r_180__48_ <= r_n_180__48_;
      r_180__47_ <= r_n_180__47_;
      r_180__46_ <= r_n_180__46_;
      r_180__45_ <= r_n_180__45_;
      r_180__44_ <= r_n_180__44_;
      r_180__43_ <= r_n_180__43_;
      r_180__42_ <= r_n_180__42_;
      r_180__41_ <= r_n_180__41_;
      r_180__40_ <= r_n_180__40_;
      r_180__39_ <= r_n_180__39_;
      r_180__38_ <= r_n_180__38_;
      r_180__37_ <= r_n_180__37_;
      r_180__36_ <= r_n_180__36_;
      r_180__35_ <= r_n_180__35_;
      r_180__34_ <= r_n_180__34_;
      r_180__33_ <= r_n_180__33_;
      r_180__32_ <= r_n_180__32_;
      r_180__31_ <= r_n_180__31_;
      r_180__30_ <= r_n_180__30_;
      r_180__29_ <= r_n_180__29_;
      r_180__28_ <= r_n_180__28_;
      r_180__27_ <= r_n_180__27_;
      r_180__26_ <= r_n_180__26_;
      r_180__25_ <= r_n_180__25_;
      r_180__24_ <= r_n_180__24_;
      r_180__23_ <= r_n_180__23_;
      r_180__22_ <= r_n_180__22_;
      r_180__21_ <= r_n_180__21_;
      r_180__20_ <= r_n_180__20_;
      r_180__19_ <= r_n_180__19_;
      r_180__18_ <= r_n_180__18_;
      r_180__17_ <= r_n_180__17_;
      r_180__16_ <= r_n_180__16_;
      r_180__15_ <= r_n_180__15_;
      r_180__14_ <= r_n_180__14_;
      r_180__13_ <= r_n_180__13_;
      r_180__12_ <= r_n_180__12_;
      r_180__11_ <= r_n_180__11_;
      r_180__10_ <= r_n_180__10_;
      r_180__9_ <= r_n_180__9_;
      r_180__8_ <= r_n_180__8_;
      r_180__7_ <= r_n_180__7_;
      r_180__6_ <= r_n_180__6_;
      r_180__5_ <= r_n_180__5_;
      r_180__4_ <= r_n_180__4_;
      r_180__3_ <= r_n_180__3_;
      r_180__2_ <= r_n_180__2_;
      r_180__1_ <= r_n_180__1_;
      r_180__0_ <= r_n_180__0_;
    end 
    if(N3765) begin
      r_181__63_ <= r_n_181__63_;
      r_181__62_ <= r_n_181__62_;
      r_181__61_ <= r_n_181__61_;
      r_181__60_ <= r_n_181__60_;
      r_181__59_ <= r_n_181__59_;
      r_181__58_ <= r_n_181__58_;
      r_181__57_ <= r_n_181__57_;
      r_181__56_ <= r_n_181__56_;
      r_181__55_ <= r_n_181__55_;
      r_181__54_ <= r_n_181__54_;
      r_181__53_ <= r_n_181__53_;
      r_181__52_ <= r_n_181__52_;
      r_181__51_ <= r_n_181__51_;
      r_181__50_ <= r_n_181__50_;
      r_181__49_ <= r_n_181__49_;
      r_181__48_ <= r_n_181__48_;
      r_181__47_ <= r_n_181__47_;
      r_181__46_ <= r_n_181__46_;
      r_181__45_ <= r_n_181__45_;
      r_181__44_ <= r_n_181__44_;
      r_181__43_ <= r_n_181__43_;
      r_181__42_ <= r_n_181__42_;
      r_181__41_ <= r_n_181__41_;
      r_181__40_ <= r_n_181__40_;
      r_181__39_ <= r_n_181__39_;
      r_181__38_ <= r_n_181__38_;
      r_181__37_ <= r_n_181__37_;
      r_181__36_ <= r_n_181__36_;
      r_181__35_ <= r_n_181__35_;
      r_181__34_ <= r_n_181__34_;
      r_181__33_ <= r_n_181__33_;
      r_181__32_ <= r_n_181__32_;
      r_181__31_ <= r_n_181__31_;
      r_181__30_ <= r_n_181__30_;
      r_181__29_ <= r_n_181__29_;
      r_181__28_ <= r_n_181__28_;
      r_181__27_ <= r_n_181__27_;
      r_181__26_ <= r_n_181__26_;
      r_181__25_ <= r_n_181__25_;
      r_181__24_ <= r_n_181__24_;
      r_181__23_ <= r_n_181__23_;
      r_181__22_ <= r_n_181__22_;
      r_181__21_ <= r_n_181__21_;
      r_181__20_ <= r_n_181__20_;
      r_181__19_ <= r_n_181__19_;
      r_181__18_ <= r_n_181__18_;
      r_181__17_ <= r_n_181__17_;
      r_181__16_ <= r_n_181__16_;
      r_181__15_ <= r_n_181__15_;
      r_181__14_ <= r_n_181__14_;
      r_181__13_ <= r_n_181__13_;
      r_181__12_ <= r_n_181__12_;
      r_181__11_ <= r_n_181__11_;
      r_181__10_ <= r_n_181__10_;
      r_181__9_ <= r_n_181__9_;
      r_181__8_ <= r_n_181__8_;
      r_181__7_ <= r_n_181__7_;
      r_181__6_ <= r_n_181__6_;
      r_181__5_ <= r_n_181__5_;
      r_181__4_ <= r_n_181__4_;
      r_181__3_ <= r_n_181__3_;
      r_181__2_ <= r_n_181__2_;
      r_181__1_ <= r_n_181__1_;
      r_181__0_ <= r_n_181__0_;
    end 
    if(N3766) begin
      r_182__63_ <= r_n_182__63_;
      r_182__62_ <= r_n_182__62_;
      r_182__61_ <= r_n_182__61_;
      r_182__60_ <= r_n_182__60_;
      r_182__59_ <= r_n_182__59_;
      r_182__58_ <= r_n_182__58_;
      r_182__57_ <= r_n_182__57_;
      r_182__56_ <= r_n_182__56_;
      r_182__55_ <= r_n_182__55_;
      r_182__54_ <= r_n_182__54_;
      r_182__53_ <= r_n_182__53_;
      r_182__52_ <= r_n_182__52_;
      r_182__51_ <= r_n_182__51_;
      r_182__50_ <= r_n_182__50_;
      r_182__49_ <= r_n_182__49_;
      r_182__48_ <= r_n_182__48_;
      r_182__47_ <= r_n_182__47_;
      r_182__46_ <= r_n_182__46_;
      r_182__45_ <= r_n_182__45_;
      r_182__44_ <= r_n_182__44_;
      r_182__43_ <= r_n_182__43_;
      r_182__42_ <= r_n_182__42_;
      r_182__41_ <= r_n_182__41_;
      r_182__40_ <= r_n_182__40_;
      r_182__39_ <= r_n_182__39_;
      r_182__38_ <= r_n_182__38_;
      r_182__37_ <= r_n_182__37_;
      r_182__36_ <= r_n_182__36_;
      r_182__35_ <= r_n_182__35_;
      r_182__34_ <= r_n_182__34_;
      r_182__33_ <= r_n_182__33_;
      r_182__32_ <= r_n_182__32_;
      r_182__31_ <= r_n_182__31_;
      r_182__30_ <= r_n_182__30_;
      r_182__29_ <= r_n_182__29_;
      r_182__28_ <= r_n_182__28_;
      r_182__27_ <= r_n_182__27_;
      r_182__26_ <= r_n_182__26_;
      r_182__25_ <= r_n_182__25_;
      r_182__24_ <= r_n_182__24_;
      r_182__23_ <= r_n_182__23_;
      r_182__22_ <= r_n_182__22_;
      r_182__21_ <= r_n_182__21_;
      r_182__20_ <= r_n_182__20_;
      r_182__19_ <= r_n_182__19_;
      r_182__18_ <= r_n_182__18_;
      r_182__17_ <= r_n_182__17_;
      r_182__16_ <= r_n_182__16_;
      r_182__15_ <= r_n_182__15_;
      r_182__14_ <= r_n_182__14_;
      r_182__13_ <= r_n_182__13_;
      r_182__12_ <= r_n_182__12_;
      r_182__11_ <= r_n_182__11_;
      r_182__10_ <= r_n_182__10_;
      r_182__9_ <= r_n_182__9_;
      r_182__8_ <= r_n_182__8_;
      r_182__7_ <= r_n_182__7_;
      r_182__6_ <= r_n_182__6_;
      r_182__5_ <= r_n_182__5_;
      r_182__4_ <= r_n_182__4_;
      r_182__3_ <= r_n_182__3_;
      r_182__2_ <= r_n_182__2_;
      r_182__1_ <= r_n_182__1_;
      r_182__0_ <= r_n_182__0_;
    end 
    if(N3767) begin
      r_183__63_ <= r_n_183__63_;
      r_183__62_ <= r_n_183__62_;
      r_183__61_ <= r_n_183__61_;
      r_183__60_ <= r_n_183__60_;
      r_183__59_ <= r_n_183__59_;
      r_183__58_ <= r_n_183__58_;
      r_183__57_ <= r_n_183__57_;
      r_183__56_ <= r_n_183__56_;
      r_183__55_ <= r_n_183__55_;
      r_183__54_ <= r_n_183__54_;
      r_183__53_ <= r_n_183__53_;
      r_183__52_ <= r_n_183__52_;
      r_183__51_ <= r_n_183__51_;
      r_183__50_ <= r_n_183__50_;
      r_183__49_ <= r_n_183__49_;
      r_183__48_ <= r_n_183__48_;
      r_183__47_ <= r_n_183__47_;
      r_183__46_ <= r_n_183__46_;
      r_183__45_ <= r_n_183__45_;
      r_183__44_ <= r_n_183__44_;
      r_183__43_ <= r_n_183__43_;
      r_183__42_ <= r_n_183__42_;
      r_183__41_ <= r_n_183__41_;
      r_183__40_ <= r_n_183__40_;
      r_183__39_ <= r_n_183__39_;
      r_183__38_ <= r_n_183__38_;
      r_183__37_ <= r_n_183__37_;
      r_183__36_ <= r_n_183__36_;
      r_183__35_ <= r_n_183__35_;
      r_183__34_ <= r_n_183__34_;
      r_183__33_ <= r_n_183__33_;
      r_183__32_ <= r_n_183__32_;
      r_183__31_ <= r_n_183__31_;
      r_183__30_ <= r_n_183__30_;
      r_183__29_ <= r_n_183__29_;
      r_183__28_ <= r_n_183__28_;
      r_183__27_ <= r_n_183__27_;
      r_183__26_ <= r_n_183__26_;
      r_183__25_ <= r_n_183__25_;
      r_183__24_ <= r_n_183__24_;
      r_183__23_ <= r_n_183__23_;
      r_183__22_ <= r_n_183__22_;
      r_183__21_ <= r_n_183__21_;
      r_183__20_ <= r_n_183__20_;
      r_183__19_ <= r_n_183__19_;
      r_183__18_ <= r_n_183__18_;
      r_183__17_ <= r_n_183__17_;
      r_183__16_ <= r_n_183__16_;
      r_183__15_ <= r_n_183__15_;
      r_183__14_ <= r_n_183__14_;
      r_183__13_ <= r_n_183__13_;
      r_183__12_ <= r_n_183__12_;
      r_183__11_ <= r_n_183__11_;
      r_183__10_ <= r_n_183__10_;
      r_183__9_ <= r_n_183__9_;
      r_183__8_ <= r_n_183__8_;
      r_183__7_ <= r_n_183__7_;
      r_183__6_ <= r_n_183__6_;
      r_183__5_ <= r_n_183__5_;
      r_183__4_ <= r_n_183__4_;
      r_183__3_ <= r_n_183__3_;
      r_183__2_ <= r_n_183__2_;
      r_183__1_ <= r_n_183__1_;
      r_183__0_ <= r_n_183__0_;
    end 
    if(N3768) begin
      r_184__63_ <= r_n_184__63_;
      r_184__62_ <= r_n_184__62_;
      r_184__61_ <= r_n_184__61_;
      r_184__60_ <= r_n_184__60_;
      r_184__59_ <= r_n_184__59_;
      r_184__58_ <= r_n_184__58_;
      r_184__57_ <= r_n_184__57_;
      r_184__56_ <= r_n_184__56_;
      r_184__55_ <= r_n_184__55_;
      r_184__54_ <= r_n_184__54_;
      r_184__53_ <= r_n_184__53_;
      r_184__52_ <= r_n_184__52_;
      r_184__51_ <= r_n_184__51_;
      r_184__50_ <= r_n_184__50_;
      r_184__49_ <= r_n_184__49_;
      r_184__48_ <= r_n_184__48_;
      r_184__47_ <= r_n_184__47_;
      r_184__46_ <= r_n_184__46_;
      r_184__45_ <= r_n_184__45_;
      r_184__44_ <= r_n_184__44_;
      r_184__43_ <= r_n_184__43_;
      r_184__42_ <= r_n_184__42_;
      r_184__41_ <= r_n_184__41_;
      r_184__40_ <= r_n_184__40_;
      r_184__39_ <= r_n_184__39_;
      r_184__38_ <= r_n_184__38_;
      r_184__37_ <= r_n_184__37_;
      r_184__36_ <= r_n_184__36_;
      r_184__35_ <= r_n_184__35_;
      r_184__34_ <= r_n_184__34_;
      r_184__33_ <= r_n_184__33_;
      r_184__32_ <= r_n_184__32_;
      r_184__31_ <= r_n_184__31_;
      r_184__30_ <= r_n_184__30_;
      r_184__29_ <= r_n_184__29_;
      r_184__28_ <= r_n_184__28_;
      r_184__27_ <= r_n_184__27_;
      r_184__26_ <= r_n_184__26_;
      r_184__25_ <= r_n_184__25_;
      r_184__24_ <= r_n_184__24_;
      r_184__23_ <= r_n_184__23_;
      r_184__22_ <= r_n_184__22_;
      r_184__21_ <= r_n_184__21_;
      r_184__20_ <= r_n_184__20_;
      r_184__19_ <= r_n_184__19_;
      r_184__18_ <= r_n_184__18_;
      r_184__17_ <= r_n_184__17_;
      r_184__16_ <= r_n_184__16_;
      r_184__15_ <= r_n_184__15_;
      r_184__14_ <= r_n_184__14_;
      r_184__13_ <= r_n_184__13_;
      r_184__12_ <= r_n_184__12_;
      r_184__11_ <= r_n_184__11_;
      r_184__10_ <= r_n_184__10_;
      r_184__9_ <= r_n_184__9_;
      r_184__8_ <= r_n_184__8_;
      r_184__7_ <= r_n_184__7_;
      r_184__6_ <= r_n_184__6_;
      r_184__5_ <= r_n_184__5_;
      r_184__4_ <= r_n_184__4_;
      r_184__3_ <= r_n_184__3_;
      r_184__2_ <= r_n_184__2_;
      r_184__1_ <= r_n_184__1_;
      r_184__0_ <= r_n_184__0_;
    end 
    if(N3769) begin
      r_185__63_ <= r_n_185__63_;
      r_185__62_ <= r_n_185__62_;
      r_185__61_ <= r_n_185__61_;
      r_185__60_ <= r_n_185__60_;
      r_185__59_ <= r_n_185__59_;
      r_185__58_ <= r_n_185__58_;
      r_185__57_ <= r_n_185__57_;
      r_185__56_ <= r_n_185__56_;
      r_185__55_ <= r_n_185__55_;
      r_185__54_ <= r_n_185__54_;
      r_185__53_ <= r_n_185__53_;
      r_185__52_ <= r_n_185__52_;
      r_185__51_ <= r_n_185__51_;
      r_185__50_ <= r_n_185__50_;
      r_185__49_ <= r_n_185__49_;
      r_185__48_ <= r_n_185__48_;
      r_185__47_ <= r_n_185__47_;
      r_185__46_ <= r_n_185__46_;
      r_185__45_ <= r_n_185__45_;
      r_185__44_ <= r_n_185__44_;
      r_185__43_ <= r_n_185__43_;
      r_185__42_ <= r_n_185__42_;
      r_185__41_ <= r_n_185__41_;
      r_185__40_ <= r_n_185__40_;
      r_185__39_ <= r_n_185__39_;
      r_185__38_ <= r_n_185__38_;
      r_185__37_ <= r_n_185__37_;
      r_185__36_ <= r_n_185__36_;
      r_185__35_ <= r_n_185__35_;
      r_185__34_ <= r_n_185__34_;
      r_185__33_ <= r_n_185__33_;
      r_185__32_ <= r_n_185__32_;
      r_185__31_ <= r_n_185__31_;
      r_185__30_ <= r_n_185__30_;
      r_185__29_ <= r_n_185__29_;
      r_185__28_ <= r_n_185__28_;
      r_185__27_ <= r_n_185__27_;
      r_185__26_ <= r_n_185__26_;
      r_185__25_ <= r_n_185__25_;
      r_185__24_ <= r_n_185__24_;
      r_185__23_ <= r_n_185__23_;
      r_185__22_ <= r_n_185__22_;
      r_185__21_ <= r_n_185__21_;
      r_185__20_ <= r_n_185__20_;
      r_185__19_ <= r_n_185__19_;
      r_185__18_ <= r_n_185__18_;
      r_185__17_ <= r_n_185__17_;
      r_185__16_ <= r_n_185__16_;
      r_185__15_ <= r_n_185__15_;
      r_185__14_ <= r_n_185__14_;
      r_185__13_ <= r_n_185__13_;
      r_185__12_ <= r_n_185__12_;
      r_185__11_ <= r_n_185__11_;
      r_185__10_ <= r_n_185__10_;
      r_185__9_ <= r_n_185__9_;
      r_185__8_ <= r_n_185__8_;
      r_185__7_ <= r_n_185__7_;
      r_185__6_ <= r_n_185__6_;
      r_185__5_ <= r_n_185__5_;
      r_185__4_ <= r_n_185__4_;
      r_185__3_ <= r_n_185__3_;
      r_185__2_ <= r_n_185__2_;
      r_185__1_ <= r_n_185__1_;
      r_185__0_ <= r_n_185__0_;
    end 
    if(N3770) begin
      r_186__63_ <= r_n_186__63_;
      r_186__62_ <= r_n_186__62_;
      r_186__61_ <= r_n_186__61_;
      r_186__60_ <= r_n_186__60_;
      r_186__59_ <= r_n_186__59_;
      r_186__58_ <= r_n_186__58_;
      r_186__57_ <= r_n_186__57_;
      r_186__56_ <= r_n_186__56_;
      r_186__55_ <= r_n_186__55_;
      r_186__54_ <= r_n_186__54_;
      r_186__53_ <= r_n_186__53_;
      r_186__52_ <= r_n_186__52_;
      r_186__51_ <= r_n_186__51_;
      r_186__50_ <= r_n_186__50_;
      r_186__49_ <= r_n_186__49_;
      r_186__48_ <= r_n_186__48_;
      r_186__47_ <= r_n_186__47_;
      r_186__46_ <= r_n_186__46_;
      r_186__45_ <= r_n_186__45_;
      r_186__44_ <= r_n_186__44_;
      r_186__43_ <= r_n_186__43_;
      r_186__42_ <= r_n_186__42_;
      r_186__41_ <= r_n_186__41_;
      r_186__40_ <= r_n_186__40_;
      r_186__39_ <= r_n_186__39_;
      r_186__38_ <= r_n_186__38_;
      r_186__37_ <= r_n_186__37_;
      r_186__36_ <= r_n_186__36_;
      r_186__35_ <= r_n_186__35_;
      r_186__34_ <= r_n_186__34_;
      r_186__33_ <= r_n_186__33_;
      r_186__32_ <= r_n_186__32_;
      r_186__31_ <= r_n_186__31_;
      r_186__30_ <= r_n_186__30_;
      r_186__29_ <= r_n_186__29_;
      r_186__28_ <= r_n_186__28_;
      r_186__27_ <= r_n_186__27_;
      r_186__26_ <= r_n_186__26_;
      r_186__25_ <= r_n_186__25_;
      r_186__24_ <= r_n_186__24_;
      r_186__23_ <= r_n_186__23_;
      r_186__22_ <= r_n_186__22_;
      r_186__21_ <= r_n_186__21_;
      r_186__20_ <= r_n_186__20_;
      r_186__19_ <= r_n_186__19_;
      r_186__18_ <= r_n_186__18_;
      r_186__17_ <= r_n_186__17_;
      r_186__16_ <= r_n_186__16_;
      r_186__15_ <= r_n_186__15_;
      r_186__14_ <= r_n_186__14_;
      r_186__13_ <= r_n_186__13_;
      r_186__12_ <= r_n_186__12_;
      r_186__11_ <= r_n_186__11_;
      r_186__10_ <= r_n_186__10_;
      r_186__9_ <= r_n_186__9_;
      r_186__8_ <= r_n_186__8_;
      r_186__7_ <= r_n_186__7_;
      r_186__6_ <= r_n_186__6_;
      r_186__5_ <= r_n_186__5_;
      r_186__4_ <= r_n_186__4_;
      r_186__3_ <= r_n_186__3_;
      r_186__2_ <= r_n_186__2_;
      r_186__1_ <= r_n_186__1_;
      r_186__0_ <= r_n_186__0_;
    end 
    if(N3771) begin
      r_187__63_ <= r_n_187__63_;
      r_187__62_ <= r_n_187__62_;
      r_187__61_ <= r_n_187__61_;
      r_187__60_ <= r_n_187__60_;
      r_187__59_ <= r_n_187__59_;
      r_187__58_ <= r_n_187__58_;
      r_187__57_ <= r_n_187__57_;
      r_187__56_ <= r_n_187__56_;
      r_187__55_ <= r_n_187__55_;
      r_187__54_ <= r_n_187__54_;
      r_187__53_ <= r_n_187__53_;
      r_187__52_ <= r_n_187__52_;
      r_187__51_ <= r_n_187__51_;
      r_187__50_ <= r_n_187__50_;
      r_187__49_ <= r_n_187__49_;
      r_187__48_ <= r_n_187__48_;
      r_187__47_ <= r_n_187__47_;
      r_187__46_ <= r_n_187__46_;
      r_187__45_ <= r_n_187__45_;
      r_187__44_ <= r_n_187__44_;
      r_187__43_ <= r_n_187__43_;
      r_187__42_ <= r_n_187__42_;
      r_187__41_ <= r_n_187__41_;
      r_187__40_ <= r_n_187__40_;
      r_187__39_ <= r_n_187__39_;
      r_187__38_ <= r_n_187__38_;
      r_187__37_ <= r_n_187__37_;
      r_187__36_ <= r_n_187__36_;
      r_187__35_ <= r_n_187__35_;
      r_187__34_ <= r_n_187__34_;
      r_187__33_ <= r_n_187__33_;
      r_187__32_ <= r_n_187__32_;
      r_187__31_ <= r_n_187__31_;
      r_187__30_ <= r_n_187__30_;
      r_187__29_ <= r_n_187__29_;
      r_187__28_ <= r_n_187__28_;
      r_187__27_ <= r_n_187__27_;
      r_187__26_ <= r_n_187__26_;
      r_187__25_ <= r_n_187__25_;
      r_187__24_ <= r_n_187__24_;
      r_187__23_ <= r_n_187__23_;
      r_187__22_ <= r_n_187__22_;
      r_187__21_ <= r_n_187__21_;
      r_187__20_ <= r_n_187__20_;
      r_187__19_ <= r_n_187__19_;
      r_187__18_ <= r_n_187__18_;
      r_187__17_ <= r_n_187__17_;
      r_187__16_ <= r_n_187__16_;
      r_187__15_ <= r_n_187__15_;
      r_187__14_ <= r_n_187__14_;
      r_187__13_ <= r_n_187__13_;
      r_187__12_ <= r_n_187__12_;
      r_187__11_ <= r_n_187__11_;
      r_187__10_ <= r_n_187__10_;
      r_187__9_ <= r_n_187__9_;
      r_187__8_ <= r_n_187__8_;
      r_187__7_ <= r_n_187__7_;
      r_187__6_ <= r_n_187__6_;
      r_187__5_ <= r_n_187__5_;
      r_187__4_ <= r_n_187__4_;
      r_187__3_ <= r_n_187__3_;
      r_187__2_ <= r_n_187__2_;
      r_187__1_ <= r_n_187__1_;
      r_187__0_ <= r_n_187__0_;
    end 
    if(N3772) begin
      r_188__63_ <= r_n_188__63_;
      r_188__62_ <= r_n_188__62_;
      r_188__61_ <= r_n_188__61_;
      r_188__60_ <= r_n_188__60_;
      r_188__59_ <= r_n_188__59_;
      r_188__58_ <= r_n_188__58_;
      r_188__57_ <= r_n_188__57_;
      r_188__56_ <= r_n_188__56_;
      r_188__55_ <= r_n_188__55_;
      r_188__54_ <= r_n_188__54_;
      r_188__53_ <= r_n_188__53_;
      r_188__52_ <= r_n_188__52_;
      r_188__51_ <= r_n_188__51_;
      r_188__50_ <= r_n_188__50_;
      r_188__49_ <= r_n_188__49_;
      r_188__48_ <= r_n_188__48_;
      r_188__47_ <= r_n_188__47_;
      r_188__46_ <= r_n_188__46_;
      r_188__45_ <= r_n_188__45_;
      r_188__44_ <= r_n_188__44_;
      r_188__43_ <= r_n_188__43_;
      r_188__42_ <= r_n_188__42_;
      r_188__41_ <= r_n_188__41_;
      r_188__40_ <= r_n_188__40_;
      r_188__39_ <= r_n_188__39_;
      r_188__38_ <= r_n_188__38_;
      r_188__37_ <= r_n_188__37_;
      r_188__36_ <= r_n_188__36_;
      r_188__35_ <= r_n_188__35_;
      r_188__34_ <= r_n_188__34_;
      r_188__33_ <= r_n_188__33_;
      r_188__32_ <= r_n_188__32_;
      r_188__31_ <= r_n_188__31_;
      r_188__30_ <= r_n_188__30_;
      r_188__29_ <= r_n_188__29_;
      r_188__28_ <= r_n_188__28_;
      r_188__27_ <= r_n_188__27_;
      r_188__26_ <= r_n_188__26_;
      r_188__25_ <= r_n_188__25_;
      r_188__24_ <= r_n_188__24_;
      r_188__23_ <= r_n_188__23_;
      r_188__22_ <= r_n_188__22_;
      r_188__21_ <= r_n_188__21_;
      r_188__20_ <= r_n_188__20_;
      r_188__19_ <= r_n_188__19_;
      r_188__18_ <= r_n_188__18_;
      r_188__17_ <= r_n_188__17_;
      r_188__16_ <= r_n_188__16_;
      r_188__15_ <= r_n_188__15_;
      r_188__14_ <= r_n_188__14_;
      r_188__13_ <= r_n_188__13_;
      r_188__12_ <= r_n_188__12_;
      r_188__11_ <= r_n_188__11_;
      r_188__10_ <= r_n_188__10_;
      r_188__9_ <= r_n_188__9_;
      r_188__8_ <= r_n_188__8_;
      r_188__7_ <= r_n_188__7_;
      r_188__6_ <= r_n_188__6_;
      r_188__5_ <= r_n_188__5_;
      r_188__4_ <= r_n_188__4_;
      r_188__3_ <= r_n_188__3_;
      r_188__2_ <= r_n_188__2_;
      r_188__1_ <= r_n_188__1_;
      r_188__0_ <= r_n_188__0_;
    end 
    if(N3773) begin
      r_189__63_ <= r_n_189__63_;
      r_189__62_ <= r_n_189__62_;
      r_189__61_ <= r_n_189__61_;
      r_189__60_ <= r_n_189__60_;
      r_189__59_ <= r_n_189__59_;
      r_189__58_ <= r_n_189__58_;
      r_189__57_ <= r_n_189__57_;
      r_189__56_ <= r_n_189__56_;
      r_189__55_ <= r_n_189__55_;
      r_189__54_ <= r_n_189__54_;
      r_189__53_ <= r_n_189__53_;
      r_189__52_ <= r_n_189__52_;
      r_189__51_ <= r_n_189__51_;
      r_189__50_ <= r_n_189__50_;
      r_189__49_ <= r_n_189__49_;
      r_189__48_ <= r_n_189__48_;
      r_189__47_ <= r_n_189__47_;
      r_189__46_ <= r_n_189__46_;
      r_189__45_ <= r_n_189__45_;
      r_189__44_ <= r_n_189__44_;
      r_189__43_ <= r_n_189__43_;
      r_189__42_ <= r_n_189__42_;
      r_189__41_ <= r_n_189__41_;
      r_189__40_ <= r_n_189__40_;
      r_189__39_ <= r_n_189__39_;
      r_189__38_ <= r_n_189__38_;
      r_189__37_ <= r_n_189__37_;
      r_189__36_ <= r_n_189__36_;
      r_189__35_ <= r_n_189__35_;
      r_189__34_ <= r_n_189__34_;
      r_189__33_ <= r_n_189__33_;
      r_189__32_ <= r_n_189__32_;
      r_189__31_ <= r_n_189__31_;
      r_189__30_ <= r_n_189__30_;
      r_189__29_ <= r_n_189__29_;
      r_189__28_ <= r_n_189__28_;
      r_189__27_ <= r_n_189__27_;
      r_189__26_ <= r_n_189__26_;
      r_189__25_ <= r_n_189__25_;
      r_189__24_ <= r_n_189__24_;
      r_189__23_ <= r_n_189__23_;
      r_189__22_ <= r_n_189__22_;
      r_189__21_ <= r_n_189__21_;
      r_189__20_ <= r_n_189__20_;
      r_189__19_ <= r_n_189__19_;
      r_189__18_ <= r_n_189__18_;
      r_189__17_ <= r_n_189__17_;
      r_189__16_ <= r_n_189__16_;
      r_189__15_ <= r_n_189__15_;
      r_189__14_ <= r_n_189__14_;
      r_189__13_ <= r_n_189__13_;
      r_189__12_ <= r_n_189__12_;
      r_189__11_ <= r_n_189__11_;
      r_189__10_ <= r_n_189__10_;
      r_189__9_ <= r_n_189__9_;
      r_189__8_ <= r_n_189__8_;
      r_189__7_ <= r_n_189__7_;
      r_189__6_ <= r_n_189__6_;
      r_189__5_ <= r_n_189__5_;
      r_189__4_ <= r_n_189__4_;
      r_189__3_ <= r_n_189__3_;
      r_189__2_ <= r_n_189__2_;
      r_189__1_ <= r_n_189__1_;
      r_189__0_ <= r_n_189__0_;
    end 
    if(N3774) begin
      r_190__63_ <= r_n_190__63_;
      r_190__62_ <= r_n_190__62_;
      r_190__61_ <= r_n_190__61_;
      r_190__60_ <= r_n_190__60_;
      r_190__59_ <= r_n_190__59_;
      r_190__58_ <= r_n_190__58_;
      r_190__57_ <= r_n_190__57_;
      r_190__56_ <= r_n_190__56_;
      r_190__55_ <= r_n_190__55_;
      r_190__54_ <= r_n_190__54_;
      r_190__53_ <= r_n_190__53_;
      r_190__52_ <= r_n_190__52_;
      r_190__51_ <= r_n_190__51_;
      r_190__50_ <= r_n_190__50_;
      r_190__49_ <= r_n_190__49_;
      r_190__48_ <= r_n_190__48_;
      r_190__47_ <= r_n_190__47_;
      r_190__46_ <= r_n_190__46_;
      r_190__45_ <= r_n_190__45_;
      r_190__44_ <= r_n_190__44_;
      r_190__43_ <= r_n_190__43_;
      r_190__42_ <= r_n_190__42_;
      r_190__41_ <= r_n_190__41_;
      r_190__40_ <= r_n_190__40_;
      r_190__39_ <= r_n_190__39_;
      r_190__38_ <= r_n_190__38_;
      r_190__37_ <= r_n_190__37_;
      r_190__36_ <= r_n_190__36_;
      r_190__35_ <= r_n_190__35_;
      r_190__34_ <= r_n_190__34_;
      r_190__33_ <= r_n_190__33_;
      r_190__32_ <= r_n_190__32_;
      r_190__31_ <= r_n_190__31_;
      r_190__30_ <= r_n_190__30_;
      r_190__29_ <= r_n_190__29_;
      r_190__28_ <= r_n_190__28_;
      r_190__27_ <= r_n_190__27_;
      r_190__26_ <= r_n_190__26_;
      r_190__25_ <= r_n_190__25_;
      r_190__24_ <= r_n_190__24_;
      r_190__23_ <= r_n_190__23_;
      r_190__22_ <= r_n_190__22_;
      r_190__21_ <= r_n_190__21_;
      r_190__20_ <= r_n_190__20_;
      r_190__19_ <= r_n_190__19_;
      r_190__18_ <= r_n_190__18_;
      r_190__17_ <= r_n_190__17_;
      r_190__16_ <= r_n_190__16_;
      r_190__15_ <= r_n_190__15_;
      r_190__14_ <= r_n_190__14_;
      r_190__13_ <= r_n_190__13_;
      r_190__12_ <= r_n_190__12_;
      r_190__11_ <= r_n_190__11_;
      r_190__10_ <= r_n_190__10_;
      r_190__9_ <= r_n_190__9_;
      r_190__8_ <= r_n_190__8_;
      r_190__7_ <= r_n_190__7_;
      r_190__6_ <= r_n_190__6_;
      r_190__5_ <= r_n_190__5_;
      r_190__4_ <= r_n_190__4_;
      r_190__3_ <= r_n_190__3_;
      r_190__2_ <= r_n_190__2_;
      r_190__1_ <= r_n_190__1_;
      r_190__0_ <= r_n_190__0_;
    end 
    if(N3775) begin
      r_191__63_ <= r_n_191__63_;
      r_191__62_ <= r_n_191__62_;
      r_191__61_ <= r_n_191__61_;
      r_191__60_ <= r_n_191__60_;
      r_191__59_ <= r_n_191__59_;
      r_191__58_ <= r_n_191__58_;
      r_191__57_ <= r_n_191__57_;
      r_191__56_ <= r_n_191__56_;
      r_191__55_ <= r_n_191__55_;
      r_191__54_ <= r_n_191__54_;
      r_191__53_ <= r_n_191__53_;
      r_191__52_ <= r_n_191__52_;
      r_191__51_ <= r_n_191__51_;
      r_191__50_ <= r_n_191__50_;
      r_191__49_ <= r_n_191__49_;
      r_191__48_ <= r_n_191__48_;
      r_191__47_ <= r_n_191__47_;
      r_191__46_ <= r_n_191__46_;
      r_191__45_ <= r_n_191__45_;
      r_191__44_ <= r_n_191__44_;
      r_191__43_ <= r_n_191__43_;
      r_191__42_ <= r_n_191__42_;
      r_191__41_ <= r_n_191__41_;
      r_191__40_ <= r_n_191__40_;
      r_191__39_ <= r_n_191__39_;
      r_191__38_ <= r_n_191__38_;
      r_191__37_ <= r_n_191__37_;
      r_191__36_ <= r_n_191__36_;
      r_191__35_ <= r_n_191__35_;
      r_191__34_ <= r_n_191__34_;
      r_191__33_ <= r_n_191__33_;
      r_191__32_ <= r_n_191__32_;
      r_191__31_ <= r_n_191__31_;
      r_191__30_ <= r_n_191__30_;
      r_191__29_ <= r_n_191__29_;
      r_191__28_ <= r_n_191__28_;
      r_191__27_ <= r_n_191__27_;
      r_191__26_ <= r_n_191__26_;
      r_191__25_ <= r_n_191__25_;
      r_191__24_ <= r_n_191__24_;
      r_191__23_ <= r_n_191__23_;
      r_191__22_ <= r_n_191__22_;
      r_191__21_ <= r_n_191__21_;
      r_191__20_ <= r_n_191__20_;
      r_191__19_ <= r_n_191__19_;
      r_191__18_ <= r_n_191__18_;
      r_191__17_ <= r_n_191__17_;
      r_191__16_ <= r_n_191__16_;
      r_191__15_ <= r_n_191__15_;
      r_191__14_ <= r_n_191__14_;
      r_191__13_ <= r_n_191__13_;
      r_191__12_ <= r_n_191__12_;
      r_191__11_ <= r_n_191__11_;
      r_191__10_ <= r_n_191__10_;
      r_191__9_ <= r_n_191__9_;
      r_191__8_ <= r_n_191__8_;
      r_191__7_ <= r_n_191__7_;
      r_191__6_ <= r_n_191__6_;
      r_191__5_ <= r_n_191__5_;
      r_191__4_ <= r_n_191__4_;
      r_191__3_ <= r_n_191__3_;
      r_191__2_ <= r_n_191__2_;
      r_191__1_ <= r_n_191__1_;
      r_191__0_ <= r_n_191__0_;
    end 
    if(N3776) begin
      r_192__63_ <= r_n_192__63_;
      r_192__62_ <= r_n_192__62_;
      r_192__61_ <= r_n_192__61_;
      r_192__60_ <= r_n_192__60_;
      r_192__59_ <= r_n_192__59_;
      r_192__58_ <= r_n_192__58_;
      r_192__57_ <= r_n_192__57_;
      r_192__56_ <= r_n_192__56_;
      r_192__55_ <= r_n_192__55_;
      r_192__54_ <= r_n_192__54_;
      r_192__53_ <= r_n_192__53_;
      r_192__52_ <= r_n_192__52_;
      r_192__51_ <= r_n_192__51_;
      r_192__50_ <= r_n_192__50_;
      r_192__49_ <= r_n_192__49_;
      r_192__48_ <= r_n_192__48_;
      r_192__47_ <= r_n_192__47_;
      r_192__46_ <= r_n_192__46_;
      r_192__45_ <= r_n_192__45_;
      r_192__44_ <= r_n_192__44_;
      r_192__43_ <= r_n_192__43_;
      r_192__42_ <= r_n_192__42_;
      r_192__41_ <= r_n_192__41_;
      r_192__40_ <= r_n_192__40_;
      r_192__39_ <= r_n_192__39_;
      r_192__38_ <= r_n_192__38_;
      r_192__37_ <= r_n_192__37_;
      r_192__36_ <= r_n_192__36_;
      r_192__35_ <= r_n_192__35_;
      r_192__34_ <= r_n_192__34_;
      r_192__33_ <= r_n_192__33_;
      r_192__32_ <= r_n_192__32_;
      r_192__31_ <= r_n_192__31_;
      r_192__30_ <= r_n_192__30_;
      r_192__29_ <= r_n_192__29_;
      r_192__28_ <= r_n_192__28_;
      r_192__27_ <= r_n_192__27_;
      r_192__26_ <= r_n_192__26_;
      r_192__25_ <= r_n_192__25_;
      r_192__24_ <= r_n_192__24_;
      r_192__23_ <= r_n_192__23_;
      r_192__22_ <= r_n_192__22_;
      r_192__21_ <= r_n_192__21_;
      r_192__20_ <= r_n_192__20_;
      r_192__19_ <= r_n_192__19_;
      r_192__18_ <= r_n_192__18_;
      r_192__17_ <= r_n_192__17_;
      r_192__16_ <= r_n_192__16_;
      r_192__15_ <= r_n_192__15_;
      r_192__14_ <= r_n_192__14_;
      r_192__13_ <= r_n_192__13_;
      r_192__12_ <= r_n_192__12_;
      r_192__11_ <= r_n_192__11_;
      r_192__10_ <= r_n_192__10_;
      r_192__9_ <= r_n_192__9_;
      r_192__8_ <= r_n_192__8_;
      r_192__7_ <= r_n_192__7_;
      r_192__6_ <= r_n_192__6_;
      r_192__5_ <= r_n_192__5_;
      r_192__4_ <= r_n_192__4_;
      r_192__3_ <= r_n_192__3_;
      r_192__2_ <= r_n_192__2_;
      r_192__1_ <= r_n_192__1_;
      r_192__0_ <= r_n_192__0_;
    end 
    if(N3777) begin
      r_193__63_ <= r_n_193__63_;
      r_193__62_ <= r_n_193__62_;
      r_193__61_ <= r_n_193__61_;
      r_193__60_ <= r_n_193__60_;
      r_193__59_ <= r_n_193__59_;
      r_193__58_ <= r_n_193__58_;
      r_193__57_ <= r_n_193__57_;
      r_193__56_ <= r_n_193__56_;
      r_193__55_ <= r_n_193__55_;
      r_193__54_ <= r_n_193__54_;
      r_193__53_ <= r_n_193__53_;
      r_193__52_ <= r_n_193__52_;
      r_193__51_ <= r_n_193__51_;
      r_193__50_ <= r_n_193__50_;
      r_193__49_ <= r_n_193__49_;
      r_193__48_ <= r_n_193__48_;
      r_193__47_ <= r_n_193__47_;
      r_193__46_ <= r_n_193__46_;
      r_193__45_ <= r_n_193__45_;
      r_193__44_ <= r_n_193__44_;
      r_193__43_ <= r_n_193__43_;
      r_193__42_ <= r_n_193__42_;
      r_193__41_ <= r_n_193__41_;
      r_193__40_ <= r_n_193__40_;
      r_193__39_ <= r_n_193__39_;
      r_193__38_ <= r_n_193__38_;
      r_193__37_ <= r_n_193__37_;
      r_193__36_ <= r_n_193__36_;
      r_193__35_ <= r_n_193__35_;
      r_193__34_ <= r_n_193__34_;
      r_193__33_ <= r_n_193__33_;
      r_193__32_ <= r_n_193__32_;
      r_193__31_ <= r_n_193__31_;
      r_193__30_ <= r_n_193__30_;
      r_193__29_ <= r_n_193__29_;
      r_193__28_ <= r_n_193__28_;
      r_193__27_ <= r_n_193__27_;
      r_193__26_ <= r_n_193__26_;
      r_193__25_ <= r_n_193__25_;
      r_193__24_ <= r_n_193__24_;
      r_193__23_ <= r_n_193__23_;
      r_193__22_ <= r_n_193__22_;
      r_193__21_ <= r_n_193__21_;
      r_193__20_ <= r_n_193__20_;
      r_193__19_ <= r_n_193__19_;
      r_193__18_ <= r_n_193__18_;
      r_193__17_ <= r_n_193__17_;
      r_193__16_ <= r_n_193__16_;
      r_193__15_ <= r_n_193__15_;
      r_193__14_ <= r_n_193__14_;
      r_193__13_ <= r_n_193__13_;
      r_193__12_ <= r_n_193__12_;
      r_193__11_ <= r_n_193__11_;
      r_193__10_ <= r_n_193__10_;
      r_193__9_ <= r_n_193__9_;
      r_193__8_ <= r_n_193__8_;
      r_193__7_ <= r_n_193__7_;
      r_193__6_ <= r_n_193__6_;
      r_193__5_ <= r_n_193__5_;
      r_193__4_ <= r_n_193__4_;
      r_193__3_ <= r_n_193__3_;
      r_193__2_ <= r_n_193__2_;
      r_193__1_ <= r_n_193__1_;
      r_193__0_ <= r_n_193__0_;
    end 
    if(N3778) begin
      r_194__63_ <= r_n_194__63_;
      r_194__62_ <= r_n_194__62_;
      r_194__61_ <= r_n_194__61_;
      r_194__60_ <= r_n_194__60_;
      r_194__59_ <= r_n_194__59_;
      r_194__58_ <= r_n_194__58_;
      r_194__57_ <= r_n_194__57_;
      r_194__56_ <= r_n_194__56_;
      r_194__55_ <= r_n_194__55_;
      r_194__54_ <= r_n_194__54_;
      r_194__53_ <= r_n_194__53_;
      r_194__52_ <= r_n_194__52_;
      r_194__51_ <= r_n_194__51_;
      r_194__50_ <= r_n_194__50_;
      r_194__49_ <= r_n_194__49_;
      r_194__48_ <= r_n_194__48_;
      r_194__47_ <= r_n_194__47_;
      r_194__46_ <= r_n_194__46_;
      r_194__45_ <= r_n_194__45_;
      r_194__44_ <= r_n_194__44_;
      r_194__43_ <= r_n_194__43_;
      r_194__42_ <= r_n_194__42_;
      r_194__41_ <= r_n_194__41_;
      r_194__40_ <= r_n_194__40_;
      r_194__39_ <= r_n_194__39_;
      r_194__38_ <= r_n_194__38_;
      r_194__37_ <= r_n_194__37_;
      r_194__36_ <= r_n_194__36_;
      r_194__35_ <= r_n_194__35_;
      r_194__34_ <= r_n_194__34_;
      r_194__33_ <= r_n_194__33_;
      r_194__32_ <= r_n_194__32_;
      r_194__31_ <= r_n_194__31_;
      r_194__30_ <= r_n_194__30_;
      r_194__29_ <= r_n_194__29_;
      r_194__28_ <= r_n_194__28_;
      r_194__27_ <= r_n_194__27_;
      r_194__26_ <= r_n_194__26_;
      r_194__25_ <= r_n_194__25_;
      r_194__24_ <= r_n_194__24_;
      r_194__23_ <= r_n_194__23_;
      r_194__22_ <= r_n_194__22_;
      r_194__21_ <= r_n_194__21_;
      r_194__20_ <= r_n_194__20_;
      r_194__19_ <= r_n_194__19_;
      r_194__18_ <= r_n_194__18_;
      r_194__17_ <= r_n_194__17_;
      r_194__16_ <= r_n_194__16_;
      r_194__15_ <= r_n_194__15_;
      r_194__14_ <= r_n_194__14_;
      r_194__13_ <= r_n_194__13_;
      r_194__12_ <= r_n_194__12_;
      r_194__11_ <= r_n_194__11_;
      r_194__10_ <= r_n_194__10_;
      r_194__9_ <= r_n_194__9_;
      r_194__8_ <= r_n_194__8_;
      r_194__7_ <= r_n_194__7_;
      r_194__6_ <= r_n_194__6_;
      r_194__5_ <= r_n_194__5_;
      r_194__4_ <= r_n_194__4_;
      r_194__3_ <= r_n_194__3_;
      r_194__2_ <= r_n_194__2_;
      r_194__1_ <= r_n_194__1_;
      r_194__0_ <= r_n_194__0_;
    end 
    if(N3779) begin
      r_195__63_ <= r_n_195__63_;
      r_195__62_ <= r_n_195__62_;
      r_195__61_ <= r_n_195__61_;
      r_195__60_ <= r_n_195__60_;
      r_195__59_ <= r_n_195__59_;
      r_195__58_ <= r_n_195__58_;
      r_195__57_ <= r_n_195__57_;
      r_195__56_ <= r_n_195__56_;
      r_195__55_ <= r_n_195__55_;
      r_195__54_ <= r_n_195__54_;
      r_195__53_ <= r_n_195__53_;
      r_195__52_ <= r_n_195__52_;
      r_195__51_ <= r_n_195__51_;
      r_195__50_ <= r_n_195__50_;
      r_195__49_ <= r_n_195__49_;
      r_195__48_ <= r_n_195__48_;
      r_195__47_ <= r_n_195__47_;
      r_195__46_ <= r_n_195__46_;
      r_195__45_ <= r_n_195__45_;
      r_195__44_ <= r_n_195__44_;
      r_195__43_ <= r_n_195__43_;
      r_195__42_ <= r_n_195__42_;
      r_195__41_ <= r_n_195__41_;
      r_195__40_ <= r_n_195__40_;
      r_195__39_ <= r_n_195__39_;
      r_195__38_ <= r_n_195__38_;
      r_195__37_ <= r_n_195__37_;
      r_195__36_ <= r_n_195__36_;
      r_195__35_ <= r_n_195__35_;
      r_195__34_ <= r_n_195__34_;
      r_195__33_ <= r_n_195__33_;
      r_195__32_ <= r_n_195__32_;
      r_195__31_ <= r_n_195__31_;
      r_195__30_ <= r_n_195__30_;
      r_195__29_ <= r_n_195__29_;
      r_195__28_ <= r_n_195__28_;
      r_195__27_ <= r_n_195__27_;
      r_195__26_ <= r_n_195__26_;
      r_195__25_ <= r_n_195__25_;
      r_195__24_ <= r_n_195__24_;
      r_195__23_ <= r_n_195__23_;
      r_195__22_ <= r_n_195__22_;
      r_195__21_ <= r_n_195__21_;
      r_195__20_ <= r_n_195__20_;
      r_195__19_ <= r_n_195__19_;
      r_195__18_ <= r_n_195__18_;
      r_195__17_ <= r_n_195__17_;
      r_195__16_ <= r_n_195__16_;
      r_195__15_ <= r_n_195__15_;
      r_195__14_ <= r_n_195__14_;
      r_195__13_ <= r_n_195__13_;
      r_195__12_ <= r_n_195__12_;
      r_195__11_ <= r_n_195__11_;
      r_195__10_ <= r_n_195__10_;
      r_195__9_ <= r_n_195__9_;
      r_195__8_ <= r_n_195__8_;
      r_195__7_ <= r_n_195__7_;
      r_195__6_ <= r_n_195__6_;
      r_195__5_ <= r_n_195__5_;
      r_195__4_ <= r_n_195__4_;
      r_195__3_ <= r_n_195__3_;
      r_195__2_ <= r_n_195__2_;
      r_195__1_ <= r_n_195__1_;
      r_195__0_ <= r_n_195__0_;
    end 
    if(N3780) begin
      r_196__63_ <= r_n_196__63_;
      r_196__62_ <= r_n_196__62_;
      r_196__61_ <= r_n_196__61_;
      r_196__60_ <= r_n_196__60_;
      r_196__59_ <= r_n_196__59_;
      r_196__58_ <= r_n_196__58_;
      r_196__57_ <= r_n_196__57_;
      r_196__56_ <= r_n_196__56_;
      r_196__55_ <= r_n_196__55_;
      r_196__54_ <= r_n_196__54_;
      r_196__53_ <= r_n_196__53_;
      r_196__52_ <= r_n_196__52_;
      r_196__51_ <= r_n_196__51_;
      r_196__50_ <= r_n_196__50_;
      r_196__49_ <= r_n_196__49_;
      r_196__48_ <= r_n_196__48_;
      r_196__47_ <= r_n_196__47_;
      r_196__46_ <= r_n_196__46_;
      r_196__45_ <= r_n_196__45_;
      r_196__44_ <= r_n_196__44_;
      r_196__43_ <= r_n_196__43_;
      r_196__42_ <= r_n_196__42_;
      r_196__41_ <= r_n_196__41_;
      r_196__40_ <= r_n_196__40_;
      r_196__39_ <= r_n_196__39_;
      r_196__38_ <= r_n_196__38_;
      r_196__37_ <= r_n_196__37_;
      r_196__36_ <= r_n_196__36_;
      r_196__35_ <= r_n_196__35_;
      r_196__34_ <= r_n_196__34_;
      r_196__33_ <= r_n_196__33_;
      r_196__32_ <= r_n_196__32_;
      r_196__31_ <= r_n_196__31_;
      r_196__30_ <= r_n_196__30_;
      r_196__29_ <= r_n_196__29_;
      r_196__28_ <= r_n_196__28_;
      r_196__27_ <= r_n_196__27_;
      r_196__26_ <= r_n_196__26_;
      r_196__25_ <= r_n_196__25_;
      r_196__24_ <= r_n_196__24_;
      r_196__23_ <= r_n_196__23_;
      r_196__22_ <= r_n_196__22_;
      r_196__21_ <= r_n_196__21_;
      r_196__20_ <= r_n_196__20_;
      r_196__19_ <= r_n_196__19_;
      r_196__18_ <= r_n_196__18_;
      r_196__17_ <= r_n_196__17_;
      r_196__16_ <= r_n_196__16_;
      r_196__15_ <= r_n_196__15_;
      r_196__14_ <= r_n_196__14_;
      r_196__13_ <= r_n_196__13_;
      r_196__12_ <= r_n_196__12_;
      r_196__11_ <= r_n_196__11_;
      r_196__10_ <= r_n_196__10_;
      r_196__9_ <= r_n_196__9_;
      r_196__8_ <= r_n_196__8_;
      r_196__7_ <= r_n_196__7_;
      r_196__6_ <= r_n_196__6_;
      r_196__5_ <= r_n_196__5_;
      r_196__4_ <= r_n_196__4_;
      r_196__3_ <= r_n_196__3_;
      r_196__2_ <= r_n_196__2_;
      r_196__1_ <= r_n_196__1_;
      r_196__0_ <= r_n_196__0_;
    end 
    if(N3781) begin
      r_197__63_ <= r_n_197__63_;
      r_197__62_ <= r_n_197__62_;
      r_197__61_ <= r_n_197__61_;
      r_197__60_ <= r_n_197__60_;
      r_197__59_ <= r_n_197__59_;
      r_197__58_ <= r_n_197__58_;
      r_197__57_ <= r_n_197__57_;
      r_197__56_ <= r_n_197__56_;
      r_197__55_ <= r_n_197__55_;
      r_197__54_ <= r_n_197__54_;
      r_197__53_ <= r_n_197__53_;
      r_197__52_ <= r_n_197__52_;
      r_197__51_ <= r_n_197__51_;
      r_197__50_ <= r_n_197__50_;
      r_197__49_ <= r_n_197__49_;
      r_197__48_ <= r_n_197__48_;
      r_197__47_ <= r_n_197__47_;
      r_197__46_ <= r_n_197__46_;
      r_197__45_ <= r_n_197__45_;
      r_197__44_ <= r_n_197__44_;
      r_197__43_ <= r_n_197__43_;
      r_197__42_ <= r_n_197__42_;
      r_197__41_ <= r_n_197__41_;
      r_197__40_ <= r_n_197__40_;
      r_197__39_ <= r_n_197__39_;
      r_197__38_ <= r_n_197__38_;
      r_197__37_ <= r_n_197__37_;
      r_197__36_ <= r_n_197__36_;
      r_197__35_ <= r_n_197__35_;
      r_197__34_ <= r_n_197__34_;
      r_197__33_ <= r_n_197__33_;
      r_197__32_ <= r_n_197__32_;
      r_197__31_ <= r_n_197__31_;
      r_197__30_ <= r_n_197__30_;
      r_197__29_ <= r_n_197__29_;
      r_197__28_ <= r_n_197__28_;
      r_197__27_ <= r_n_197__27_;
      r_197__26_ <= r_n_197__26_;
      r_197__25_ <= r_n_197__25_;
      r_197__24_ <= r_n_197__24_;
      r_197__23_ <= r_n_197__23_;
      r_197__22_ <= r_n_197__22_;
      r_197__21_ <= r_n_197__21_;
      r_197__20_ <= r_n_197__20_;
      r_197__19_ <= r_n_197__19_;
      r_197__18_ <= r_n_197__18_;
      r_197__17_ <= r_n_197__17_;
      r_197__16_ <= r_n_197__16_;
      r_197__15_ <= r_n_197__15_;
      r_197__14_ <= r_n_197__14_;
      r_197__13_ <= r_n_197__13_;
      r_197__12_ <= r_n_197__12_;
      r_197__11_ <= r_n_197__11_;
      r_197__10_ <= r_n_197__10_;
      r_197__9_ <= r_n_197__9_;
      r_197__8_ <= r_n_197__8_;
      r_197__7_ <= r_n_197__7_;
      r_197__6_ <= r_n_197__6_;
      r_197__5_ <= r_n_197__5_;
      r_197__4_ <= r_n_197__4_;
      r_197__3_ <= r_n_197__3_;
      r_197__2_ <= r_n_197__2_;
      r_197__1_ <= r_n_197__1_;
      r_197__0_ <= r_n_197__0_;
    end 
    if(N3782) begin
      r_198__63_ <= r_n_198__63_;
      r_198__62_ <= r_n_198__62_;
      r_198__61_ <= r_n_198__61_;
      r_198__60_ <= r_n_198__60_;
      r_198__59_ <= r_n_198__59_;
      r_198__58_ <= r_n_198__58_;
      r_198__57_ <= r_n_198__57_;
      r_198__56_ <= r_n_198__56_;
      r_198__55_ <= r_n_198__55_;
      r_198__54_ <= r_n_198__54_;
      r_198__53_ <= r_n_198__53_;
      r_198__52_ <= r_n_198__52_;
      r_198__51_ <= r_n_198__51_;
      r_198__50_ <= r_n_198__50_;
      r_198__49_ <= r_n_198__49_;
      r_198__48_ <= r_n_198__48_;
      r_198__47_ <= r_n_198__47_;
      r_198__46_ <= r_n_198__46_;
      r_198__45_ <= r_n_198__45_;
      r_198__44_ <= r_n_198__44_;
      r_198__43_ <= r_n_198__43_;
      r_198__42_ <= r_n_198__42_;
      r_198__41_ <= r_n_198__41_;
      r_198__40_ <= r_n_198__40_;
      r_198__39_ <= r_n_198__39_;
      r_198__38_ <= r_n_198__38_;
      r_198__37_ <= r_n_198__37_;
      r_198__36_ <= r_n_198__36_;
      r_198__35_ <= r_n_198__35_;
      r_198__34_ <= r_n_198__34_;
      r_198__33_ <= r_n_198__33_;
      r_198__32_ <= r_n_198__32_;
      r_198__31_ <= r_n_198__31_;
      r_198__30_ <= r_n_198__30_;
      r_198__29_ <= r_n_198__29_;
      r_198__28_ <= r_n_198__28_;
      r_198__27_ <= r_n_198__27_;
      r_198__26_ <= r_n_198__26_;
      r_198__25_ <= r_n_198__25_;
      r_198__24_ <= r_n_198__24_;
      r_198__23_ <= r_n_198__23_;
      r_198__22_ <= r_n_198__22_;
      r_198__21_ <= r_n_198__21_;
      r_198__20_ <= r_n_198__20_;
      r_198__19_ <= r_n_198__19_;
      r_198__18_ <= r_n_198__18_;
      r_198__17_ <= r_n_198__17_;
      r_198__16_ <= r_n_198__16_;
      r_198__15_ <= r_n_198__15_;
      r_198__14_ <= r_n_198__14_;
      r_198__13_ <= r_n_198__13_;
      r_198__12_ <= r_n_198__12_;
      r_198__11_ <= r_n_198__11_;
      r_198__10_ <= r_n_198__10_;
      r_198__9_ <= r_n_198__9_;
      r_198__8_ <= r_n_198__8_;
      r_198__7_ <= r_n_198__7_;
      r_198__6_ <= r_n_198__6_;
      r_198__5_ <= r_n_198__5_;
      r_198__4_ <= r_n_198__4_;
      r_198__3_ <= r_n_198__3_;
      r_198__2_ <= r_n_198__2_;
      r_198__1_ <= r_n_198__1_;
      r_198__0_ <= r_n_198__0_;
    end 
    if(N3783) begin
      r_199__63_ <= r_n_199__63_;
      r_199__62_ <= r_n_199__62_;
      r_199__61_ <= r_n_199__61_;
      r_199__60_ <= r_n_199__60_;
      r_199__59_ <= r_n_199__59_;
      r_199__58_ <= r_n_199__58_;
      r_199__57_ <= r_n_199__57_;
      r_199__56_ <= r_n_199__56_;
      r_199__55_ <= r_n_199__55_;
      r_199__54_ <= r_n_199__54_;
      r_199__53_ <= r_n_199__53_;
      r_199__52_ <= r_n_199__52_;
      r_199__51_ <= r_n_199__51_;
      r_199__50_ <= r_n_199__50_;
      r_199__49_ <= r_n_199__49_;
      r_199__48_ <= r_n_199__48_;
      r_199__47_ <= r_n_199__47_;
      r_199__46_ <= r_n_199__46_;
      r_199__45_ <= r_n_199__45_;
      r_199__44_ <= r_n_199__44_;
      r_199__43_ <= r_n_199__43_;
      r_199__42_ <= r_n_199__42_;
      r_199__41_ <= r_n_199__41_;
      r_199__40_ <= r_n_199__40_;
      r_199__39_ <= r_n_199__39_;
      r_199__38_ <= r_n_199__38_;
      r_199__37_ <= r_n_199__37_;
      r_199__36_ <= r_n_199__36_;
      r_199__35_ <= r_n_199__35_;
      r_199__34_ <= r_n_199__34_;
      r_199__33_ <= r_n_199__33_;
      r_199__32_ <= r_n_199__32_;
      r_199__31_ <= r_n_199__31_;
      r_199__30_ <= r_n_199__30_;
      r_199__29_ <= r_n_199__29_;
      r_199__28_ <= r_n_199__28_;
      r_199__27_ <= r_n_199__27_;
      r_199__26_ <= r_n_199__26_;
      r_199__25_ <= r_n_199__25_;
      r_199__24_ <= r_n_199__24_;
      r_199__23_ <= r_n_199__23_;
      r_199__22_ <= r_n_199__22_;
      r_199__21_ <= r_n_199__21_;
      r_199__20_ <= r_n_199__20_;
      r_199__19_ <= r_n_199__19_;
      r_199__18_ <= r_n_199__18_;
      r_199__17_ <= r_n_199__17_;
      r_199__16_ <= r_n_199__16_;
      r_199__15_ <= r_n_199__15_;
      r_199__14_ <= r_n_199__14_;
      r_199__13_ <= r_n_199__13_;
      r_199__12_ <= r_n_199__12_;
      r_199__11_ <= r_n_199__11_;
      r_199__10_ <= r_n_199__10_;
      r_199__9_ <= r_n_199__9_;
      r_199__8_ <= r_n_199__8_;
      r_199__7_ <= r_n_199__7_;
      r_199__6_ <= r_n_199__6_;
      r_199__5_ <= r_n_199__5_;
      r_199__4_ <= r_n_199__4_;
      r_199__3_ <= r_n_199__3_;
      r_199__2_ <= r_n_199__2_;
      r_199__1_ <= r_n_199__1_;
      r_199__0_ <= r_n_199__0_;
    end 
    if(N3784) begin
      r_200__63_ <= r_n_200__63_;
      r_200__62_ <= r_n_200__62_;
      r_200__61_ <= r_n_200__61_;
      r_200__60_ <= r_n_200__60_;
      r_200__59_ <= r_n_200__59_;
      r_200__58_ <= r_n_200__58_;
      r_200__57_ <= r_n_200__57_;
      r_200__56_ <= r_n_200__56_;
      r_200__55_ <= r_n_200__55_;
      r_200__54_ <= r_n_200__54_;
      r_200__53_ <= r_n_200__53_;
      r_200__52_ <= r_n_200__52_;
      r_200__51_ <= r_n_200__51_;
      r_200__50_ <= r_n_200__50_;
      r_200__49_ <= r_n_200__49_;
      r_200__48_ <= r_n_200__48_;
      r_200__47_ <= r_n_200__47_;
      r_200__46_ <= r_n_200__46_;
      r_200__45_ <= r_n_200__45_;
      r_200__44_ <= r_n_200__44_;
      r_200__43_ <= r_n_200__43_;
      r_200__42_ <= r_n_200__42_;
      r_200__41_ <= r_n_200__41_;
      r_200__40_ <= r_n_200__40_;
      r_200__39_ <= r_n_200__39_;
      r_200__38_ <= r_n_200__38_;
      r_200__37_ <= r_n_200__37_;
      r_200__36_ <= r_n_200__36_;
      r_200__35_ <= r_n_200__35_;
      r_200__34_ <= r_n_200__34_;
      r_200__33_ <= r_n_200__33_;
      r_200__32_ <= r_n_200__32_;
      r_200__31_ <= r_n_200__31_;
      r_200__30_ <= r_n_200__30_;
      r_200__29_ <= r_n_200__29_;
      r_200__28_ <= r_n_200__28_;
      r_200__27_ <= r_n_200__27_;
      r_200__26_ <= r_n_200__26_;
      r_200__25_ <= r_n_200__25_;
      r_200__24_ <= r_n_200__24_;
      r_200__23_ <= r_n_200__23_;
      r_200__22_ <= r_n_200__22_;
      r_200__21_ <= r_n_200__21_;
      r_200__20_ <= r_n_200__20_;
      r_200__19_ <= r_n_200__19_;
      r_200__18_ <= r_n_200__18_;
      r_200__17_ <= r_n_200__17_;
      r_200__16_ <= r_n_200__16_;
      r_200__15_ <= r_n_200__15_;
      r_200__14_ <= r_n_200__14_;
      r_200__13_ <= r_n_200__13_;
      r_200__12_ <= r_n_200__12_;
      r_200__11_ <= r_n_200__11_;
      r_200__10_ <= r_n_200__10_;
      r_200__9_ <= r_n_200__9_;
      r_200__8_ <= r_n_200__8_;
      r_200__7_ <= r_n_200__7_;
      r_200__6_ <= r_n_200__6_;
      r_200__5_ <= r_n_200__5_;
      r_200__4_ <= r_n_200__4_;
      r_200__3_ <= r_n_200__3_;
      r_200__2_ <= r_n_200__2_;
      r_200__1_ <= r_n_200__1_;
      r_200__0_ <= r_n_200__0_;
    end 
    if(N3785) begin
      r_201__63_ <= r_n_201__63_;
      r_201__62_ <= r_n_201__62_;
      r_201__61_ <= r_n_201__61_;
      r_201__60_ <= r_n_201__60_;
      r_201__59_ <= r_n_201__59_;
      r_201__58_ <= r_n_201__58_;
      r_201__57_ <= r_n_201__57_;
      r_201__56_ <= r_n_201__56_;
      r_201__55_ <= r_n_201__55_;
      r_201__54_ <= r_n_201__54_;
      r_201__53_ <= r_n_201__53_;
      r_201__52_ <= r_n_201__52_;
      r_201__51_ <= r_n_201__51_;
      r_201__50_ <= r_n_201__50_;
      r_201__49_ <= r_n_201__49_;
      r_201__48_ <= r_n_201__48_;
      r_201__47_ <= r_n_201__47_;
      r_201__46_ <= r_n_201__46_;
      r_201__45_ <= r_n_201__45_;
      r_201__44_ <= r_n_201__44_;
      r_201__43_ <= r_n_201__43_;
      r_201__42_ <= r_n_201__42_;
      r_201__41_ <= r_n_201__41_;
      r_201__40_ <= r_n_201__40_;
      r_201__39_ <= r_n_201__39_;
      r_201__38_ <= r_n_201__38_;
      r_201__37_ <= r_n_201__37_;
      r_201__36_ <= r_n_201__36_;
      r_201__35_ <= r_n_201__35_;
      r_201__34_ <= r_n_201__34_;
      r_201__33_ <= r_n_201__33_;
      r_201__32_ <= r_n_201__32_;
      r_201__31_ <= r_n_201__31_;
      r_201__30_ <= r_n_201__30_;
      r_201__29_ <= r_n_201__29_;
      r_201__28_ <= r_n_201__28_;
      r_201__27_ <= r_n_201__27_;
      r_201__26_ <= r_n_201__26_;
      r_201__25_ <= r_n_201__25_;
      r_201__24_ <= r_n_201__24_;
      r_201__23_ <= r_n_201__23_;
      r_201__22_ <= r_n_201__22_;
      r_201__21_ <= r_n_201__21_;
      r_201__20_ <= r_n_201__20_;
      r_201__19_ <= r_n_201__19_;
      r_201__18_ <= r_n_201__18_;
      r_201__17_ <= r_n_201__17_;
      r_201__16_ <= r_n_201__16_;
      r_201__15_ <= r_n_201__15_;
      r_201__14_ <= r_n_201__14_;
      r_201__13_ <= r_n_201__13_;
      r_201__12_ <= r_n_201__12_;
      r_201__11_ <= r_n_201__11_;
      r_201__10_ <= r_n_201__10_;
      r_201__9_ <= r_n_201__9_;
      r_201__8_ <= r_n_201__8_;
      r_201__7_ <= r_n_201__7_;
      r_201__6_ <= r_n_201__6_;
      r_201__5_ <= r_n_201__5_;
      r_201__4_ <= r_n_201__4_;
      r_201__3_ <= r_n_201__3_;
      r_201__2_ <= r_n_201__2_;
      r_201__1_ <= r_n_201__1_;
      r_201__0_ <= r_n_201__0_;
    end 
    if(N3786) begin
      r_202__63_ <= r_n_202__63_;
      r_202__62_ <= r_n_202__62_;
      r_202__61_ <= r_n_202__61_;
      r_202__60_ <= r_n_202__60_;
      r_202__59_ <= r_n_202__59_;
      r_202__58_ <= r_n_202__58_;
      r_202__57_ <= r_n_202__57_;
      r_202__56_ <= r_n_202__56_;
      r_202__55_ <= r_n_202__55_;
      r_202__54_ <= r_n_202__54_;
      r_202__53_ <= r_n_202__53_;
      r_202__52_ <= r_n_202__52_;
      r_202__51_ <= r_n_202__51_;
      r_202__50_ <= r_n_202__50_;
      r_202__49_ <= r_n_202__49_;
      r_202__48_ <= r_n_202__48_;
      r_202__47_ <= r_n_202__47_;
      r_202__46_ <= r_n_202__46_;
      r_202__45_ <= r_n_202__45_;
      r_202__44_ <= r_n_202__44_;
      r_202__43_ <= r_n_202__43_;
      r_202__42_ <= r_n_202__42_;
      r_202__41_ <= r_n_202__41_;
      r_202__40_ <= r_n_202__40_;
      r_202__39_ <= r_n_202__39_;
      r_202__38_ <= r_n_202__38_;
      r_202__37_ <= r_n_202__37_;
      r_202__36_ <= r_n_202__36_;
      r_202__35_ <= r_n_202__35_;
      r_202__34_ <= r_n_202__34_;
      r_202__33_ <= r_n_202__33_;
      r_202__32_ <= r_n_202__32_;
      r_202__31_ <= r_n_202__31_;
      r_202__30_ <= r_n_202__30_;
      r_202__29_ <= r_n_202__29_;
      r_202__28_ <= r_n_202__28_;
      r_202__27_ <= r_n_202__27_;
      r_202__26_ <= r_n_202__26_;
      r_202__25_ <= r_n_202__25_;
      r_202__24_ <= r_n_202__24_;
      r_202__23_ <= r_n_202__23_;
      r_202__22_ <= r_n_202__22_;
      r_202__21_ <= r_n_202__21_;
      r_202__20_ <= r_n_202__20_;
      r_202__19_ <= r_n_202__19_;
      r_202__18_ <= r_n_202__18_;
      r_202__17_ <= r_n_202__17_;
      r_202__16_ <= r_n_202__16_;
      r_202__15_ <= r_n_202__15_;
      r_202__14_ <= r_n_202__14_;
      r_202__13_ <= r_n_202__13_;
      r_202__12_ <= r_n_202__12_;
      r_202__11_ <= r_n_202__11_;
      r_202__10_ <= r_n_202__10_;
      r_202__9_ <= r_n_202__9_;
      r_202__8_ <= r_n_202__8_;
      r_202__7_ <= r_n_202__7_;
      r_202__6_ <= r_n_202__6_;
      r_202__5_ <= r_n_202__5_;
      r_202__4_ <= r_n_202__4_;
      r_202__3_ <= r_n_202__3_;
      r_202__2_ <= r_n_202__2_;
      r_202__1_ <= r_n_202__1_;
      r_202__0_ <= r_n_202__0_;
    end 
    if(N3787) begin
      r_203__63_ <= r_n_203__63_;
      r_203__62_ <= r_n_203__62_;
      r_203__61_ <= r_n_203__61_;
      r_203__60_ <= r_n_203__60_;
      r_203__59_ <= r_n_203__59_;
      r_203__58_ <= r_n_203__58_;
      r_203__57_ <= r_n_203__57_;
      r_203__56_ <= r_n_203__56_;
      r_203__55_ <= r_n_203__55_;
      r_203__54_ <= r_n_203__54_;
      r_203__53_ <= r_n_203__53_;
      r_203__52_ <= r_n_203__52_;
      r_203__51_ <= r_n_203__51_;
      r_203__50_ <= r_n_203__50_;
      r_203__49_ <= r_n_203__49_;
      r_203__48_ <= r_n_203__48_;
      r_203__47_ <= r_n_203__47_;
      r_203__46_ <= r_n_203__46_;
      r_203__45_ <= r_n_203__45_;
      r_203__44_ <= r_n_203__44_;
      r_203__43_ <= r_n_203__43_;
      r_203__42_ <= r_n_203__42_;
      r_203__41_ <= r_n_203__41_;
      r_203__40_ <= r_n_203__40_;
      r_203__39_ <= r_n_203__39_;
      r_203__38_ <= r_n_203__38_;
      r_203__37_ <= r_n_203__37_;
      r_203__36_ <= r_n_203__36_;
      r_203__35_ <= r_n_203__35_;
      r_203__34_ <= r_n_203__34_;
      r_203__33_ <= r_n_203__33_;
      r_203__32_ <= r_n_203__32_;
      r_203__31_ <= r_n_203__31_;
      r_203__30_ <= r_n_203__30_;
      r_203__29_ <= r_n_203__29_;
      r_203__28_ <= r_n_203__28_;
      r_203__27_ <= r_n_203__27_;
      r_203__26_ <= r_n_203__26_;
      r_203__25_ <= r_n_203__25_;
      r_203__24_ <= r_n_203__24_;
      r_203__23_ <= r_n_203__23_;
      r_203__22_ <= r_n_203__22_;
      r_203__21_ <= r_n_203__21_;
      r_203__20_ <= r_n_203__20_;
      r_203__19_ <= r_n_203__19_;
      r_203__18_ <= r_n_203__18_;
      r_203__17_ <= r_n_203__17_;
      r_203__16_ <= r_n_203__16_;
      r_203__15_ <= r_n_203__15_;
      r_203__14_ <= r_n_203__14_;
      r_203__13_ <= r_n_203__13_;
      r_203__12_ <= r_n_203__12_;
      r_203__11_ <= r_n_203__11_;
      r_203__10_ <= r_n_203__10_;
      r_203__9_ <= r_n_203__9_;
      r_203__8_ <= r_n_203__8_;
      r_203__7_ <= r_n_203__7_;
      r_203__6_ <= r_n_203__6_;
      r_203__5_ <= r_n_203__5_;
      r_203__4_ <= r_n_203__4_;
      r_203__3_ <= r_n_203__3_;
      r_203__2_ <= r_n_203__2_;
      r_203__1_ <= r_n_203__1_;
      r_203__0_ <= r_n_203__0_;
    end 
    if(N3788) begin
      r_204__63_ <= r_n_204__63_;
      r_204__62_ <= r_n_204__62_;
      r_204__61_ <= r_n_204__61_;
      r_204__60_ <= r_n_204__60_;
      r_204__59_ <= r_n_204__59_;
      r_204__58_ <= r_n_204__58_;
      r_204__57_ <= r_n_204__57_;
      r_204__56_ <= r_n_204__56_;
      r_204__55_ <= r_n_204__55_;
      r_204__54_ <= r_n_204__54_;
      r_204__53_ <= r_n_204__53_;
      r_204__52_ <= r_n_204__52_;
      r_204__51_ <= r_n_204__51_;
      r_204__50_ <= r_n_204__50_;
      r_204__49_ <= r_n_204__49_;
      r_204__48_ <= r_n_204__48_;
      r_204__47_ <= r_n_204__47_;
      r_204__46_ <= r_n_204__46_;
      r_204__45_ <= r_n_204__45_;
      r_204__44_ <= r_n_204__44_;
      r_204__43_ <= r_n_204__43_;
      r_204__42_ <= r_n_204__42_;
      r_204__41_ <= r_n_204__41_;
      r_204__40_ <= r_n_204__40_;
      r_204__39_ <= r_n_204__39_;
      r_204__38_ <= r_n_204__38_;
      r_204__37_ <= r_n_204__37_;
      r_204__36_ <= r_n_204__36_;
      r_204__35_ <= r_n_204__35_;
      r_204__34_ <= r_n_204__34_;
      r_204__33_ <= r_n_204__33_;
      r_204__32_ <= r_n_204__32_;
      r_204__31_ <= r_n_204__31_;
      r_204__30_ <= r_n_204__30_;
      r_204__29_ <= r_n_204__29_;
      r_204__28_ <= r_n_204__28_;
      r_204__27_ <= r_n_204__27_;
      r_204__26_ <= r_n_204__26_;
      r_204__25_ <= r_n_204__25_;
      r_204__24_ <= r_n_204__24_;
      r_204__23_ <= r_n_204__23_;
      r_204__22_ <= r_n_204__22_;
      r_204__21_ <= r_n_204__21_;
      r_204__20_ <= r_n_204__20_;
      r_204__19_ <= r_n_204__19_;
      r_204__18_ <= r_n_204__18_;
      r_204__17_ <= r_n_204__17_;
      r_204__16_ <= r_n_204__16_;
      r_204__15_ <= r_n_204__15_;
      r_204__14_ <= r_n_204__14_;
      r_204__13_ <= r_n_204__13_;
      r_204__12_ <= r_n_204__12_;
      r_204__11_ <= r_n_204__11_;
      r_204__10_ <= r_n_204__10_;
      r_204__9_ <= r_n_204__9_;
      r_204__8_ <= r_n_204__8_;
      r_204__7_ <= r_n_204__7_;
      r_204__6_ <= r_n_204__6_;
      r_204__5_ <= r_n_204__5_;
      r_204__4_ <= r_n_204__4_;
      r_204__3_ <= r_n_204__3_;
      r_204__2_ <= r_n_204__2_;
      r_204__1_ <= r_n_204__1_;
      r_204__0_ <= r_n_204__0_;
    end 
    if(N3789) begin
      r_205__63_ <= r_n_205__63_;
      r_205__62_ <= r_n_205__62_;
      r_205__61_ <= r_n_205__61_;
      r_205__60_ <= r_n_205__60_;
      r_205__59_ <= r_n_205__59_;
      r_205__58_ <= r_n_205__58_;
      r_205__57_ <= r_n_205__57_;
      r_205__56_ <= r_n_205__56_;
      r_205__55_ <= r_n_205__55_;
      r_205__54_ <= r_n_205__54_;
      r_205__53_ <= r_n_205__53_;
      r_205__52_ <= r_n_205__52_;
      r_205__51_ <= r_n_205__51_;
      r_205__50_ <= r_n_205__50_;
      r_205__49_ <= r_n_205__49_;
      r_205__48_ <= r_n_205__48_;
      r_205__47_ <= r_n_205__47_;
      r_205__46_ <= r_n_205__46_;
      r_205__45_ <= r_n_205__45_;
      r_205__44_ <= r_n_205__44_;
      r_205__43_ <= r_n_205__43_;
      r_205__42_ <= r_n_205__42_;
      r_205__41_ <= r_n_205__41_;
      r_205__40_ <= r_n_205__40_;
      r_205__39_ <= r_n_205__39_;
      r_205__38_ <= r_n_205__38_;
      r_205__37_ <= r_n_205__37_;
      r_205__36_ <= r_n_205__36_;
      r_205__35_ <= r_n_205__35_;
      r_205__34_ <= r_n_205__34_;
      r_205__33_ <= r_n_205__33_;
      r_205__32_ <= r_n_205__32_;
      r_205__31_ <= r_n_205__31_;
      r_205__30_ <= r_n_205__30_;
      r_205__29_ <= r_n_205__29_;
      r_205__28_ <= r_n_205__28_;
      r_205__27_ <= r_n_205__27_;
      r_205__26_ <= r_n_205__26_;
      r_205__25_ <= r_n_205__25_;
      r_205__24_ <= r_n_205__24_;
      r_205__23_ <= r_n_205__23_;
      r_205__22_ <= r_n_205__22_;
      r_205__21_ <= r_n_205__21_;
      r_205__20_ <= r_n_205__20_;
      r_205__19_ <= r_n_205__19_;
      r_205__18_ <= r_n_205__18_;
      r_205__17_ <= r_n_205__17_;
      r_205__16_ <= r_n_205__16_;
      r_205__15_ <= r_n_205__15_;
      r_205__14_ <= r_n_205__14_;
      r_205__13_ <= r_n_205__13_;
      r_205__12_ <= r_n_205__12_;
      r_205__11_ <= r_n_205__11_;
      r_205__10_ <= r_n_205__10_;
      r_205__9_ <= r_n_205__9_;
      r_205__8_ <= r_n_205__8_;
      r_205__7_ <= r_n_205__7_;
      r_205__6_ <= r_n_205__6_;
      r_205__5_ <= r_n_205__5_;
      r_205__4_ <= r_n_205__4_;
      r_205__3_ <= r_n_205__3_;
      r_205__2_ <= r_n_205__2_;
      r_205__1_ <= r_n_205__1_;
      r_205__0_ <= r_n_205__0_;
    end 
    if(N3790) begin
      r_206__63_ <= r_n_206__63_;
      r_206__62_ <= r_n_206__62_;
      r_206__61_ <= r_n_206__61_;
      r_206__60_ <= r_n_206__60_;
      r_206__59_ <= r_n_206__59_;
      r_206__58_ <= r_n_206__58_;
      r_206__57_ <= r_n_206__57_;
      r_206__56_ <= r_n_206__56_;
      r_206__55_ <= r_n_206__55_;
      r_206__54_ <= r_n_206__54_;
      r_206__53_ <= r_n_206__53_;
      r_206__52_ <= r_n_206__52_;
      r_206__51_ <= r_n_206__51_;
      r_206__50_ <= r_n_206__50_;
      r_206__49_ <= r_n_206__49_;
      r_206__48_ <= r_n_206__48_;
      r_206__47_ <= r_n_206__47_;
      r_206__46_ <= r_n_206__46_;
      r_206__45_ <= r_n_206__45_;
      r_206__44_ <= r_n_206__44_;
      r_206__43_ <= r_n_206__43_;
      r_206__42_ <= r_n_206__42_;
      r_206__41_ <= r_n_206__41_;
      r_206__40_ <= r_n_206__40_;
      r_206__39_ <= r_n_206__39_;
      r_206__38_ <= r_n_206__38_;
      r_206__37_ <= r_n_206__37_;
      r_206__36_ <= r_n_206__36_;
      r_206__35_ <= r_n_206__35_;
      r_206__34_ <= r_n_206__34_;
      r_206__33_ <= r_n_206__33_;
      r_206__32_ <= r_n_206__32_;
      r_206__31_ <= r_n_206__31_;
      r_206__30_ <= r_n_206__30_;
      r_206__29_ <= r_n_206__29_;
      r_206__28_ <= r_n_206__28_;
      r_206__27_ <= r_n_206__27_;
      r_206__26_ <= r_n_206__26_;
      r_206__25_ <= r_n_206__25_;
      r_206__24_ <= r_n_206__24_;
      r_206__23_ <= r_n_206__23_;
      r_206__22_ <= r_n_206__22_;
      r_206__21_ <= r_n_206__21_;
      r_206__20_ <= r_n_206__20_;
      r_206__19_ <= r_n_206__19_;
      r_206__18_ <= r_n_206__18_;
      r_206__17_ <= r_n_206__17_;
      r_206__16_ <= r_n_206__16_;
      r_206__15_ <= r_n_206__15_;
      r_206__14_ <= r_n_206__14_;
      r_206__13_ <= r_n_206__13_;
      r_206__12_ <= r_n_206__12_;
      r_206__11_ <= r_n_206__11_;
      r_206__10_ <= r_n_206__10_;
      r_206__9_ <= r_n_206__9_;
      r_206__8_ <= r_n_206__8_;
      r_206__7_ <= r_n_206__7_;
      r_206__6_ <= r_n_206__6_;
      r_206__5_ <= r_n_206__5_;
      r_206__4_ <= r_n_206__4_;
      r_206__3_ <= r_n_206__3_;
      r_206__2_ <= r_n_206__2_;
      r_206__1_ <= r_n_206__1_;
      r_206__0_ <= r_n_206__0_;
    end 
    if(N3791) begin
      r_207__63_ <= r_n_207__63_;
      r_207__62_ <= r_n_207__62_;
      r_207__61_ <= r_n_207__61_;
      r_207__60_ <= r_n_207__60_;
      r_207__59_ <= r_n_207__59_;
      r_207__58_ <= r_n_207__58_;
      r_207__57_ <= r_n_207__57_;
      r_207__56_ <= r_n_207__56_;
      r_207__55_ <= r_n_207__55_;
      r_207__54_ <= r_n_207__54_;
      r_207__53_ <= r_n_207__53_;
      r_207__52_ <= r_n_207__52_;
      r_207__51_ <= r_n_207__51_;
      r_207__50_ <= r_n_207__50_;
      r_207__49_ <= r_n_207__49_;
      r_207__48_ <= r_n_207__48_;
      r_207__47_ <= r_n_207__47_;
      r_207__46_ <= r_n_207__46_;
      r_207__45_ <= r_n_207__45_;
      r_207__44_ <= r_n_207__44_;
      r_207__43_ <= r_n_207__43_;
      r_207__42_ <= r_n_207__42_;
      r_207__41_ <= r_n_207__41_;
      r_207__40_ <= r_n_207__40_;
      r_207__39_ <= r_n_207__39_;
      r_207__38_ <= r_n_207__38_;
      r_207__37_ <= r_n_207__37_;
      r_207__36_ <= r_n_207__36_;
      r_207__35_ <= r_n_207__35_;
      r_207__34_ <= r_n_207__34_;
      r_207__33_ <= r_n_207__33_;
      r_207__32_ <= r_n_207__32_;
      r_207__31_ <= r_n_207__31_;
      r_207__30_ <= r_n_207__30_;
      r_207__29_ <= r_n_207__29_;
      r_207__28_ <= r_n_207__28_;
      r_207__27_ <= r_n_207__27_;
      r_207__26_ <= r_n_207__26_;
      r_207__25_ <= r_n_207__25_;
      r_207__24_ <= r_n_207__24_;
      r_207__23_ <= r_n_207__23_;
      r_207__22_ <= r_n_207__22_;
      r_207__21_ <= r_n_207__21_;
      r_207__20_ <= r_n_207__20_;
      r_207__19_ <= r_n_207__19_;
      r_207__18_ <= r_n_207__18_;
      r_207__17_ <= r_n_207__17_;
      r_207__16_ <= r_n_207__16_;
      r_207__15_ <= r_n_207__15_;
      r_207__14_ <= r_n_207__14_;
      r_207__13_ <= r_n_207__13_;
      r_207__12_ <= r_n_207__12_;
      r_207__11_ <= r_n_207__11_;
      r_207__10_ <= r_n_207__10_;
      r_207__9_ <= r_n_207__9_;
      r_207__8_ <= r_n_207__8_;
      r_207__7_ <= r_n_207__7_;
      r_207__6_ <= r_n_207__6_;
      r_207__5_ <= r_n_207__5_;
      r_207__4_ <= r_n_207__4_;
      r_207__3_ <= r_n_207__3_;
      r_207__2_ <= r_n_207__2_;
      r_207__1_ <= r_n_207__1_;
      r_207__0_ <= r_n_207__0_;
    end 
    if(N3792) begin
      r_208__63_ <= r_n_208__63_;
      r_208__62_ <= r_n_208__62_;
      r_208__61_ <= r_n_208__61_;
      r_208__60_ <= r_n_208__60_;
      r_208__59_ <= r_n_208__59_;
      r_208__58_ <= r_n_208__58_;
      r_208__57_ <= r_n_208__57_;
      r_208__56_ <= r_n_208__56_;
      r_208__55_ <= r_n_208__55_;
      r_208__54_ <= r_n_208__54_;
      r_208__53_ <= r_n_208__53_;
      r_208__52_ <= r_n_208__52_;
      r_208__51_ <= r_n_208__51_;
      r_208__50_ <= r_n_208__50_;
      r_208__49_ <= r_n_208__49_;
      r_208__48_ <= r_n_208__48_;
      r_208__47_ <= r_n_208__47_;
      r_208__46_ <= r_n_208__46_;
      r_208__45_ <= r_n_208__45_;
      r_208__44_ <= r_n_208__44_;
      r_208__43_ <= r_n_208__43_;
      r_208__42_ <= r_n_208__42_;
      r_208__41_ <= r_n_208__41_;
      r_208__40_ <= r_n_208__40_;
      r_208__39_ <= r_n_208__39_;
      r_208__38_ <= r_n_208__38_;
      r_208__37_ <= r_n_208__37_;
      r_208__36_ <= r_n_208__36_;
      r_208__35_ <= r_n_208__35_;
      r_208__34_ <= r_n_208__34_;
      r_208__33_ <= r_n_208__33_;
      r_208__32_ <= r_n_208__32_;
      r_208__31_ <= r_n_208__31_;
      r_208__30_ <= r_n_208__30_;
      r_208__29_ <= r_n_208__29_;
      r_208__28_ <= r_n_208__28_;
      r_208__27_ <= r_n_208__27_;
      r_208__26_ <= r_n_208__26_;
      r_208__25_ <= r_n_208__25_;
      r_208__24_ <= r_n_208__24_;
      r_208__23_ <= r_n_208__23_;
      r_208__22_ <= r_n_208__22_;
      r_208__21_ <= r_n_208__21_;
      r_208__20_ <= r_n_208__20_;
      r_208__19_ <= r_n_208__19_;
      r_208__18_ <= r_n_208__18_;
      r_208__17_ <= r_n_208__17_;
      r_208__16_ <= r_n_208__16_;
      r_208__15_ <= r_n_208__15_;
      r_208__14_ <= r_n_208__14_;
      r_208__13_ <= r_n_208__13_;
      r_208__12_ <= r_n_208__12_;
      r_208__11_ <= r_n_208__11_;
      r_208__10_ <= r_n_208__10_;
      r_208__9_ <= r_n_208__9_;
      r_208__8_ <= r_n_208__8_;
      r_208__7_ <= r_n_208__7_;
      r_208__6_ <= r_n_208__6_;
      r_208__5_ <= r_n_208__5_;
      r_208__4_ <= r_n_208__4_;
      r_208__3_ <= r_n_208__3_;
      r_208__2_ <= r_n_208__2_;
      r_208__1_ <= r_n_208__1_;
      r_208__0_ <= r_n_208__0_;
    end 
    if(N3793) begin
      r_209__63_ <= r_n_209__63_;
      r_209__62_ <= r_n_209__62_;
      r_209__61_ <= r_n_209__61_;
      r_209__60_ <= r_n_209__60_;
      r_209__59_ <= r_n_209__59_;
      r_209__58_ <= r_n_209__58_;
      r_209__57_ <= r_n_209__57_;
      r_209__56_ <= r_n_209__56_;
      r_209__55_ <= r_n_209__55_;
      r_209__54_ <= r_n_209__54_;
      r_209__53_ <= r_n_209__53_;
      r_209__52_ <= r_n_209__52_;
      r_209__51_ <= r_n_209__51_;
      r_209__50_ <= r_n_209__50_;
      r_209__49_ <= r_n_209__49_;
      r_209__48_ <= r_n_209__48_;
      r_209__47_ <= r_n_209__47_;
      r_209__46_ <= r_n_209__46_;
      r_209__45_ <= r_n_209__45_;
      r_209__44_ <= r_n_209__44_;
      r_209__43_ <= r_n_209__43_;
      r_209__42_ <= r_n_209__42_;
      r_209__41_ <= r_n_209__41_;
      r_209__40_ <= r_n_209__40_;
      r_209__39_ <= r_n_209__39_;
      r_209__38_ <= r_n_209__38_;
      r_209__37_ <= r_n_209__37_;
      r_209__36_ <= r_n_209__36_;
      r_209__35_ <= r_n_209__35_;
      r_209__34_ <= r_n_209__34_;
      r_209__33_ <= r_n_209__33_;
      r_209__32_ <= r_n_209__32_;
      r_209__31_ <= r_n_209__31_;
      r_209__30_ <= r_n_209__30_;
      r_209__29_ <= r_n_209__29_;
      r_209__28_ <= r_n_209__28_;
      r_209__27_ <= r_n_209__27_;
      r_209__26_ <= r_n_209__26_;
      r_209__25_ <= r_n_209__25_;
      r_209__24_ <= r_n_209__24_;
      r_209__23_ <= r_n_209__23_;
      r_209__22_ <= r_n_209__22_;
      r_209__21_ <= r_n_209__21_;
      r_209__20_ <= r_n_209__20_;
      r_209__19_ <= r_n_209__19_;
      r_209__18_ <= r_n_209__18_;
      r_209__17_ <= r_n_209__17_;
      r_209__16_ <= r_n_209__16_;
      r_209__15_ <= r_n_209__15_;
      r_209__14_ <= r_n_209__14_;
      r_209__13_ <= r_n_209__13_;
      r_209__12_ <= r_n_209__12_;
      r_209__11_ <= r_n_209__11_;
      r_209__10_ <= r_n_209__10_;
      r_209__9_ <= r_n_209__9_;
      r_209__8_ <= r_n_209__8_;
      r_209__7_ <= r_n_209__7_;
      r_209__6_ <= r_n_209__6_;
      r_209__5_ <= r_n_209__5_;
      r_209__4_ <= r_n_209__4_;
      r_209__3_ <= r_n_209__3_;
      r_209__2_ <= r_n_209__2_;
      r_209__1_ <= r_n_209__1_;
      r_209__0_ <= r_n_209__0_;
    end 
    if(N3794) begin
      r_210__63_ <= r_n_210__63_;
      r_210__62_ <= r_n_210__62_;
      r_210__61_ <= r_n_210__61_;
      r_210__60_ <= r_n_210__60_;
      r_210__59_ <= r_n_210__59_;
      r_210__58_ <= r_n_210__58_;
      r_210__57_ <= r_n_210__57_;
      r_210__56_ <= r_n_210__56_;
      r_210__55_ <= r_n_210__55_;
      r_210__54_ <= r_n_210__54_;
      r_210__53_ <= r_n_210__53_;
      r_210__52_ <= r_n_210__52_;
      r_210__51_ <= r_n_210__51_;
      r_210__50_ <= r_n_210__50_;
      r_210__49_ <= r_n_210__49_;
      r_210__48_ <= r_n_210__48_;
      r_210__47_ <= r_n_210__47_;
      r_210__46_ <= r_n_210__46_;
      r_210__45_ <= r_n_210__45_;
      r_210__44_ <= r_n_210__44_;
      r_210__43_ <= r_n_210__43_;
      r_210__42_ <= r_n_210__42_;
      r_210__41_ <= r_n_210__41_;
      r_210__40_ <= r_n_210__40_;
      r_210__39_ <= r_n_210__39_;
      r_210__38_ <= r_n_210__38_;
      r_210__37_ <= r_n_210__37_;
      r_210__36_ <= r_n_210__36_;
      r_210__35_ <= r_n_210__35_;
      r_210__34_ <= r_n_210__34_;
      r_210__33_ <= r_n_210__33_;
      r_210__32_ <= r_n_210__32_;
      r_210__31_ <= r_n_210__31_;
      r_210__30_ <= r_n_210__30_;
      r_210__29_ <= r_n_210__29_;
      r_210__28_ <= r_n_210__28_;
      r_210__27_ <= r_n_210__27_;
      r_210__26_ <= r_n_210__26_;
      r_210__25_ <= r_n_210__25_;
      r_210__24_ <= r_n_210__24_;
      r_210__23_ <= r_n_210__23_;
      r_210__22_ <= r_n_210__22_;
      r_210__21_ <= r_n_210__21_;
      r_210__20_ <= r_n_210__20_;
      r_210__19_ <= r_n_210__19_;
      r_210__18_ <= r_n_210__18_;
      r_210__17_ <= r_n_210__17_;
      r_210__16_ <= r_n_210__16_;
      r_210__15_ <= r_n_210__15_;
      r_210__14_ <= r_n_210__14_;
      r_210__13_ <= r_n_210__13_;
      r_210__12_ <= r_n_210__12_;
      r_210__11_ <= r_n_210__11_;
      r_210__10_ <= r_n_210__10_;
      r_210__9_ <= r_n_210__9_;
      r_210__8_ <= r_n_210__8_;
      r_210__7_ <= r_n_210__7_;
      r_210__6_ <= r_n_210__6_;
      r_210__5_ <= r_n_210__5_;
      r_210__4_ <= r_n_210__4_;
      r_210__3_ <= r_n_210__3_;
      r_210__2_ <= r_n_210__2_;
      r_210__1_ <= r_n_210__1_;
      r_210__0_ <= r_n_210__0_;
    end 
    if(N3795) begin
      r_211__63_ <= r_n_211__63_;
      r_211__62_ <= r_n_211__62_;
      r_211__61_ <= r_n_211__61_;
      r_211__60_ <= r_n_211__60_;
      r_211__59_ <= r_n_211__59_;
      r_211__58_ <= r_n_211__58_;
      r_211__57_ <= r_n_211__57_;
      r_211__56_ <= r_n_211__56_;
      r_211__55_ <= r_n_211__55_;
      r_211__54_ <= r_n_211__54_;
      r_211__53_ <= r_n_211__53_;
      r_211__52_ <= r_n_211__52_;
      r_211__51_ <= r_n_211__51_;
      r_211__50_ <= r_n_211__50_;
      r_211__49_ <= r_n_211__49_;
      r_211__48_ <= r_n_211__48_;
      r_211__47_ <= r_n_211__47_;
      r_211__46_ <= r_n_211__46_;
      r_211__45_ <= r_n_211__45_;
      r_211__44_ <= r_n_211__44_;
      r_211__43_ <= r_n_211__43_;
      r_211__42_ <= r_n_211__42_;
      r_211__41_ <= r_n_211__41_;
      r_211__40_ <= r_n_211__40_;
      r_211__39_ <= r_n_211__39_;
      r_211__38_ <= r_n_211__38_;
      r_211__37_ <= r_n_211__37_;
      r_211__36_ <= r_n_211__36_;
      r_211__35_ <= r_n_211__35_;
      r_211__34_ <= r_n_211__34_;
      r_211__33_ <= r_n_211__33_;
      r_211__32_ <= r_n_211__32_;
      r_211__31_ <= r_n_211__31_;
      r_211__30_ <= r_n_211__30_;
      r_211__29_ <= r_n_211__29_;
      r_211__28_ <= r_n_211__28_;
      r_211__27_ <= r_n_211__27_;
      r_211__26_ <= r_n_211__26_;
      r_211__25_ <= r_n_211__25_;
      r_211__24_ <= r_n_211__24_;
      r_211__23_ <= r_n_211__23_;
      r_211__22_ <= r_n_211__22_;
      r_211__21_ <= r_n_211__21_;
      r_211__20_ <= r_n_211__20_;
      r_211__19_ <= r_n_211__19_;
      r_211__18_ <= r_n_211__18_;
      r_211__17_ <= r_n_211__17_;
      r_211__16_ <= r_n_211__16_;
      r_211__15_ <= r_n_211__15_;
      r_211__14_ <= r_n_211__14_;
      r_211__13_ <= r_n_211__13_;
      r_211__12_ <= r_n_211__12_;
      r_211__11_ <= r_n_211__11_;
      r_211__10_ <= r_n_211__10_;
      r_211__9_ <= r_n_211__9_;
      r_211__8_ <= r_n_211__8_;
      r_211__7_ <= r_n_211__7_;
      r_211__6_ <= r_n_211__6_;
      r_211__5_ <= r_n_211__5_;
      r_211__4_ <= r_n_211__4_;
      r_211__3_ <= r_n_211__3_;
      r_211__2_ <= r_n_211__2_;
      r_211__1_ <= r_n_211__1_;
      r_211__0_ <= r_n_211__0_;
    end 
    if(N3796) begin
      r_212__63_ <= r_n_212__63_;
      r_212__62_ <= r_n_212__62_;
      r_212__61_ <= r_n_212__61_;
      r_212__60_ <= r_n_212__60_;
      r_212__59_ <= r_n_212__59_;
      r_212__58_ <= r_n_212__58_;
      r_212__57_ <= r_n_212__57_;
      r_212__56_ <= r_n_212__56_;
      r_212__55_ <= r_n_212__55_;
      r_212__54_ <= r_n_212__54_;
      r_212__53_ <= r_n_212__53_;
      r_212__52_ <= r_n_212__52_;
      r_212__51_ <= r_n_212__51_;
      r_212__50_ <= r_n_212__50_;
      r_212__49_ <= r_n_212__49_;
      r_212__48_ <= r_n_212__48_;
      r_212__47_ <= r_n_212__47_;
      r_212__46_ <= r_n_212__46_;
      r_212__45_ <= r_n_212__45_;
      r_212__44_ <= r_n_212__44_;
      r_212__43_ <= r_n_212__43_;
      r_212__42_ <= r_n_212__42_;
      r_212__41_ <= r_n_212__41_;
      r_212__40_ <= r_n_212__40_;
      r_212__39_ <= r_n_212__39_;
      r_212__38_ <= r_n_212__38_;
      r_212__37_ <= r_n_212__37_;
      r_212__36_ <= r_n_212__36_;
      r_212__35_ <= r_n_212__35_;
      r_212__34_ <= r_n_212__34_;
      r_212__33_ <= r_n_212__33_;
      r_212__32_ <= r_n_212__32_;
      r_212__31_ <= r_n_212__31_;
      r_212__30_ <= r_n_212__30_;
      r_212__29_ <= r_n_212__29_;
      r_212__28_ <= r_n_212__28_;
      r_212__27_ <= r_n_212__27_;
      r_212__26_ <= r_n_212__26_;
      r_212__25_ <= r_n_212__25_;
      r_212__24_ <= r_n_212__24_;
      r_212__23_ <= r_n_212__23_;
      r_212__22_ <= r_n_212__22_;
      r_212__21_ <= r_n_212__21_;
      r_212__20_ <= r_n_212__20_;
      r_212__19_ <= r_n_212__19_;
      r_212__18_ <= r_n_212__18_;
      r_212__17_ <= r_n_212__17_;
      r_212__16_ <= r_n_212__16_;
      r_212__15_ <= r_n_212__15_;
      r_212__14_ <= r_n_212__14_;
      r_212__13_ <= r_n_212__13_;
      r_212__12_ <= r_n_212__12_;
      r_212__11_ <= r_n_212__11_;
      r_212__10_ <= r_n_212__10_;
      r_212__9_ <= r_n_212__9_;
      r_212__8_ <= r_n_212__8_;
      r_212__7_ <= r_n_212__7_;
      r_212__6_ <= r_n_212__6_;
      r_212__5_ <= r_n_212__5_;
      r_212__4_ <= r_n_212__4_;
      r_212__3_ <= r_n_212__3_;
      r_212__2_ <= r_n_212__2_;
      r_212__1_ <= r_n_212__1_;
      r_212__0_ <= r_n_212__0_;
    end 
    if(N3797) begin
      r_213__63_ <= r_n_213__63_;
      r_213__62_ <= r_n_213__62_;
      r_213__61_ <= r_n_213__61_;
      r_213__60_ <= r_n_213__60_;
      r_213__59_ <= r_n_213__59_;
      r_213__58_ <= r_n_213__58_;
      r_213__57_ <= r_n_213__57_;
      r_213__56_ <= r_n_213__56_;
      r_213__55_ <= r_n_213__55_;
      r_213__54_ <= r_n_213__54_;
      r_213__53_ <= r_n_213__53_;
      r_213__52_ <= r_n_213__52_;
      r_213__51_ <= r_n_213__51_;
      r_213__50_ <= r_n_213__50_;
      r_213__49_ <= r_n_213__49_;
      r_213__48_ <= r_n_213__48_;
      r_213__47_ <= r_n_213__47_;
      r_213__46_ <= r_n_213__46_;
      r_213__45_ <= r_n_213__45_;
      r_213__44_ <= r_n_213__44_;
      r_213__43_ <= r_n_213__43_;
      r_213__42_ <= r_n_213__42_;
      r_213__41_ <= r_n_213__41_;
      r_213__40_ <= r_n_213__40_;
      r_213__39_ <= r_n_213__39_;
      r_213__38_ <= r_n_213__38_;
      r_213__37_ <= r_n_213__37_;
      r_213__36_ <= r_n_213__36_;
      r_213__35_ <= r_n_213__35_;
      r_213__34_ <= r_n_213__34_;
      r_213__33_ <= r_n_213__33_;
      r_213__32_ <= r_n_213__32_;
      r_213__31_ <= r_n_213__31_;
      r_213__30_ <= r_n_213__30_;
      r_213__29_ <= r_n_213__29_;
      r_213__28_ <= r_n_213__28_;
      r_213__27_ <= r_n_213__27_;
      r_213__26_ <= r_n_213__26_;
      r_213__25_ <= r_n_213__25_;
      r_213__24_ <= r_n_213__24_;
      r_213__23_ <= r_n_213__23_;
      r_213__22_ <= r_n_213__22_;
      r_213__21_ <= r_n_213__21_;
      r_213__20_ <= r_n_213__20_;
      r_213__19_ <= r_n_213__19_;
      r_213__18_ <= r_n_213__18_;
      r_213__17_ <= r_n_213__17_;
      r_213__16_ <= r_n_213__16_;
      r_213__15_ <= r_n_213__15_;
      r_213__14_ <= r_n_213__14_;
      r_213__13_ <= r_n_213__13_;
      r_213__12_ <= r_n_213__12_;
      r_213__11_ <= r_n_213__11_;
      r_213__10_ <= r_n_213__10_;
      r_213__9_ <= r_n_213__9_;
      r_213__8_ <= r_n_213__8_;
      r_213__7_ <= r_n_213__7_;
      r_213__6_ <= r_n_213__6_;
      r_213__5_ <= r_n_213__5_;
      r_213__4_ <= r_n_213__4_;
      r_213__3_ <= r_n_213__3_;
      r_213__2_ <= r_n_213__2_;
      r_213__1_ <= r_n_213__1_;
      r_213__0_ <= r_n_213__0_;
    end 
    if(N3798) begin
      r_214__63_ <= r_n_214__63_;
      r_214__62_ <= r_n_214__62_;
      r_214__61_ <= r_n_214__61_;
      r_214__60_ <= r_n_214__60_;
      r_214__59_ <= r_n_214__59_;
      r_214__58_ <= r_n_214__58_;
      r_214__57_ <= r_n_214__57_;
      r_214__56_ <= r_n_214__56_;
      r_214__55_ <= r_n_214__55_;
      r_214__54_ <= r_n_214__54_;
      r_214__53_ <= r_n_214__53_;
      r_214__52_ <= r_n_214__52_;
      r_214__51_ <= r_n_214__51_;
      r_214__50_ <= r_n_214__50_;
      r_214__49_ <= r_n_214__49_;
      r_214__48_ <= r_n_214__48_;
      r_214__47_ <= r_n_214__47_;
      r_214__46_ <= r_n_214__46_;
      r_214__45_ <= r_n_214__45_;
      r_214__44_ <= r_n_214__44_;
      r_214__43_ <= r_n_214__43_;
      r_214__42_ <= r_n_214__42_;
      r_214__41_ <= r_n_214__41_;
      r_214__40_ <= r_n_214__40_;
      r_214__39_ <= r_n_214__39_;
      r_214__38_ <= r_n_214__38_;
      r_214__37_ <= r_n_214__37_;
      r_214__36_ <= r_n_214__36_;
      r_214__35_ <= r_n_214__35_;
      r_214__34_ <= r_n_214__34_;
      r_214__33_ <= r_n_214__33_;
      r_214__32_ <= r_n_214__32_;
      r_214__31_ <= r_n_214__31_;
      r_214__30_ <= r_n_214__30_;
      r_214__29_ <= r_n_214__29_;
      r_214__28_ <= r_n_214__28_;
      r_214__27_ <= r_n_214__27_;
      r_214__26_ <= r_n_214__26_;
      r_214__25_ <= r_n_214__25_;
      r_214__24_ <= r_n_214__24_;
      r_214__23_ <= r_n_214__23_;
      r_214__22_ <= r_n_214__22_;
      r_214__21_ <= r_n_214__21_;
      r_214__20_ <= r_n_214__20_;
      r_214__19_ <= r_n_214__19_;
      r_214__18_ <= r_n_214__18_;
      r_214__17_ <= r_n_214__17_;
      r_214__16_ <= r_n_214__16_;
      r_214__15_ <= r_n_214__15_;
      r_214__14_ <= r_n_214__14_;
      r_214__13_ <= r_n_214__13_;
      r_214__12_ <= r_n_214__12_;
      r_214__11_ <= r_n_214__11_;
      r_214__10_ <= r_n_214__10_;
      r_214__9_ <= r_n_214__9_;
      r_214__8_ <= r_n_214__8_;
      r_214__7_ <= r_n_214__7_;
      r_214__6_ <= r_n_214__6_;
      r_214__5_ <= r_n_214__5_;
      r_214__4_ <= r_n_214__4_;
      r_214__3_ <= r_n_214__3_;
      r_214__2_ <= r_n_214__2_;
      r_214__1_ <= r_n_214__1_;
      r_214__0_ <= r_n_214__0_;
    end 
    if(N3799) begin
      r_215__63_ <= r_n_215__63_;
      r_215__62_ <= r_n_215__62_;
      r_215__61_ <= r_n_215__61_;
      r_215__60_ <= r_n_215__60_;
      r_215__59_ <= r_n_215__59_;
      r_215__58_ <= r_n_215__58_;
      r_215__57_ <= r_n_215__57_;
      r_215__56_ <= r_n_215__56_;
      r_215__55_ <= r_n_215__55_;
      r_215__54_ <= r_n_215__54_;
      r_215__53_ <= r_n_215__53_;
      r_215__52_ <= r_n_215__52_;
      r_215__51_ <= r_n_215__51_;
      r_215__50_ <= r_n_215__50_;
      r_215__49_ <= r_n_215__49_;
      r_215__48_ <= r_n_215__48_;
      r_215__47_ <= r_n_215__47_;
      r_215__46_ <= r_n_215__46_;
      r_215__45_ <= r_n_215__45_;
      r_215__44_ <= r_n_215__44_;
      r_215__43_ <= r_n_215__43_;
      r_215__42_ <= r_n_215__42_;
      r_215__41_ <= r_n_215__41_;
      r_215__40_ <= r_n_215__40_;
      r_215__39_ <= r_n_215__39_;
      r_215__38_ <= r_n_215__38_;
      r_215__37_ <= r_n_215__37_;
      r_215__36_ <= r_n_215__36_;
      r_215__35_ <= r_n_215__35_;
      r_215__34_ <= r_n_215__34_;
      r_215__33_ <= r_n_215__33_;
      r_215__32_ <= r_n_215__32_;
      r_215__31_ <= r_n_215__31_;
      r_215__30_ <= r_n_215__30_;
      r_215__29_ <= r_n_215__29_;
      r_215__28_ <= r_n_215__28_;
      r_215__27_ <= r_n_215__27_;
      r_215__26_ <= r_n_215__26_;
      r_215__25_ <= r_n_215__25_;
      r_215__24_ <= r_n_215__24_;
      r_215__23_ <= r_n_215__23_;
      r_215__22_ <= r_n_215__22_;
      r_215__21_ <= r_n_215__21_;
      r_215__20_ <= r_n_215__20_;
      r_215__19_ <= r_n_215__19_;
      r_215__18_ <= r_n_215__18_;
      r_215__17_ <= r_n_215__17_;
      r_215__16_ <= r_n_215__16_;
      r_215__15_ <= r_n_215__15_;
      r_215__14_ <= r_n_215__14_;
      r_215__13_ <= r_n_215__13_;
      r_215__12_ <= r_n_215__12_;
      r_215__11_ <= r_n_215__11_;
      r_215__10_ <= r_n_215__10_;
      r_215__9_ <= r_n_215__9_;
      r_215__8_ <= r_n_215__8_;
      r_215__7_ <= r_n_215__7_;
      r_215__6_ <= r_n_215__6_;
      r_215__5_ <= r_n_215__5_;
      r_215__4_ <= r_n_215__4_;
      r_215__3_ <= r_n_215__3_;
      r_215__2_ <= r_n_215__2_;
      r_215__1_ <= r_n_215__1_;
      r_215__0_ <= r_n_215__0_;
    end 
    if(N3800) begin
      r_216__63_ <= r_n_216__63_;
      r_216__62_ <= r_n_216__62_;
      r_216__61_ <= r_n_216__61_;
      r_216__60_ <= r_n_216__60_;
      r_216__59_ <= r_n_216__59_;
      r_216__58_ <= r_n_216__58_;
      r_216__57_ <= r_n_216__57_;
      r_216__56_ <= r_n_216__56_;
      r_216__55_ <= r_n_216__55_;
      r_216__54_ <= r_n_216__54_;
      r_216__53_ <= r_n_216__53_;
      r_216__52_ <= r_n_216__52_;
      r_216__51_ <= r_n_216__51_;
      r_216__50_ <= r_n_216__50_;
      r_216__49_ <= r_n_216__49_;
      r_216__48_ <= r_n_216__48_;
      r_216__47_ <= r_n_216__47_;
      r_216__46_ <= r_n_216__46_;
      r_216__45_ <= r_n_216__45_;
      r_216__44_ <= r_n_216__44_;
      r_216__43_ <= r_n_216__43_;
      r_216__42_ <= r_n_216__42_;
      r_216__41_ <= r_n_216__41_;
      r_216__40_ <= r_n_216__40_;
      r_216__39_ <= r_n_216__39_;
      r_216__38_ <= r_n_216__38_;
      r_216__37_ <= r_n_216__37_;
      r_216__36_ <= r_n_216__36_;
      r_216__35_ <= r_n_216__35_;
      r_216__34_ <= r_n_216__34_;
      r_216__33_ <= r_n_216__33_;
      r_216__32_ <= r_n_216__32_;
      r_216__31_ <= r_n_216__31_;
      r_216__30_ <= r_n_216__30_;
      r_216__29_ <= r_n_216__29_;
      r_216__28_ <= r_n_216__28_;
      r_216__27_ <= r_n_216__27_;
      r_216__26_ <= r_n_216__26_;
      r_216__25_ <= r_n_216__25_;
      r_216__24_ <= r_n_216__24_;
      r_216__23_ <= r_n_216__23_;
      r_216__22_ <= r_n_216__22_;
      r_216__21_ <= r_n_216__21_;
      r_216__20_ <= r_n_216__20_;
      r_216__19_ <= r_n_216__19_;
      r_216__18_ <= r_n_216__18_;
      r_216__17_ <= r_n_216__17_;
      r_216__16_ <= r_n_216__16_;
      r_216__15_ <= r_n_216__15_;
      r_216__14_ <= r_n_216__14_;
      r_216__13_ <= r_n_216__13_;
      r_216__12_ <= r_n_216__12_;
      r_216__11_ <= r_n_216__11_;
      r_216__10_ <= r_n_216__10_;
      r_216__9_ <= r_n_216__9_;
      r_216__8_ <= r_n_216__8_;
      r_216__7_ <= r_n_216__7_;
      r_216__6_ <= r_n_216__6_;
      r_216__5_ <= r_n_216__5_;
      r_216__4_ <= r_n_216__4_;
      r_216__3_ <= r_n_216__3_;
      r_216__2_ <= r_n_216__2_;
      r_216__1_ <= r_n_216__1_;
      r_216__0_ <= r_n_216__0_;
    end 
    if(N3801) begin
      r_217__63_ <= r_n_217__63_;
      r_217__62_ <= r_n_217__62_;
      r_217__61_ <= r_n_217__61_;
      r_217__60_ <= r_n_217__60_;
      r_217__59_ <= r_n_217__59_;
      r_217__58_ <= r_n_217__58_;
      r_217__57_ <= r_n_217__57_;
      r_217__56_ <= r_n_217__56_;
      r_217__55_ <= r_n_217__55_;
      r_217__54_ <= r_n_217__54_;
      r_217__53_ <= r_n_217__53_;
      r_217__52_ <= r_n_217__52_;
      r_217__51_ <= r_n_217__51_;
      r_217__50_ <= r_n_217__50_;
      r_217__49_ <= r_n_217__49_;
      r_217__48_ <= r_n_217__48_;
      r_217__47_ <= r_n_217__47_;
      r_217__46_ <= r_n_217__46_;
      r_217__45_ <= r_n_217__45_;
      r_217__44_ <= r_n_217__44_;
      r_217__43_ <= r_n_217__43_;
      r_217__42_ <= r_n_217__42_;
      r_217__41_ <= r_n_217__41_;
      r_217__40_ <= r_n_217__40_;
      r_217__39_ <= r_n_217__39_;
      r_217__38_ <= r_n_217__38_;
      r_217__37_ <= r_n_217__37_;
      r_217__36_ <= r_n_217__36_;
      r_217__35_ <= r_n_217__35_;
      r_217__34_ <= r_n_217__34_;
      r_217__33_ <= r_n_217__33_;
      r_217__32_ <= r_n_217__32_;
      r_217__31_ <= r_n_217__31_;
      r_217__30_ <= r_n_217__30_;
      r_217__29_ <= r_n_217__29_;
      r_217__28_ <= r_n_217__28_;
      r_217__27_ <= r_n_217__27_;
      r_217__26_ <= r_n_217__26_;
      r_217__25_ <= r_n_217__25_;
      r_217__24_ <= r_n_217__24_;
      r_217__23_ <= r_n_217__23_;
      r_217__22_ <= r_n_217__22_;
      r_217__21_ <= r_n_217__21_;
      r_217__20_ <= r_n_217__20_;
      r_217__19_ <= r_n_217__19_;
      r_217__18_ <= r_n_217__18_;
      r_217__17_ <= r_n_217__17_;
      r_217__16_ <= r_n_217__16_;
      r_217__15_ <= r_n_217__15_;
      r_217__14_ <= r_n_217__14_;
      r_217__13_ <= r_n_217__13_;
      r_217__12_ <= r_n_217__12_;
      r_217__11_ <= r_n_217__11_;
      r_217__10_ <= r_n_217__10_;
      r_217__9_ <= r_n_217__9_;
      r_217__8_ <= r_n_217__8_;
      r_217__7_ <= r_n_217__7_;
      r_217__6_ <= r_n_217__6_;
      r_217__5_ <= r_n_217__5_;
      r_217__4_ <= r_n_217__4_;
      r_217__3_ <= r_n_217__3_;
      r_217__2_ <= r_n_217__2_;
      r_217__1_ <= r_n_217__1_;
      r_217__0_ <= r_n_217__0_;
    end 
    if(N3802) begin
      r_218__63_ <= r_n_218__63_;
      r_218__62_ <= r_n_218__62_;
      r_218__61_ <= r_n_218__61_;
      r_218__60_ <= r_n_218__60_;
      r_218__59_ <= r_n_218__59_;
      r_218__58_ <= r_n_218__58_;
      r_218__57_ <= r_n_218__57_;
      r_218__56_ <= r_n_218__56_;
      r_218__55_ <= r_n_218__55_;
      r_218__54_ <= r_n_218__54_;
      r_218__53_ <= r_n_218__53_;
      r_218__52_ <= r_n_218__52_;
      r_218__51_ <= r_n_218__51_;
      r_218__50_ <= r_n_218__50_;
      r_218__49_ <= r_n_218__49_;
      r_218__48_ <= r_n_218__48_;
      r_218__47_ <= r_n_218__47_;
      r_218__46_ <= r_n_218__46_;
      r_218__45_ <= r_n_218__45_;
      r_218__44_ <= r_n_218__44_;
      r_218__43_ <= r_n_218__43_;
      r_218__42_ <= r_n_218__42_;
      r_218__41_ <= r_n_218__41_;
      r_218__40_ <= r_n_218__40_;
      r_218__39_ <= r_n_218__39_;
      r_218__38_ <= r_n_218__38_;
      r_218__37_ <= r_n_218__37_;
      r_218__36_ <= r_n_218__36_;
      r_218__35_ <= r_n_218__35_;
      r_218__34_ <= r_n_218__34_;
      r_218__33_ <= r_n_218__33_;
      r_218__32_ <= r_n_218__32_;
      r_218__31_ <= r_n_218__31_;
      r_218__30_ <= r_n_218__30_;
      r_218__29_ <= r_n_218__29_;
      r_218__28_ <= r_n_218__28_;
      r_218__27_ <= r_n_218__27_;
      r_218__26_ <= r_n_218__26_;
      r_218__25_ <= r_n_218__25_;
      r_218__24_ <= r_n_218__24_;
      r_218__23_ <= r_n_218__23_;
      r_218__22_ <= r_n_218__22_;
      r_218__21_ <= r_n_218__21_;
      r_218__20_ <= r_n_218__20_;
      r_218__19_ <= r_n_218__19_;
      r_218__18_ <= r_n_218__18_;
      r_218__17_ <= r_n_218__17_;
      r_218__16_ <= r_n_218__16_;
      r_218__15_ <= r_n_218__15_;
      r_218__14_ <= r_n_218__14_;
      r_218__13_ <= r_n_218__13_;
      r_218__12_ <= r_n_218__12_;
      r_218__11_ <= r_n_218__11_;
      r_218__10_ <= r_n_218__10_;
      r_218__9_ <= r_n_218__9_;
      r_218__8_ <= r_n_218__8_;
      r_218__7_ <= r_n_218__7_;
      r_218__6_ <= r_n_218__6_;
      r_218__5_ <= r_n_218__5_;
      r_218__4_ <= r_n_218__4_;
      r_218__3_ <= r_n_218__3_;
      r_218__2_ <= r_n_218__2_;
      r_218__1_ <= r_n_218__1_;
      r_218__0_ <= r_n_218__0_;
    end 
    if(N3803) begin
      r_219__63_ <= r_n_219__63_;
      r_219__62_ <= r_n_219__62_;
      r_219__61_ <= r_n_219__61_;
      r_219__60_ <= r_n_219__60_;
      r_219__59_ <= r_n_219__59_;
      r_219__58_ <= r_n_219__58_;
      r_219__57_ <= r_n_219__57_;
      r_219__56_ <= r_n_219__56_;
      r_219__55_ <= r_n_219__55_;
      r_219__54_ <= r_n_219__54_;
      r_219__53_ <= r_n_219__53_;
      r_219__52_ <= r_n_219__52_;
      r_219__51_ <= r_n_219__51_;
      r_219__50_ <= r_n_219__50_;
      r_219__49_ <= r_n_219__49_;
      r_219__48_ <= r_n_219__48_;
      r_219__47_ <= r_n_219__47_;
      r_219__46_ <= r_n_219__46_;
      r_219__45_ <= r_n_219__45_;
      r_219__44_ <= r_n_219__44_;
      r_219__43_ <= r_n_219__43_;
      r_219__42_ <= r_n_219__42_;
      r_219__41_ <= r_n_219__41_;
      r_219__40_ <= r_n_219__40_;
      r_219__39_ <= r_n_219__39_;
      r_219__38_ <= r_n_219__38_;
      r_219__37_ <= r_n_219__37_;
      r_219__36_ <= r_n_219__36_;
      r_219__35_ <= r_n_219__35_;
      r_219__34_ <= r_n_219__34_;
      r_219__33_ <= r_n_219__33_;
      r_219__32_ <= r_n_219__32_;
      r_219__31_ <= r_n_219__31_;
      r_219__30_ <= r_n_219__30_;
      r_219__29_ <= r_n_219__29_;
      r_219__28_ <= r_n_219__28_;
      r_219__27_ <= r_n_219__27_;
      r_219__26_ <= r_n_219__26_;
      r_219__25_ <= r_n_219__25_;
      r_219__24_ <= r_n_219__24_;
      r_219__23_ <= r_n_219__23_;
      r_219__22_ <= r_n_219__22_;
      r_219__21_ <= r_n_219__21_;
      r_219__20_ <= r_n_219__20_;
      r_219__19_ <= r_n_219__19_;
      r_219__18_ <= r_n_219__18_;
      r_219__17_ <= r_n_219__17_;
      r_219__16_ <= r_n_219__16_;
      r_219__15_ <= r_n_219__15_;
      r_219__14_ <= r_n_219__14_;
      r_219__13_ <= r_n_219__13_;
      r_219__12_ <= r_n_219__12_;
      r_219__11_ <= r_n_219__11_;
      r_219__10_ <= r_n_219__10_;
      r_219__9_ <= r_n_219__9_;
      r_219__8_ <= r_n_219__8_;
      r_219__7_ <= r_n_219__7_;
      r_219__6_ <= r_n_219__6_;
      r_219__5_ <= r_n_219__5_;
      r_219__4_ <= r_n_219__4_;
      r_219__3_ <= r_n_219__3_;
      r_219__2_ <= r_n_219__2_;
      r_219__1_ <= r_n_219__1_;
      r_219__0_ <= r_n_219__0_;
    end 
    if(N3804) begin
      r_220__63_ <= r_n_220__63_;
      r_220__62_ <= r_n_220__62_;
      r_220__61_ <= r_n_220__61_;
      r_220__60_ <= r_n_220__60_;
      r_220__59_ <= r_n_220__59_;
      r_220__58_ <= r_n_220__58_;
      r_220__57_ <= r_n_220__57_;
      r_220__56_ <= r_n_220__56_;
      r_220__55_ <= r_n_220__55_;
      r_220__54_ <= r_n_220__54_;
      r_220__53_ <= r_n_220__53_;
      r_220__52_ <= r_n_220__52_;
      r_220__51_ <= r_n_220__51_;
      r_220__50_ <= r_n_220__50_;
      r_220__49_ <= r_n_220__49_;
      r_220__48_ <= r_n_220__48_;
      r_220__47_ <= r_n_220__47_;
      r_220__46_ <= r_n_220__46_;
      r_220__45_ <= r_n_220__45_;
      r_220__44_ <= r_n_220__44_;
      r_220__43_ <= r_n_220__43_;
      r_220__42_ <= r_n_220__42_;
      r_220__41_ <= r_n_220__41_;
      r_220__40_ <= r_n_220__40_;
      r_220__39_ <= r_n_220__39_;
      r_220__38_ <= r_n_220__38_;
      r_220__37_ <= r_n_220__37_;
      r_220__36_ <= r_n_220__36_;
      r_220__35_ <= r_n_220__35_;
      r_220__34_ <= r_n_220__34_;
      r_220__33_ <= r_n_220__33_;
      r_220__32_ <= r_n_220__32_;
      r_220__31_ <= r_n_220__31_;
      r_220__30_ <= r_n_220__30_;
      r_220__29_ <= r_n_220__29_;
      r_220__28_ <= r_n_220__28_;
      r_220__27_ <= r_n_220__27_;
      r_220__26_ <= r_n_220__26_;
      r_220__25_ <= r_n_220__25_;
      r_220__24_ <= r_n_220__24_;
      r_220__23_ <= r_n_220__23_;
      r_220__22_ <= r_n_220__22_;
      r_220__21_ <= r_n_220__21_;
      r_220__20_ <= r_n_220__20_;
      r_220__19_ <= r_n_220__19_;
      r_220__18_ <= r_n_220__18_;
      r_220__17_ <= r_n_220__17_;
      r_220__16_ <= r_n_220__16_;
      r_220__15_ <= r_n_220__15_;
      r_220__14_ <= r_n_220__14_;
      r_220__13_ <= r_n_220__13_;
      r_220__12_ <= r_n_220__12_;
      r_220__11_ <= r_n_220__11_;
      r_220__10_ <= r_n_220__10_;
      r_220__9_ <= r_n_220__9_;
      r_220__8_ <= r_n_220__8_;
      r_220__7_ <= r_n_220__7_;
      r_220__6_ <= r_n_220__6_;
      r_220__5_ <= r_n_220__5_;
      r_220__4_ <= r_n_220__4_;
      r_220__3_ <= r_n_220__3_;
      r_220__2_ <= r_n_220__2_;
      r_220__1_ <= r_n_220__1_;
      r_220__0_ <= r_n_220__0_;
    end 
    if(N3805) begin
      r_221__63_ <= r_n_221__63_;
      r_221__62_ <= r_n_221__62_;
      r_221__61_ <= r_n_221__61_;
      r_221__60_ <= r_n_221__60_;
      r_221__59_ <= r_n_221__59_;
      r_221__58_ <= r_n_221__58_;
      r_221__57_ <= r_n_221__57_;
      r_221__56_ <= r_n_221__56_;
      r_221__55_ <= r_n_221__55_;
      r_221__54_ <= r_n_221__54_;
      r_221__53_ <= r_n_221__53_;
      r_221__52_ <= r_n_221__52_;
      r_221__51_ <= r_n_221__51_;
      r_221__50_ <= r_n_221__50_;
      r_221__49_ <= r_n_221__49_;
      r_221__48_ <= r_n_221__48_;
      r_221__47_ <= r_n_221__47_;
      r_221__46_ <= r_n_221__46_;
      r_221__45_ <= r_n_221__45_;
      r_221__44_ <= r_n_221__44_;
      r_221__43_ <= r_n_221__43_;
      r_221__42_ <= r_n_221__42_;
      r_221__41_ <= r_n_221__41_;
      r_221__40_ <= r_n_221__40_;
      r_221__39_ <= r_n_221__39_;
      r_221__38_ <= r_n_221__38_;
      r_221__37_ <= r_n_221__37_;
      r_221__36_ <= r_n_221__36_;
      r_221__35_ <= r_n_221__35_;
      r_221__34_ <= r_n_221__34_;
      r_221__33_ <= r_n_221__33_;
      r_221__32_ <= r_n_221__32_;
      r_221__31_ <= r_n_221__31_;
      r_221__30_ <= r_n_221__30_;
      r_221__29_ <= r_n_221__29_;
      r_221__28_ <= r_n_221__28_;
      r_221__27_ <= r_n_221__27_;
      r_221__26_ <= r_n_221__26_;
      r_221__25_ <= r_n_221__25_;
      r_221__24_ <= r_n_221__24_;
      r_221__23_ <= r_n_221__23_;
      r_221__22_ <= r_n_221__22_;
      r_221__21_ <= r_n_221__21_;
      r_221__20_ <= r_n_221__20_;
      r_221__19_ <= r_n_221__19_;
      r_221__18_ <= r_n_221__18_;
      r_221__17_ <= r_n_221__17_;
      r_221__16_ <= r_n_221__16_;
      r_221__15_ <= r_n_221__15_;
      r_221__14_ <= r_n_221__14_;
      r_221__13_ <= r_n_221__13_;
      r_221__12_ <= r_n_221__12_;
      r_221__11_ <= r_n_221__11_;
      r_221__10_ <= r_n_221__10_;
      r_221__9_ <= r_n_221__9_;
      r_221__8_ <= r_n_221__8_;
      r_221__7_ <= r_n_221__7_;
      r_221__6_ <= r_n_221__6_;
      r_221__5_ <= r_n_221__5_;
      r_221__4_ <= r_n_221__4_;
      r_221__3_ <= r_n_221__3_;
      r_221__2_ <= r_n_221__2_;
      r_221__1_ <= r_n_221__1_;
      r_221__0_ <= r_n_221__0_;
    end 
    if(N3806) begin
      r_222__63_ <= r_n_222__63_;
      r_222__62_ <= r_n_222__62_;
      r_222__61_ <= r_n_222__61_;
      r_222__60_ <= r_n_222__60_;
      r_222__59_ <= r_n_222__59_;
      r_222__58_ <= r_n_222__58_;
      r_222__57_ <= r_n_222__57_;
      r_222__56_ <= r_n_222__56_;
      r_222__55_ <= r_n_222__55_;
      r_222__54_ <= r_n_222__54_;
      r_222__53_ <= r_n_222__53_;
      r_222__52_ <= r_n_222__52_;
      r_222__51_ <= r_n_222__51_;
      r_222__50_ <= r_n_222__50_;
      r_222__49_ <= r_n_222__49_;
      r_222__48_ <= r_n_222__48_;
      r_222__47_ <= r_n_222__47_;
      r_222__46_ <= r_n_222__46_;
      r_222__45_ <= r_n_222__45_;
      r_222__44_ <= r_n_222__44_;
      r_222__43_ <= r_n_222__43_;
      r_222__42_ <= r_n_222__42_;
      r_222__41_ <= r_n_222__41_;
      r_222__40_ <= r_n_222__40_;
      r_222__39_ <= r_n_222__39_;
      r_222__38_ <= r_n_222__38_;
      r_222__37_ <= r_n_222__37_;
      r_222__36_ <= r_n_222__36_;
      r_222__35_ <= r_n_222__35_;
      r_222__34_ <= r_n_222__34_;
      r_222__33_ <= r_n_222__33_;
      r_222__32_ <= r_n_222__32_;
      r_222__31_ <= r_n_222__31_;
      r_222__30_ <= r_n_222__30_;
      r_222__29_ <= r_n_222__29_;
      r_222__28_ <= r_n_222__28_;
      r_222__27_ <= r_n_222__27_;
      r_222__26_ <= r_n_222__26_;
      r_222__25_ <= r_n_222__25_;
      r_222__24_ <= r_n_222__24_;
      r_222__23_ <= r_n_222__23_;
      r_222__22_ <= r_n_222__22_;
      r_222__21_ <= r_n_222__21_;
      r_222__20_ <= r_n_222__20_;
      r_222__19_ <= r_n_222__19_;
      r_222__18_ <= r_n_222__18_;
      r_222__17_ <= r_n_222__17_;
      r_222__16_ <= r_n_222__16_;
      r_222__15_ <= r_n_222__15_;
      r_222__14_ <= r_n_222__14_;
      r_222__13_ <= r_n_222__13_;
      r_222__12_ <= r_n_222__12_;
      r_222__11_ <= r_n_222__11_;
      r_222__10_ <= r_n_222__10_;
      r_222__9_ <= r_n_222__9_;
      r_222__8_ <= r_n_222__8_;
      r_222__7_ <= r_n_222__7_;
      r_222__6_ <= r_n_222__6_;
      r_222__5_ <= r_n_222__5_;
      r_222__4_ <= r_n_222__4_;
      r_222__3_ <= r_n_222__3_;
      r_222__2_ <= r_n_222__2_;
      r_222__1_ <= r_n_222__1_;
      r_222__0_ <= r_n_222__0_;
    end 
    if(N3807) begin
      r_223__63_ <= r_n_223__63_;
      r_223__62_ <= r_n_223__62_;
      r_223__61_ <= r_n_223__61_;
      r_223__60_ <= r_n_223__60_;
      r_223__59_ <= r_n_223__59_;
      r_223__58_ <= r_n_223__58_;
      r_223__57_ <= r_n_223__57_;
      r_223__56_ <= r_n_223__56_;
      r_223__55_ <= r_n_223__55_;
      r_223__54_ <= r_n_223__54_;
      r_223__53_ <= r_n_223__53_;
      r_223__52_ <= r_n_223__52_;
      r_223__51_ <= r_n_223__51_;
      r_223__50_ <= r_n_223__50_;
      r_223__49_ <= r_n_223__49_;
      r_223__48_ <= r_n_223__48_;
      r_223__47_ <= r_n_223__47_;
      r_223__46_ <= r_n_223__46_;
      r_223__45_ <= r_n_223__45_;
      r_223__44_ <= r_n_223__44_;
      r_223__43_ <= r_n_223__43_;
      r_223__42_ <= r_n_223__42_;
      r_223__41_ <= r_n_223__41_;
      r_223__40_ <= r_n_223__40_;
      r_223__39_ <= r_n_223__39_;
      r_223__38_ <= r_n_223__38_;
      r_223__37_ <= r_n_223__37_;
      r_223__36_ <= r_n_223__36_;
      r_223__35_ <= r_n_223__35_;
      r_223__34_ <= r_n_223__34_;
      r_223__33_ <= r_n_223__33_;
      r_223__32_ <= r_n_223__32_;
      r_223__31_ <= r_n_223__31_;
      r_223__30_ <= r_n_223__30_;
      r_223__29_ <= r_n_223__29_;
      r_223__28_ <= r_n_223__28_;
      r_223__27_ <= r_n_223__27_;
      r_223__26_ <= r_n_223__26_;
      r_223__25_ <= r_n_223__25_;
      r_223__24_ <= r_n_223__24_;
      r_223__23_ <= r_n_223__23_;
      r_223__22_ <= r_n_223__22_;
      r_223__21_ <= r_n_223__21_;
      r_223__20_ <= r_n_223__20_;
      r_223__19_ <= r_n_223__19_;
      r_223__18_ <= r_n_223__18_;
      r_223__17_ <= r_n_223__17_;
      r_223__16_ <= r_n_223__16_;
      r_223__15_ <= r_n_223__15_;
      r_223__14_ <= r_n_223__14_;
      r_223__13_ <= r_n_223__13_;
      r_223__12_ <= r_n_223__12_;
      r_223__11_ <= r_n_223__11_;
      r_223__10_ <= r_n_223__10_;
      r_223__9_ <= r_n_223__9_;
      r_223__8_ <= r_n_223__8_;
      r_223__7_ <= r_n_223__7_;
      r_223__6_ <= r_n_223__6_;
      r_223__5_ <= r_n_223__5_;
      r_223__4_ <= r_n_223__4_;
      r_223__3_ <= r_n_223__3_;
      r_223__2_ <= r_n_223__2_;
      r_223__1_ <= r_n_223__1_;
      r_223__0_ <= r_n_223__0_;
    end 
    if(N3808) begin
      r_224__63_ <= r_n_224__63_;
      r_224__62_ <= r_n_224__62_;
      r_224__61_ <= r_n_224__61_;
      r_224__60_ <= r_n_224__60_;
      r_224__59_ <= r_n_224__59_;
      r_224__58_ <= r_n_224__58_;
      r_224__57_ <= r_n_224__57_;
      r_224__56_ <= r_n_224__56_;
      r_224__55_ <= r_n_224__55_;
      r_224__54_ <= r_n_224__54_;
      r_224__53_ <= r_n_224__53_;
      r_224__52_ <= r_n_224__52_;
      r_224__51_ <= r_n_224__51_;
      r_224__50_ <= r_n_224__50_;
      r_224__49_ <= r_n_224__49_;
      r_224__48_ <= r_n_224__48_;
      r_224__47_ <= r_n_224__47_;
      r_224__46_ <= r_n_224__46_;
      r_224__45_ <= r_n_224__45_;
      r_224__44_ <= r_n_224__44_;
      r_224__43_ <= r_n_224__43_;
      r_224__42_ <= r_n_224__42_;
      r_224__41_ <= r_n_224__41_;
      r_224__40_ <= r_n_224__40_;
      r_224__39_ <= r_n_224__39_;
      r_224__38_ <= r_n_224__38_;
      r_224__37_ <= r_n_224__37_;
      r_224__36_ <= r_n_224__36_;
      r_224__35_ <= r_n_224__35_;
      r_224__34_ <= r_n_224__34_;
      r_224__33_ <= r_n_224__33_;
      r_224__32_ <= r_n_224__32_;
      r_224__31_ <= r_n_224__31_;
      r_224__30_ <= r_n_224__30_;
      r_224__29_ <= r_n_224__29_;
      r_224__28_ <= r_n_224__28_;
      r_224__27_ <= r_n_224__27_;
      r_224__26_ <= r_n_224__26_;
      r_224__25_ <= r_n_224__25_;
      r_224__24_ <= r_n_224__24_;
      r_224__23_ <= r_n_224__23_;
      r_224__22_ <= r_n_224__22_;
      r_224__21_ <= r_n_224__21_;
      r_224__20_ <= r_n_224__20_;
      r_224__19_ <= r_n_224__19_;
      r_224__18_ <= r_n_224__18_;
      r_224__17_ <= r_n_224__17_;
      r_224__16_ <= r_n_224__16_;
      r_224__15_ <= r_n_224__15_;
      r_224__14_ <= r_n_224__14_;
      r_224__13_ <= r_n_224__13_;
      r_224__12_ <= r_n_224__12_;
      r_224__11_ <= r_n_224__11_;
      r_224__10_ <= r_n_224__10_;
      r_224__9_ <= r_n_224__9_;
      r_224__8_ <= r_n_224__8_;
      r_224__7_ <= r_n_224__7_;
      r_224__6_ <= r_n_224__6_;
      r_224__5_ <= r_n_224__5_;
      r_224__4_ <= r_n_224__4_;
      r_224__3_ <= r_n_224__3_;
      r_224__2_ <= r_n_224__2_;
      r_224__1_ <= r_n_224__1_;
      r_224__0_ <= r_n_224__0_;
    end 
    if(N3809) begin
      r_225__63_ <= r_n_225__63_;
      r_225__62_ <= r_n_225__62_;
      r_225__61_ <= r_n_225__61_;
      r_225__60_ <= r_n_225__60_;
      r_225__59_ <= r_n_225__59_;
      r_225__58_ <= r_n_225__58_;
      r_225__57_ <= r_n_225__57_;
      r_225__56_ <= r_n_225__56_;
      r_225__55_ <= r_n_225__55_;
      r_225__54_ <= r_n_225__54_;
      r_225__53_ <= r_n_225__53_;
      r_225__52_ <= r_n_225__52_;
      r_225__51_ <= r_n_225__51_;
      r_225__50_ <= r_n_225__50_;
      r_225__49_ <= r_n_225__49_;
      r_225__48_ <= r_n_225__48_;
      r_225__47_ <= r_n_225__47_;
      r_225__46_ <= r_n_225__46_;
      r_225__45_ <= r_n_225__45_;
      r_225__44_ <= r_n_225__44_;
      r_225__43_ <= r_n_225__43_;
      r_225__42_ <= r_n_225__42_;
      r_225__41_ <= r_n_225__41_;
      r_225__40_ <= r_n_225__40_;
      r_225__39_ <= r_n_225__39_;
      r_225__38_ <= r_n_225__38_;
      r_225__37_ <= r_n_225__37_;
      r_225__36_ <= r_n_225__36_;
      r_225__35_ <= r_n_225__35_;
      r_225__34_ <= r_n_225__34_;
      r_225__33_ <= r_n_225__33_;
      r_225__32_ <= r_n_225__32_;
      r_225__31_ <= r_n_225__31_;
      r_225__30_ <= r_n_225__30_;
      r_225__29_ <= r_n_225__29_;
      r_225__28_ <= r_n_225__28_;
      r_225__27_ <= r_n_225__27_;
      r_225__26_ <= r_n_225__26_;
      r_225__25_ <= r_n_225__25_;
      r_225__24_ <= r_n_225__24_;
      r_225__23_ <= r_n_225__23_;
      r_225__22_ <= r_n_225__22_;
      r_225__21_ <= r_n_225__21_;
      r_225__20_ <= r_n_225__20_;
      r_225__19_ <= r_n_225__19_;
      r_225__18_ <= r_n_225__18_;
      r_225__17_ <= r_n_225__17_;
      r_225__16_ <= r_n_225__16_;
      r_225__15_ <= r_n_225__15_;
      r_225__14_ <= r_n_225__14_;
      r_225__13_ <= r_n_225__13_;
      r_225__12_ <= r_n_225__12_;
      r_225__11_ <= r_n_225__11_;
      r_225__10_ <= r_n_225__10_;
      r_225__9_ <= r_n_225__9_;
      r_225__8_ <= r_n_225__8_;
      r_225__7_ <= r_n_225__7_;
      r_225__6_ <= r_n_225__6_;
      r_225__5_ <= r_n_225__5_;
      r_225__4_ <= r_n_225__4_;
      r_225__3_ <= r_n_225__3_;
      r_225__2_ <= r_n_225__2_;
      r_225__1_ <= r_n_225__1_;
      r_225__0_ <= r_n_225__0_;
    end 
    if(N3810) begin
      r_226__63_ <= r_n_226__63_;
      r_226__62_ <= r_n_226__62_;
      r_226__61_ <= r_n_226__61_;
      r_226__60_ <= r_n_226__60_;
      r_226__59_ <= r_n_226__59_;
      r_226__58_ <= r_n_226__58_;
      r_226__57_ <= r_n_226__57_;
      r_226__56_ <= r_n_226__56_;
      r_226__55_ <= r_n_226__55_;
      r_226__54_ <= r_n_226__54_;
      r_226__53_ <= r_n_226__53_;
      r_226__52_ <= r_n_226__52_;
      r_226__51_ <= r_n_226__51_;
      r_226__50_ <= r_n_226__50_;
      r_226__49_ <= r_n_226__49_;
      r_226__48_ <= r_n_226__48_;
      r_226__47_ <= r_n_226__47_;
      r_226__46_ <= r_n_226__46_;
      r_226__45_ <= r_n_226__45_;
      r_226__44_ <= r_n_226__44_;
      r_226__43_ <= r_n_226__43_;
      r_226__42_ <= r_n_226__42_;
      r_226__41_ <= r_n_226__41_;
      r_226__40_ <= r_n_226__40_;
      r_226__39_ <= r_n_226__39_;
      r_226__38_ <= r_n_226__38_;
      r_226__37_ <= r_n_226__37_;
      r_226__36_ <= r_n_226__36_;
      r_226__35_ <= r_n_226__35_;
      r_226__34_ <= r_n_226__34_;
      r_226__33_ <= r_n_226__33_;
      r_226__32_ <= r_n_226__32_;
      r_226__31_ <= r_n_226__31_;
      r_226__30_ <= r_n_226__30_;
      r_226__29_ <= r_n_226__29_;
      r_226__28_ <= r_n_226__28_;
      r_226__27_ <= r_n_226__27_;
      r_226__26_ <= r_n_226__26_;
      r_226__25_ <= r_n_226__25_;
      r_226__24_ <= r_n_226__24_;
      r_226__23_ <= r_n_226__23_;
      r_226__22_ <= r_n_226__22_;
      r_226__21_ <= r_n_226__21_;
      r_226__20_ <= r_n_226__20_;
      r_226__19_ <= r_n_226__19_;
      r_226__18_ <= r_n_226__18_;
      r_226__17_ <= r_n_226__17_;
      r_226__16_ <= r_n_226__16_;
      r_226__15_ <= r_n_226__15_;
      r_226__14_ <= r_n_226__14_;
      r_226__13_ <= r_n_226__13_;
      r_226__12_ <= r_n_226__12_;
      r_226__11_ <= r_n_226__11_;
      r_226__10_ <= r_n_226__10_;
      r_226__9_ <= r_n_226__9_;
      r_226__8_ <= r_n_226__8_;
      r_226__7_ <= r_n_226__7_;
      r_226__6_ <= r_n_226__6_;
      r_226__5_ <= r_n_226__5_;
      r_226__4_ <= r_n_226__4_;
      r_226__3_ <= r_n_226__3_;
      r_226__2_ <= r_n_226__2_;
      r_226__1_ <= r_n_226__1_;
      r_226__0_ <= r_n_226__0_;
    end 
    if(N3811) begin
      r_227__63_ <= r_n_227__63_;
      r_227__62_ <= r_n_227__62_;
      r_227__61_ <= r_n_227__61_;
      r_227__60_ <= r_n_227__60_;
      r_227__59_ <= r_n_227__59_;
      r_227__58_ <= r_n_227__58_;
      r_227__57_ <= r_n_227__57_;
      r_227__56_ <= r_n_227__56_;
      r_227__55_ <= r_n_227__55_;
      r_227__54_ <= r_n_227__54_;
      r_227__53_ <= r_n_227__53_;
      r_227__52_ <= r_n_227__52_;
      r_227__51_ <= r_n_227__51_;
      r_227__50_ <= r_n_227__50_;
      r_227__49_ <= r_n_227__49_;
      r_227__48_ <= r_n_227__48_;
      r_227__47_ <= r_n_227__47_;
      r_227__46_ <= r_n_227__46_;
      r_227__45_ <= r_n_227__45_;
      r_227__44_ <= r_n_227__44_;
      r_227__43_ <= r_n_227__43_;
      r_227__42_ <= r_n_227__42_;
      r_227__41_ <= r_n_227__41_;
      r_227__40_ <= r_n_227__40_;
      r_227__39_ <= r_n_227__39_;
      r_227__38_ <= r_n_227__38_;
      r_227__37_ <= r_n_227__37_;
      r_227__36_ <= r_n_227__36_;
      r_227__35_ <= r_n_227__35_;
      r_227__34_ <= r_n_227__34_;
      r_227__33_ <= r_n_227__33_;
      r_227__32_ <= r_n_227__32_;
      r_227__31_ <= r_n_227__31_;
      r_227__30_ <= r_n_227__30_;
      r_227__29_ <= r_n_227__29_;
      r_227__28_ <= r_n_227__28_;
      r_227__27_ <= r_n_227__27_;
      r_227__26_ <= r_n_227__26_;
      r_227__25_ <= r_n_227__25_;
      r_227__24_ <= r_n_227__24_;
      r_227__23_ <= r_n_227__23_;
      r_227__22_ <= r_n_227__22_;
      r_227__21_ <= r_n_227__21_;
      r_227__20_ <= r_n_227__20_;
      r_227__19_ <= r_n_227__19_;
      r_227__18_ <= r_n_227__18_;
      r_227__17_ <= r_n_227__17_;
      r_227__16_ <= r_n_227__16_;
      r_227__15_ <= r_n_227__15_;
      r_227__14_ <= r_n_227__14_;
      r_227__13_ <= r_n_227__13_;
      r_227__12_ <= r_n_227__12_;
      r_227__11_ <= r_n_227__11_;
      r_227__10_ <= r_n_227__10_;
      r_227__9_ <= r_n_227__9_;
      r_227__8_ <= r_n_227__8_;
      r_227__7_ <= r_n_227__7_;
      r_227__6_ <= r_n_227__6_;
      r_227__5_ <= r_n_227__5_;
      r_227__4_ <= r_n_227__4_;
      r_227__3_ <= r_n_227__3_;
      r_227__2_ <= r_n_227__2_;
      r_227__1_ <= r_n_227__1_;
      r_227__0_ <= r_n_227__0_;
    end 
    if(N3812) begin
      r_228__63_ <= r_n_228__63_;
      r_228__62_ <= r_n_228__62_;
      r_228__61_ <= r_n_228__61_;
      r_228__60_ <= r_n_228__60_;
      r_228__59_ <= r_n_228__59_;
      r_228__58_ <= r_n_228__58_;
      r_228__57_ <= r_n_228__57_;
      r_228__56_ <= r_n_228__56_;
      r_228__55_ <= r_n_228__55_;
      r_228__54_ <= r_n_228__54_;
      r_228__53_ <= r_n_228__53_;
      r_228__52_ <= r_n_228__52_;
      r_228__51_ <= r_n_228__51_;
      r_228__50_ <= r_n_228__50_;
      r_228__49_ <= r_n_228__49_;
      r_228__48_ <= r_n_228__48_;
      r_228__47_ <= r_n_228__47_;
      r_228__46_ <= r_n_228__46_;
      r_228__45_ <= r_n_228__45_;
      r_228__44_ <= r_n_228__44_;
      r_228__43_ <= r_n_228__43_;
      r_228__42_ <= r_n_228__42_;
      r_228__41_ <= r_n_228__41_;
      r_228__40_ <= r_n_228__40_;
      r_228__39_ <= r_n_228__39_;
      r_228__38_ <= r_n_228__38_;
      r_228__37_ <= r_n_228__37_;
      r_228__36_ <= r_n_228__36_;
      r_228__35_ <= r_n_228__35_;
      r_228__34_ <= r_n_228__34_;
      r_228__33_ <= r_n_228__33_;
      r_228__32_ <= r_n_228__32_;
      r_228__31_ <= r_n_228__31_;
      r_228__30_ <= r_n_228__30_;
      r_228__29_ <= r_n_228__29_;
      r_228__28_ <= r_n_228__28_;
      r_228__27_ <= r_n_228__27_;
      r_228__26_ <= r_n_228__26_;
      r_228__25_ <= r_n_228__25_;
      r_228__24_ <= r_n_228__24_;
      r_228__23_ <= r_n_228__23_;
      r_228__22_ <= r_n_228__22_;
      r_228__21_ <= r_n_228__21_;
      r_228__20_ <= r_n_228__20_;
      r_228__19_ <= r_n_228__19_;
      r_228__18_ <= r_n_228__18_;
      r_228__17_ <= r_n_228__17_;
      r_228__16_ <= r_n_228__16_;
      r_228__15_ <= r_n_228__15_;
      r_228__14_ <= r_n_228__14_;
      r_228__13_ <= r_n_228__13_;
      r_228__12_ <= r_n_228__12_;
      r_228__11_ <= r_n_228__11_;
      r_228__10_ <= r_n_228__10_;
      r_228__9_ <= r_n_228__9_;
      r_228__8_ <= r_n_228__8_;
      r_228__7_ <= r_n_228__7_;
      r_228__6_ <= r_n_228__6_;
      r_228__5_ <= r_n_228__5_;
      r_228__4_ <= r_n_228__4_;
      r_228__3_ <= r_n_228__3_;
      r_228__2_ <= r_n_228__2_;
      r_228__1_ <= r_n_228__1_;
      r_228__0_ <= r_n_228__0_;
    end 
    if(N3813) begin
      r_229__63_ <= r_n_229__63_;
      r_229__62_ <= r_n_229__62_;
      r_229__61_ <= r_n_229__61_;
      r_229__60_ <= r_n_229__60_;
      r_229__59_ <= r_n_229__59_;
      r_229__58_ <= r_n_229__58_;
      r_229__57_ <= r_n_229__57_;
      r_229__56_ <= r_n_229__56_;
      r_229__55_ <= r_n_229__55_;
      r_229__54_ <= r_n_229__54_;
      r_229__53_ <= r_n_229__53_;
      r_229__52_ <= r_n_229__52_;
      r_229__51_ <= r_n_229__51_;
      r_229__50_ <= r_n_229__50_;
      r_229__49_ <= r_n_229__49_;
      r_229__48_ <= r_n_229__48_;
      r_229__47_ <= r_n_229__47_;
      r_229__46_ <= r_n_229__46_;
      r_229__45_ <= r_n_229__45_;
      r_229__44_ <= r_n_229__44_;
      r_229__43_ <= r_n_229__43_;
      r_229__42_ <= r_n_229__42_;
      r_229__41_ <= r_n_229__41_;
      r_229__40_ <= r_n_229__40_;
      r_229__39_ <= r_n_229__39_;
      r_229__38_ <= r_n_229__38_;
      r_229__37_ <= r_n_229__37_;
      r_229__36_ <= r_n_229__36_;
      r_229__35_ <= r_n_229__35_;
      r_229__34_ <= r_n_229__34_;
      r_229__33_ <= r_n_229__33_;
      r_229__32_ <= r_n_229__32_;
      r_229__31_ <= r_n_229__31_;
      r_229__30_ <= r_n_229__30_;
      r_229__29_ <= r_n_229__29_;
      r_229__28_ <= r_n_229__28_;
      r_229__27_ <= r_n_229__27_;
      r_229__26_ <= r_n_229__26_;
      r_229__25_ <= r_n_229__25_;
      r_229__24_ <= r_n_229__24_;
      r_229__23_ <= r_n_229__23_;
      r_229__22_ <= r_n_229__22_;
      r_229__21_ <= r_n_229__21_;
      r_229__20_ <= r_n_229__20_;
      r_229__19_ <= r_n_229__19_;
      r_229__18_ <= r_n_229__18_;
      r_229__17_ <= r_n_229__17_;
      r_229__16_ <= r_n_229__16_;
      r_229__15_ <= r_n_229__15_;
      r_229__14_ <= r_n_229__14_;
      r_229__13_ <= r_n_229__13_;
      r_229__12_ <= r_n_229__12_;
      r_229__11_ <= r_n_229__11_;
      r_229__10_ <= r_n_229__10_;
      r_229__9_ <= r_n_229__9_;
      r_229__8_ <= r_n_229__8_;
      r_229__7_ <= r_n_229__7_;
      r_229__6_ <= r_n_229__6_;
      r_229__5_ <= r_n_229__5_;
      r_229__4_ <= r_n_229__4_;
      r_229__3_ <= r_n_229__3_;
      r_229__2_ <= r_n_229__2_;
      r_229__1_ <= r_n_229__1_;
      r_229__0_ <= r_n_229__0_;
    end 
    if(N3814) begin
      r_230__63_ <= r_n_230__63_;
      r_230__62_ <= r_n_230__62_;
      r_230__61_ <= r_n_230__61_;
      r_230__60_ <= r_n_230__60_;
      r_230__59_ <= r_n_230__59_;
      r_230__58_ <= r_n_230__58_;
      r_230__57_ <= r_n_230__57_;
      r_230__56_ <= r_n_230__56_;
      r_230__55_ <= r_n_230__55_;
      r_230__54_ <= r_n_230__54_;
      r_230__53_ <= r_n_230__53_;
      r_230__52_ <= r_n_230__52_;
      r_230__51_ <= r_n_230__51_;
      r_230__50_ <= r_n_230__50_;
      r_230__49_ <= r_n_230__49_;
      r_230__48_ <= r_n_230__48_;
      r_230__47_ <= r_n_230__47_;
      r_230__46_ <= r_n_230__46_;
      r_230__45_ <= r_n_230__45_;
      r_230__44_ <= r_n_230__44_;
      r_230__43_ <= r_n_230__43_;
      r_230__42_ <= r_n_230__42_;
      r_230__41_ <= r_n_230__41_;
      r_230__40_ <= r_n_230__40_;
      r_230__39_ <= r_n_230__39_;
      r_230__38_ <= r_n_230__38_;
      r_230__37_ <= r_n_230__37_;
      r_230__36_ <= r_n_230__36_;
      r_230__35_ <= r_n_230__35_;
      r_230__34_ <= r_n_230__34_;
      r_230__33_ <= r_n_230__33_;
      r_230__32_ <= r_n_230__32_;
      r_230__31_ <= r_n_230__31_;
      r_230__30_ <= r_n_230__30_;
      r_230__29_ <= r_n_230__29_;
      r_230__28_ <= r_n_230__28_;
      r_230__27_ <= r_n_230__27_;
      r_230__26_ <= r_n_230__26_;
      r_230__25_ <= r_n_230__25_;
      r_230__24_ <= r_n_230__24_;
      r_230__23_ <= r_n_230__23_;
      r_230__22_ <= r_n_230__22_;
      r_230__21_ <= r_n_230__21_;
      r_230__20_ <= r_n_230__20_;
      r_230__19_ <= r_n_230__19_;
      r_230__18_ <= r_n_230__18_;
      r_230__17_ <= r_n_230__17_;
      r_230__16_ <= r_n_230__16_;
      r_230__15_ <= r_n_230__15_;
      r_230__14_ <= r_n_230__14_;
      r_230__13_ <= r_n_230__13_;
      r_230__12_ <= r_n_230__12_;
      r_230__11_ <= r_n_230__11_;
      r_230__10_ <= r_n_230__10_;
      r_230__9_ <= r_n_230__9_;
      r_230__8_ <= r_n_230__8_;
      r_230__7_ <= r_n_230__7_;
      r_230__6_ <= r_n_230__6_;
      r_230__5_ <= r_n_230__5_;
      r_230__4_ <= r_n_230__4_;
      r_230__3_ <= r_n_230__3_;
      r_230__2_ <= r_n_230__2_;
      r_230__1_ <= r_n_230__1_;
      r_230__0_ <= r_n_230__0_;
    end 
    if(N3815) begin
      r_231__63_ <= r_n_231__63_;
      r_231__62_ <= r_n_231__62_;
      r_231__61_ <= r_n_231__61_;
      r_231__60_ <= r_n_231__60_;
      r_231__59_ <= r_n_231__59_;
      r_231__58_ <= r_n_231__58_;
      r_231__57_ <= r_n_231__57_;
      r_231__56_ <= r_n_231__56_;
      r_231__55_ <= r_n_231__55_;
      r_231__54_ <= r_n_231__54_;
      r_231__53_ <= r_n_231__53_;
      r_231__52_ <= r_n_231__52_;
      r_231__51_ <= r_n_231__51_;
      r_231__50_ <= r_n_231__50_;
      r_231__49_ <= r_n_231__49_;
      r_231__48_ <= r_n_231__48_;
      r_231__47_ <= r_n_231__47_;
      r_231__46_ <= r_n_231__46_;
      r_231__45_ <= r_n_231__45_;
      r_231__44_ <= r_n_231__44_;
      r_231__43_ <= r_n_231__43_;
      r_231__42_ <= r_n_231__42_;
      r_231__41_ <= r_n_231__41_;
      r_231__40_ <= r_n_231__40_;
      r_231__39_ <= r_n_231__39_;
      r_231__38_ <= r_n_231__38_;
      r_231__37_ <= r_n_231__37_;
      r_231__36_ <= r_n_231__36_;
      r_231__35_ <= r_n_231__35_;
      r_231__34_ <= r_n_231__34_;
      r_231__33_ <= r_n_231__33_;
      r_231__32_ <= r_n_231__32_;
      r_231__31_ <= r_n_231__31_;
      r_231__30_ <= r_n_231__30_;
      r_231__29_ <= r_n_231__29_;
      r_231__28_ <= r_n_231__28_;
      r_231__27_ <= r_n_231__27_;
      r_231__26_ <= r_n_231__26_;
      r_231__25_ <= r_n_231__25_;
      r_231__24_ <= r_n_231__24_;
      r_231__23_ <= r_n_231__23_;
      r_231__22_ <= r_n_231__22_;
      r_231__21_ <= r_n_231__21_;
      r_231__20_ <= r_n_231__20_;
      r_231__19_ <= r_n_231__19_;
      r_231__18_ <= r_n_231__18_;
      r_231__17_ <= r_n_231__17_;
      r_231__16_ <= r_n_231__16_;
      r_231__15_ <= r_n_231__15_;
      r_231__14_ <= r_n_231__14_;
      r_231__13_ <= r_n_231__13_;
      r_231__12_ <= r_n_231__12_;
      r_231__11_ <= r_n_231__11_;
      r_231__10_ <= r_n_231__10_;
      r_231__9_ <= r_n_231__9_;
      r_231__8_ <= r_n_231__8_;
      r_231__7_ <= r_n_231__7_;
      r_231__6_ <= r_n_231__6_;
      r_231__5_ <= r_n_231__5_;
      r_231__4_ <= r_n_231__4_;
      r_231__3_ <= r_n_231__3_;
      r_231__2_ <= r_n_231__2_;
      r_231__1_ <= r_n_231__1_;
      r_231__0_ <= r_n_231__0_;
    end 
    if(N3816) begin
      r_232__63_ <= r_n_232__63_;
      r_232__62_ <= r_n_232__62_;
      r_232__61_ <= r_n_232__61_;
      r_232__60_ <= r_n_232__60_;
      r_232__59_ <= r_n_232__59_;
      r_232__58_ <= r_n_232__58_;
      r_232__57_ <= r_n_232__57_;
      r_232__56_ <= r_n_232__56_;
      r_232__55_ <= r_n_232__55_;
      r_232__54_ <= r_n_232__54_;
      r_232__53_ <= r_n_232__53_;
      r_232__52_ <= r_n_232__52_;
      r_232__51_ <= r_n_232__51_;
      r_232__50_ <= r_n_232__50_;
      r_232__49_ <= r_n_232__49_;
      r_232__48_ <= r_n_232__48_;
      r_232__47_ <= r_n_232__47_;
      r_232__46_ <= r_n_232__46_;
      r_232__45_ <= r_n_232__45_;
      r_232__44_ <= r_n_232__44_;
      r_232__43_ <= r_n_232__43_;
      r_232__42_ <= r_n_232__42_;
      r_232__41_ <= r_n_232__41_;
      r_232__40_ <= r_n_232__40_;
      r_232__39_ <= r_n_232__39_;
      r_232__38_ <= r_n_232__38_;
      r_232__37_ <= r_n_232__37_;
      r_232__36_ <= r_n_232__36_;
      r_232__35_ <= r_n_232__35_;
      r_232__34_ <= r_n_232__34_;
      r_232__33_ <= r_n_232__33_;
      r_232__32_ <= r_n_232__32_;
      r_232__31_ <= r_n_232__31_;
      r_232__30_ <= r_n_232__30_;
      r_232__29_ <= r_n_232__29_;
      r_232__28_ <= r_n_232__28_;
      r_232__27_ <= r_n_232__27_;
      r_232__26_ <= r_n_232__26_;
      r_232__25_ <= r_n_232__25_;
      r_232__24_ <= r_n_232__24_;
      r_232__23_ <= r_n_232__23_;
      r_232__22_ <= r_n_232__22_;
      r_232__21_ <= r_n_232__21_;
      r_232__20_ <= r_n_232__20_;
      r_232__19_ <= r_n_232__19_;
      r_232__18_ <= r_n_232__18_;
      r_232__17_ <= r_n_232__17_;
      r_232__16_ <= r_n_232__16_;
      r_232__15_ <= r_n_232__15_;
      r_232__14_ <= r_n_232__14_;
      r_232__13_ <= r_n_232__13_;
      r_232__12_ <= r_n_232__12_;
      r_232__11_ <= r_n_232__11_;
      r_232__10_ <= r_n_232__10_;
      r_232__9_ <= r_n_232__9_;
      r_232__8_ <= r_n_232__8_;
      r_232__7_ <= r_n_232__7_;
      r_232__6_ <= r_n_232__6_;
      r_232__5_ <= r_n_232__5_;
      r_232__4_ <= r_n_232__4_;
      r_232__3_ <= r_n_232__3_;
      r_232__2_ <= r_n_232__2_;
      r_232__1_ <= r_n_232__1_;
      r_232__0_ <= r_n_232__0_;
    end 
    if(N3817) begin
      r_233__63_ <= r_n_233__63_;
      r_233__62_ <= r_n_233__62_;
      r_233__61_ <= r_n_233__61_;
      r_233__60_ <= r_n_233__60_;
      r_233__59_ <= r_n_233__59_;
      r_233__58_ <= r_n_233__58_;
      r_233__57_ <= r_n_233__57_;
      r_233__56_ <= r_n_233__56_;
      r_233__55_ <= r_n_233__55_;
      r_233__54_ <= r_n_233__54_;
      r_233__53_ <= r_n_233__53_;
      r_233__52_ <= r_n_233__52_;
      r_233__51_ <= r_n_233__51_;
      r_233__50_ <= r_n_233__50_;
      r_233__49_ <= r_n_233__49_;
      r_233__48_ <= r_n_233__48_;
      r_233__47_ <= r_n_233__47_;
      r_233__46_ <= r_n_233__46_;
      r_233__45_ <= r_n_233__45_;
      r_233__44_ <= r_n_233__44_;
      r_233__43_ <= r_n_233__43_;
      r_233__42_ <= r_n_233__42_;
      r_233__41_ <= r_n_233__41_;
      r_233__40_ <= r_n_233__40_;
      r_233__39_ <= r_n_233__39_;
      r_233__38_ <= r_n_233__38_;
      r_233__37_ <= r_n_233__37_;
      r_233__36_ <= r_n_233__36_;
      r_233__35_ <= r_n_233__35_;
      r_233__34_ <= r_n_233__34_;
      r_233__33_ <= r_n_233__33_;
      r_233__32_ <= r_n_233__32_;
      r_233__31_ <= r_n_233__31_;
      r_233__30_ <= r_n_233__30_;
      r_233__29_ <= r_n_233__29_;
      r_233__28_ <= r_n_233__28_;
      r_233__27_ <= r_n_233__27_;
      r_233__26_ <= r_n_233__26_;
      r_233__25_ <= r_n_233__25_;
      r_233__24_ <= r_n_233__24_;
      r_233__23_ <= r_n_233__23_;
      r_233__22_ <= r_n_233__22_;
      r_233__21_ <= r_n_233__21_;
      r_233__20_ <= r_n_233__20_;
      r_233__19_ <= r_n_233__19_;
      r_233__18_ <= r_n_233__18_;
      r_233__17_ <= r_n_233__17_;
      r_233__16_ <= r_n_233__16_;
      r_233__15_ <= r_n_233__15_;
      r_233__14_ <= r_n_233__14_;
      r_233__13_ <= r_n_233__13_;
      r_233__12_ <= r_n_233__12_;
      r_233__11_ <= r_n_233__11_;
      r_233__10_ <= r_n_233__10_;
      r_233__9_ <= r_n_233__9_;
      r_233__8_ <= r_n_233__8_;
      r_233__7_ <= r_n_233__7_;
      r_233__6_ <= r_n_233__6_;
      r_233__5_ <= r_n_233__5_;
      r_233__4_ <= r_n_233__4_;
      r_233__3_ <= r_n_233__3_;
      r_233__2_ <= r_n_233__2_;
      r_233__1_ <= r_n_233__1_;
      r_233__0_ <= r_n_233__0_;
    end 
    if(N3818) begin
      r_234__63_ <= r_n_234__63_;
      r_234__62_ <= r_n_234__62_;
      r_234__61_ <= r_n_234__61_;
      r_234__60_ <= r_n_234__60_;
      r_234__59_ <= r_n_234__59_;
      r_234__58_ <= r_n_234__58_;
      r_234__57_ <= r_n_234__57_;
      r_234__56_ <= r_n_234__56_;
      r_234__55_ <= r_n_234__55_;
      r_234__54_ <= r_n_234__54_;
      r_234__53_ <= r_n_234__53_;
      r_234__52_ <= r_n_234__52_;
      r_234__51_ <= r_n_234__51_;
      r_234__50_ <= r_n_234__50_;
      r_234__49_ <= r_n_234__49_;
      r_234__48_ <= r_n_234__48_;
      r_234__47_ <= r_n_234__47_;
      r_234__46_ <= r_n_234__46_;
      r_234__45_ <= r_n_234__45_;
      r_234__44_ <= r_n_234__44_;
      r_234__43_ <= r_n_234__43_;
      r_234__42_ <= r_n_234__42_;
      r_234__41_ <= r_n_234__41_;
      r_234__40_ <= r_n_234__40_;
      r_234__39_ <= r_n_234__39_;
      r_234__38_ <= r_n_234__38_;
      r_234__37_ <= r_n_234__37_;
      r_234__36_ <= r_n_234__36_;
      r_234__35_ <= r_n_234__35_;
      r_234__34_ <= r_n_234__34_;
      r_234__33_ <= r_n_234__33_;
      r_234__32_ <= r_n_234__32_;
      r_234__31_ <= r_n_234__31_;
      r_234__30_ <= r_n_234__30_;
      r_234__29_ <= r_n_234__29_;
      r_234__28_ <= r_n_234__28_;
      r_234__27_ <= r_n_234__27_;
      r_234__26_ <= r_n_234__26_;
      r_234__25_ <= r_n_234__25_;
      r_234__24_ <= r_n_234__24_;
      r_234__23_ <= r_n_234__23_;
      r_234__22_ <= r_n_234__22_;
      r_234__21_ <= r_n_234__21_;
      r_234__20_ <= r_n_234__20_;
      r_234__19_ <= r_n_234__19_;
      r_234__18_ <= r_n_234__18_;
      r_234__17_ <= r_n_234__17_;
      r_234__16_ <= r_n_234__16_;
      r_234__15_ <= r_n_234__15_;
      r_234__14_ <= r_n_234__14_;
      r_234__13_ <= r_n_234__13_;
      r_234__12_ <= r_n_234__12_;
      r_234__11_ <= r_n_234__11_;
      r_234__10_ <= r_n_234__10_;
      r_234__9_ <= r_n_234__9_;
      r_234__8_ <= r_n_234__8_;
      r_234__7_ <= r_n_234__7_;
      r_234__6_ <= r_n_234__6_;
      r_234__5_ <= r_n_234__5_;
      r_234__4_ <= r_n_234__4_;
      r_234__3_ <= r_n_234__3_;
      r_234__2_ <= r_n_234__2_;
      r_234__1_ <= r_n_234__1_;
      r_234__0_ <= r_n_234__0_;
    end 
    if(N3819) begin
      r_235__63_ <= r_n_235__63_;
      r_235__62_ <= r_n_235__62_;
      r_235__61_ <= r_n_235__61_;
      r_235__60_ <= r_n_235__60_;
      r_235__59_ <= r_n_235__59_;
      r_235__58_ <= r_n_235__58_;
      r_235__57_ <= r_n_235__57_;
      r_235__56_ <= r_n_235__56_;
      r_235__55_ <= r_n_235__55_;
      r_235__54_ <= r_n_235__54_;
      r_235__53_ <= r_n_235__53_;
      r_235__52_ <= r_n_235__52_;
      r_235__51_ <= r_n_235__51_;
      r_235__50_ <= r_n_235__50_;
      r_235__49_ <= r_n_235__49_;
      r_235__48_ <= r_n_235__48_;
      r_235__47_ <= r_n_235__47_;
      r_235__46_ <= r_n_235__46_;
      r_235__45_ <= r_n_235__45_;
      r_235__44_ <= r_n_235__44_;
      r_235__43_ <= r_n_235__43_;
      r_235__42_ <= r_n_235__42_;
      r_235__41_ <= r_n_235__41_;
      r_235__40_ <= r_n_235__40_;
      r_235__39_ <= r_n_235__39_;
      r_235__38_ <= r_n_235__38_;
      r_235__37_ <= r_n_235__37_;
      r_235__36_ <= r_n_235__36_;
      r_235__35_ <= r_n_235__35_;
      r_235__34_ <= r_n_235__34_;
      r_235__33_ <= r_n_235__33_;
      r_235__32_ <= r_n_235__32_;
      r_235__31_ <= r_n_235__31_;
      r_235__30_ <= r_n_235__30_;
      r_235__29_ <= r_n_235__29_;
      r_235__28_ <= r_n_235__28_;
      r_235__27_ <= r_n_235__27_;
      r_235__26_ <= r_n_235__26_;
      r_235__25_ <= r_n_235__25_;
      r_235__24_ <= r_n_235__24_;
      r_235__23_ <= r_n_235__23_;
      r_235__22_ <= r_n_235__22_;
      r_235__21_ <= r_n_235__21_;
      r_235__20_ <= r_n_235__20_;
      r_235__19_ <= r_n_235__19_;
      r_235__18_ <= r_n_235__18_;
      r_235__17_ <= r_n_235__17_;
      r_235__16_ <= r_n_235__16_;
      r_235__15_ <= r_n_235__15_;
      r_235__14_ <= r_n_235__14_;
      r_235__13_ <= r_n_235__13_;
      r_235__12_ <= r_n_235__12_;
      r_235__11_ <= r_n_235__11_;
      r_235__10_ <= r_n_235__10_;
      r_235__9_ <= r_n_235__9_;
      r_235__8_ <= r_n_235__8_;
      r_235__7_ <= r_n_235__7_;
      r_235__6_ <= r_n_235__6_;
      r_235__5_ <= r_n_235__5_;
      r_235__4_ <= r_n_235__4_;
      r_235__3_ <= r_n_235__3_;
      r_235__2_ <= r_n_235__2_;
      r_235__1_ <= r_n_235__1_;
      r_235__0_ <= r_n_235__0_;
    end 
    if(N3820) begin
      r_236__63_ <= r_n_236__63_;
      r_236__62_ <= r_n_236__62_;
      r_236__61_ <= r_n_236__61_;
      r_236__60_ <= r_n_236__60_;
      r_236__59_ <= r_n_236__59_;
      r_236__58_ <= r_n_236__58_;
      r_236__57_ <= r_n_236__57_;
      r_236__56_ <= r_n_236__56_;
      r_236__55_ <= r_n_236__55_;
      r_236__54_ <= r_n_236__54_;
      r_236__53_ <= r_n_236__53_;
      r_236__52_ <= r_n_236__52_;
      r_236__51_ <= r_n_236__51_;
      r_236__50_ <= r_n_236__50_;
      r_236__49_ <= r_n_236__49_;
      r_236__48_ <= r_n_236__48_;
      r_236__47_ <= r_n_236__47_;
      r_236__46_ <= r_n_236__46_;
      r_236__45_ <= r_n_236__45_;
      r_236__44_ <= r_n_236__44_;
      r_236__43_ <= r_n_236__43_;
      r_236__42_ <= r_n_236__42_;
      r_236__41_ <= r_n_236__41_;
      r_236__40_ <= r_n_236__40_;
      r_236__39_ <= r_n_236__39_;
      r_236__38_ <= r_n_236__38_;
      r_236__37_ <= r_n_236__37_;
      r_236__36_ <= r_n_236__36_;
      r_236__35_ <= r_n_236__35_;
      r_236__34_ <= r_n_236__34_;
      r_236__33_ <= r_n_236__33_;
      r_236__32_ <= r_n_236__32_;
      r_236__31_ <= r_n_236__31_;
      r_236__30_ <= r_n_236__30_;
      r_236__29_ <= r_n_236__29_;
      r_236__28_ <= r_n_236__28_;
      r_236__27_ <= r_n_236__27_;
      r_236__26_ <= r_n_236__26_;
      r_236__25_ <= r_n_236__25_;
      r_236__24_ <= r_n_236__24_;
      r_236__23_ <= r_n_236__23_;
      r_236__22_ <= r_n_236__22_;
      r_236__21_ <= r_n_236__21_;
      r_236__20_ <= r_n_236__20_;
      r_236__19_ <= r_n_236__19_;
      r_236__18_ <= r_n_236__18_;
      r_236__17_ <= r_n_236__17_;
      r_236__16_ <= r_n_236__16_;
      r_236__15_ <= r_n_236__15_;
      r_236__14_ <= r_n_236__14_;
      r_236__13_ <= r_n_236__13_;
      r_236__12_ <= r_n_236__12_;
      r_236__11_ <= r_n_236__11_;
      r_236__10_ <= r_n_236__10_;
      r_236__9_ <= r_n_236__9_;
      r_236__8_ <= r_n_236__8_;
      r_236__7_ <= r_n_236__7_;
      r_236__6_ <= r_n_236__6_;
      r_236__5_ <= r_n_236__5_;
      r_236__4_ <= r_n_236__4_;
      r_236__3_ <= r_n_236__3_;
      r_236__2_ <= r_n_236__2_;
      r_236__1_ <= r_n_236__1_;
      r_236__0_ <= r_n_236__0_;
    end 
    if(N3821) begin
      r_237__63_ <= r_n_237__63_;
      r_237__62_ <= r_n_237__62_;
      r_237__61_ <= r_n_237__61_;
      r_237__60_ <= r_n_237__60_;
      r_237__59_ <= r_n_237__59_;
      r_237__58_ <= r_n_237__58_;
      r_237__57_ <= r_n_237__57_;
      r_237__56_ <= r_n_237__56_;
      r_237__55_ <= r_n_237__55_;
      r_237__54_ <= r_n_237__54_;
      r_237__53_ <= r_n_237__53_;
      r_237__52_ <= r_n_237__52_;
      r_237__51_ <= r_n_237__51_;
      r_237__50_ <= r_n_237__50_;
      r_237__49_ <= r_n_237__49_;
      r_237__48_ <= r_n_237__48_;
      r_237__47_ <= r_n_237__47_;
      r_237__46_ <= r_n_237__46_;
      r_237__45_ <= r_n_237__45_;
      r_237__44_ <= r_n_237__44_;
      r_237__43_ <= r_n_237__43_;
      r_237__42_ <= r_n_237__42_;
      r_237__41_ <= r_n_237__41_;
      r_237__40_ <= r_n_237__40_;
      r_237__39_ <= r_n_237__39_;
      r_237__38_ <= r_n_237__38_;
      r_237__37_ <= r_n_237__37_;
      r_237__36_ <= r_n_237__36_;
      r_237__35_ <= r_n_237__35_;
      r_237__34_ <= r_n_237__34_;
      r_237__33_ <= r_n_237__33_;
      r_237__32_ <= r_n_237__32_;
      r_237__31_ <= r_n_237__31_;
      r_237__30_ <= r_n_237__30_;
      r_237__29_ <= r_n_237__29_;
      r_237__28_ <= r_n_237__28_;
      r_237__27_ <= r_n_237__27_;
      r_237__26_ <= r_n_237__26_;
      r_237__25_ <= r_n_237__25_;
      r_237__24_ <= r_n_237__24_;
      r_237__23_ <= r_n_237__23_;
      r_237__22_ <= r_n_237__22_;
      r_237__21_ <= r_n_237__21_;
      r_237__20_ <= r_n_237__20_;
      r_237__19_ <= r_n_237__19_;
      r_237__18_ <= r_n_237__18_;
      r_237__17_ <= r_n_237__17_;
      r_237__16_ <= r_n_237__16_;
      r_237__15_ <= r_n_237__15_;
      r_237__14_ <= r_n_237__14_;
      r_237__13_ <= r_n_237__13_;
      r_237__12_ <= r_n_237__12_;
      r_237__11_ <= r_n_237__11_;
      r_237__10_ <= r_n_237__10_;
      r_237__9_ <= r_n_237__9_;
      r_237__8_ <= r_n_237__8_;
      r_237__7_ <= r_n_237__7_;
      r_237__6_ <= r_n_237__6_;
      r_237__5_ <= r_n_237__5_;
      r_237__4_ <= r_n_237__4_;
      r_237__3_ <= r_n_237__3_;
      r_237__2_ <= r_n_237__2_;
      r_237__1_ <= r_n_237__1_;
      r_237__0_ <= r_n_237__0_;
    end 
    if(N3822) begin
      r_238__63_ <= r_n_238__63_;
      r_238__62_ <= r_n_238__62_;
      r_238__61_ <= r_n_238__61_;
      r_238__60_ <= r_n_238__60_;
      r_238__59_ <= r_n_238__59_;
      r_238__58_ <= r_n_238__58_;
      r_238__57_ <= r_n_238__57_;
      r_238__56_ <= r_n_238__56_;
      r_238__55_ <= r_n_238__55_;
      r_238__54_ <= r_n_238__54_;
      r_238__53_ <= r_n_238__53_;
      r_238__52_ <= r_n_238__52_;
      r_238__51_ <= r_n_238__51_;
      r_238__50_ <= r_n_238__50_;
      r_238__49_ <= r_n_238__49_;
      r_238__48_ <= r_n_238__48_;
      r_238__47_ <= r_n_238__47_;
      r_238__46_ <= r_n_238__46_;
      r_238__45_ <= r_n_238__45_;
      r_238__44_ <= r_n_238__44_;
      r_238__43_ <= r_n_238__43_;
      r_238__42_ <= r_n_238__42_;
      r_238__41_ <= r_n_238__41_;
      r_238__40_ <= r_n_238__40_;
      r_238__39_ <= r_n_238__39_;
      r_238__38_ <= r_n_238__38_;
      r_238__37_ <= r_n_238__37_;
      r_238__36_ <= r_n_238__36_;
      r_238__35_ <= r_n_238__35_;
      r_238__34_ <= r_n_238__34_;
      r_238__33_ <= r_n_238__33_;
      r_238__32_ <= r_n_238__32_;
      r_238__31_ <= r_n_238__31_;
      r_238__30_ <= r_n_238__30_;
      r_238__29_ <= r_n_238__29_;
      r_238__28_ <= r_n_238__28_;
      r_238__27_ <= r_n_238__27_;
      r_238__26_ <= r_n_238__26_;
      r_238__25_ <= r_n_238__25_;
      r_238__24_ <= r_n_238__24_;
      r_238__23_ <= r_n_238__23_;
      r_238__22_ <= r_n_238__22_;
      r_238__21_ <= r_n_238__21_;
      r_238__20_ <= r_n_238__20_;
      r_238__19_ <= r_n_238__19_;
      r_238__18_ <= r_n_238__18_;
      r_238__17_ <= r_n_238__17_;
      r_238__16_ <= r_n_238__16_;
      r_238__15_ <= r_n_238__15_;
      r_238__14_ <= r_n_238__14_;
      r_238__13_ <= r_n_238__13_;
      r_238__12_ <= r_n_238__12_;
      r_238__11_ <= r_n_238__11_;
      r_238__10_ <= r_n_238__10_;
      r_238__9_ <= r_n_238__9_;
      r_238__8_ <= r_n_238__8_;
      r_238__7_ <= r_n_238__7_;
      r_238__6_ <= r_n_238__6_;
      r_238__5_ <= r_n_238__5_;
      r_238__4_ <= r_n_238__4_;
      r_238__3_ <= r_n_238__3_;
      r_238__2_ <= r_n_238__2_;
      r_238__1_ <= r_n_238__1_;
      r_238__0_ <= r_n_238__0_;
    end 
    if(N3823) begin
      r_239__63_ <= r_n_239__63_;
      r_239__62_ <= r_n_239__62_;
      r_239__61_ <= r_n_239__61_;
      r_239__60_ <= r_n_239__60_;
      r_239__59_ <= r_n_239__59_;
      r_239__58_ <= r_n_239__58_;
      r_239__57_ <= r_n_239__57_;
      r_239__56_ <= r_n_239__56_;
      r_239__55_ <= r_n_239__55_;
      r_239__54_ <= r_n_239__54_;
      r_239__53_ <= r_n_239__53_;
      r_239__52_ <= r_n_239__52_;
      r_239__51_ <= r_n_239__51_;
      r_239__50_ <= r_n_239__50_;
      r_239__49_ <= r_n_239__49_;
      r_239__48_ <= r_n_239__48_;
      r_239__47_ <= r_n_239__47_;
      r_239__46_ <= r_n_239__46_;
      r_239__45_ <= r_n_239__45_;
      r_239__44_ <= r_n_239__44_;
      r_239__43_ <= r_n_239__43_;
      r_239__42_ <= r_n_239__42_;
      r_239__41_ <= r_n_239__41_;
      r_239__40_ <= r_n_239__40_;
      r_239__39_ <= r_n_239__39_;
      r_239__38_ <= r_n_239__38_;
      r_239__37_ <= r_n_239__37_;
      r_239__36_ <= r_n_239__36_;
      r_239__35_ <= r_n_239__35_;
      r_239__34_ <= r_n_239__34_;
      r_239__33_ <= r_n_239__33_;
      r_239__32_ <= r_n_239__32_;
      r_239__31_ <= r_n_239__31_;
      r_239__30_ <= r_n_239__30_;
      r_239__29_ <= r_n_239__29_;
      r_239__28_ <= r_n_239__28_;
      r_239__27_ <= r_n_239__27_;
      r_239__26_ <= r_n_239__26_;
      r_239__25_ <= r_n_239__25_;
      r_239__24_ <= r_n_239__24_;
      r_239__23_ <= r_n_239__23_;
      r_239__22_ <= r_n_239__22_;
      r_239__21_ <= r_n_239__21_;
      r_239__20_ <= r_n_239__20_;
      r_239__19_ <= r_n_239__19_;
      r_239__18_ <= r_n_239__18_;
      r_239__17_ <= r_n_239__17_;
      r_239__16_ <= r_n_239__16_;
      r_239__15_ <= r_n_239__15_;
      r_239__14_ <= r_n_239__14_;
      r_239__13_ <= r_n_239__13_;
      r_239__12_ <= r_n_239__12_;
      r_239__11_ <= r_n_239__11_;
      r_239__10_ <= r_n_239__10_;
      r_239__9_ <= r_n_239__9_;
      r_239__8_ <= r_n_239__8_;
      r_239__7_ <= r_n_239__7_;
      r_239__6_ <= r_n_239__6_;
      r_239__5_ <= r_n_239__5_;
      r_239__4_ <= r_n_239__4_;
      r_239__3_ <= r_n_239__3_;
      r_239__2_ <= r_n_239__2_;
      r_239__1_ <= r_n_239__1_;
      r_239__0_ <= r_n_239__0_;
    end 
    if(N3824) begin
      r_240__63_ <= r_n_240__63_;
      r_240__62_ <= r_n_240__62_;
      r_240__61_ <= r_n_240__61_;
      r_240__60_ <= r_n_240__60_;
      r_240__59_ <= r_n_240__59_;
      r_240__58_ <= r_n_240__58_;
      r_240__57_ <= r_n_240__57_;
      r_240__56_ <= r_n_240__56_;
      r_240__55_ <= r_n_240__55_;
      r_240__54_ <= r_n_240__54_;
      r_240__53_ <= r_n_240__53_;
      r_240__52_ <= r_n_240__52_;
      r_240__51_ <= r_n_240__51_;
      r_240__50_ <= r_n_240__50_;
      r_240__49_ <= r_n_240__49_;
      r_240__48_ <= r_n_240__48_;
      r_240__47_ <= r_n_240__47_;
      r_240__46_ <= r_n_240__46_;
      r_240__45_ <= r_n_240__45_;
      r_240__44_ <= r_n_240__44_;
      r_240__43_ <= r_n_240__43_;
      r_240__42_ <= r_n_240__42_;
      r_240__41_ <= r_n_240__41_;
      r_240__40_ <= r_n_240__40_;
      r_240__39_ <= r_n_240__39_;
      r_240__38_ <= r_n_240__38_;
      r_240__37_ <= r_n_240__37_;
      r_240__36_ <= r_n_240__36_;
      r_240__35_ <= r_n_240__35_;
      r_240__34_ <= r_n_240__34_;
      r_240__33_ <= r_n_240__33_;
      r_240__32_ <= r_n_240__32_;
      r_240__31_ <= r_n_240__31_;
      r_240__30_ <= r_n_240__30_;
      r_240__29_ <= r_n_240__29_;
      r_240__28_ <= r_n_240__28_;
      r_240__27_ <= r_n_240__27_;
      r_240__26_ <= r_n_240__26_;
      r_240__25_ <= r_n_240__25_;
      r_240__24_ <= r_n_240__24_;
      r_240__23_ <= r_n_240__23_;
      r_240__22_ <= r_n_240__22_;
      r_240__21_ <= r_n_240__21_;
      r_240__20_ <= r_n_240__20_;
      r_240__19_ <= r_n_240__19_;
      r_240__18_ <= r_n_240__18_;
      r_240__17_ <= r_n_240__17_;
      r_240__16_ <= r_n_240__16_;
      r_240__15_ <= r_n_240__15_;
      r_240__14_ <= r_n_240__14_;
      r_240__13_ <= r_n_240__13_;
      r_240__12_ <= r_n_240__12_;
      r_240__11_ <= r_n_240__11_;
      r_240__10_ <= r_n_240__10_;
      r_240__9_ <= r_n_240__9_;
      r_240__8_ <= r_n_240__8_;
      r_240__7_ <= r_n_240__7_;
      r_240__6_ <= r_n_240__6_;
      r_240__5_ <= r_n_240__5_;
      r_240__4_ <= r_n_240__4_;
      r_240__3_ <= r_n_240__3_;
      r_240__2_ <= r_n_240__2_;
      r_240__1_ <= r_n_240__1_;
      r_240__0_ <= r_n_240__0_;
    end 
    if(N3825) begin
      r_241__63_ <= r_n_241__63_;
      r_241__62_ <= r_n_241__62_;
      r_241__61_ <= r_n_241__61_;
      r_241__60_ <= r_n_241__60_;
      r_241__59_ <= r_n_241__59_;
      r_241__58_ <= r_n_241__58_;
      r_241__57_ <= r_n_241__57_;
      r_241__56_ <= r_n_241__56_;
      r_241__55_ <= r_n_241__55_;
      r_241__54_ <= r_n_241__54_;
      r_241__53_ <= r_n_241__53_;
      r_241__52_ <= r_n_241__52_;
      r_241__51_ <= r_n_241__51_;
      r_241__50_ <= r_n_241__50_;
      r_241__49_ <= r_n_241__49_;
      r_241__48_ <= r_n_241__48_;
      r_241__47_ <= r_n_241__47_;
      r_241__46_ <= r_n_241__46_;
      r_241__45_ <= r_n_241__45_;
      r_241__44_ <= r_n_241__44_;
      r_241__43_ <= r_n_241__43_;
      r_241__42_ <= r_n_241__42_;
      r_241__41_ <= r_n_241__41_;
      r_241__40_ <= r_n_241__40_;
      r_241__39_ <= r_n_241__39_;
      r_241__38_ <= r_n_241__38_;
      r_241__37_ <= r_n_241__37_;
      r_241__36_ <= r_n_241__36_;
      r_241__35_ <= r_n_241__35_;
      r_241__34_ <= r_n_241__34_;
      r_241__33_ <= r_n_241__33_;
      r_241__32_ <= r_n_241__32_;
      r_241__31_ <= r_n_241__31_;
      r_241__30_ <= r_n_241__30_;
      r_241__29_ <= r_n_241__29_;
      r_241__28_ <= r_n_241__28_;
      r_241__27_ <= r_n_241__27_;
      r_241__26_ <= r_n_241__26_;
      r_241__25_ <= r_n_241__25_;
      r_241__24_ <= r_n_241__24_;
      r_241__23_ <= r_n_241__23_;
      r_241__22_ <= r_n_241__22_;
      r_241__21_ <= r_n_241__21_;
      r_241__20_ <= r_n_241__20_;
      r_241__19_ <= r_n_241__19_;
      r_241__18_ <= r_n_241__18_;
      r_241__17_ <= r_n_241__17_;
      r_241__16_ <= r_n_241__16_;
      r_241__15_ <= r_n_241__15_;
      r_241__14_ <= r_n_241__14_;
      r_241__13_ <= r_n_241__13_;
      r_241__12_ <= r_n_241__12_;
      r_241__11_ <= r_n_241__11_;
      r_241__10_ <= r_n_241__10_;
      r_241__9_ <= r_n_241__9_;
      r_241__8_ <= r_n_241__8_;
      r_241__7_ <= r_n_241__7_;
      r_241__6_ <= r_n_241__6_;
      r_241__5_ <= r_n_241__5_;
      r_241__4_ <= r_n_241__4_;
      r_241__3_ <= r_n_241__3_;
      r_241__2_ <= r_n_241__2_;
      r_241__1_ <= r_n_241__1_;
      r_241__0_ <= r_n_241__0_;
    end 
    if(N3826) begin
      r_242__63_ <= r_n_242__63_;
      r_242__62_ <= r_n_242__62_;
      r_242__61_ <= r_n_242__61_;
      r_242__60_ <= r_n_242__60_;
      r_242__59_ <= r_n_242__59_;
      r_242__58_ <= r_n_242__58_;
      r_242__57_ <= r_n_242__57_;
      r_242__56_ <= r_n_242__56_;
      r_242__55_ <= r_n_242__55_;
      r_242__54_ <= r_n_242__54_;
      r_242__53_ <= r_n_242__53_;
      r_242__52_ <= r_n_242__52_;
      r_242__51_ <= r_n_242__51_;
      r_242__50_ <= r_n_242__50_;
      r_242__49_ <= r_n_242__49_;
      r_242__48_ <= r_n_242__48_;
      r_242__47_ <= r_n_242__47_;
      r_242__46_ <= r_n_242__46_;
      r_242__45_ <= r_n_242__45_;
      r_242__44_ <= r_n_242__44_;
      r_242__43_ <= r_n_242__43_;
      r_242__42_ <= r_n_242__42_;
      r_242__41_ <= r_n_242__41_;
      r_242__40_ <= r_n_242__40_;
      r_242__39_ <= r_n_242__39_;
      r_242__38_ <= r_n_242__38_;
      r_242__37_ <= r_n_242__37_;
      r_242__36_ <= r_n_242__36_;
      r_242__35_ <= r_n_242__35_;
      r_242__34_ <= r_n_242__34_;
      r_242__33_ <= r_n_242__33_;
      r_242__32_ <= r_n_242__32_;
      r_242__31_ <= r_n_242__31_;
      r_242__30_ <= r_n_242__30_;
      r_242__29_ <= r_n_242__29_;
      r_242__28_ <= r_n_242__28_;
      r_242__27_ <= r_n_242__27_;
      r_242__26_ <= r_n_242__26_;
      r_242__25_ <= r_n_242__25_;
      r_242__24_ <= r_n_242__24_;
      r_242__23_ <= r_n_242__23_;
      r_242__22_ <= r_n_242__22_;
      r_242__21_ <= r_n_242__21_;
      r_242__20_ <= r_n_242__20_;
      r_242__19_ <= r_n_242__19_;
      r_242__18_ <= r_n_242__18_;
      r_242__17_ <= r_n_242__17_;
      r_242__16_ <= r_n_242__16_;
      r_242__15_ <= r_n_242__15_;
      r_242__14_ <= r_n_242__14_;
      r_242__13_ <= r_n_242__13_;
      r_242__12_ <= r_n_242__12_;
      r_242__11_ <= r_n_242__11_;
      r_242__10_ <= r_n_242__10_;
      r_242__9_ <= r_n_242__9_;
      r_242__8_ <= r_n_242__8_;
      r_242__7_ <= r_n_242__7_;
      r_242__6_ <= r_n_242__6_;
      r_242__5_ <= r_n_242__5_;
      r_242__4_ <= r_n_242__4_;
      r_242__3_ <= r_n_242__3_;
      r_242__2_ <= r_n_242__2_;
      r_242__1_ <= r_n_242__1_;
      r_242__0_ <= r_n_242__0_;
    end 
    if(N3827) begin
      r_243__63_ <= r_n_243__63_;
      r_243__62_ <= r_n_243__62_;
      r_243__61_ <= r_n_243__61_;
      r_243__60_ <= r_n_243__60_;
      r_243__59_ <= r_n_243__59_;
      r_243__58_ <= r_n_243__58_;
      r_243__57_ <= r_n_243__57_;
      r_243__56_ <= r_n_243__56_;
      r_243__55_ <= r_n_243__55_;
      r_243__54_ <= r_n_243__54_;
      r_243__53_ <= r_n_243__53_;
      r_243__52_ <= r_n_243__52_;
      r_243__51_ <= r_n_243__51_;
      r_243__50_ <= r_n_243__50_;
      r_243__49_ <= r_n_243__49_;
      r_243__48_ <= r_n_243__48_;
      r_243__47_ <= r_n_243__47_;
      r_243__46_ <= r_n_243__46_;
      r_243__45_ <= r_n_243__45_;
      r_243__44_ <= r_n_243__44_;
      r_243__43_ <= r_n_243__43_;
      r_243__42_ <= r_n_243__42_;
      r_243__41_ <= r_n_243__41_;
      r_243__40_ <= r_n_243__40_;
      r_243__39_ <= r_n_243__39_;
      r_243__38_ <= r_n_243__38_;
      r_243__37_ <= r_n_243__37_;
      r_243__36_ <= r_n_243__36_;
      r_243__35_ <= r_n_243__35_;
      r_243__34_ <= r_n_243__34_;
      r_243__33_ <= r_n_243__33_;
      r_243__32_ <= r_n_243__32_;
      r_243__31_ <= r_n_243__31_;
      r_243__30_ <= r_n_243__30_;
      r_243__29_ <= r_n_243__29_;
      r_243__28_ <= r_n_243__28_;
      r_243__27_ <= r_n_243__27_;
      r_243__26_ <= r_n_243__26_;
      r_243__25_ <= r_n_243__25_;
      r_243__24_ <= r_n_243__24_;
      r_243__23_ <= r_n_243__23_;
      r_243__22_ <= r_n_243__22_;
      r_243__21_ <= r_n_243__21_;
      r_243__20_ <= r_n_243__20_;
      r_243__19_ <= r_n_243__19_;
      r_243__18_ <= r_n_243__18_;
      r_243__17_ <= r_n_243__17_;
      r_243__16_ <= r_n_243__16_;
      r_243__15_ <= r_n_243__15_;
      r_243__14_ <= r_n_243__14_;
      r_243__13_ <= r_n_243__13_;
      r_243__12_ <= r_n_243__12_;
      r_243__11_ <= r_n_243__11_;
      r_243__10_ <= r_n_243__10_;
      r_243__9_ <= r_n_243__9_;
      r_243__8_ <= r_n_243__8_;
      r_243__7_ <= r_n_243__7_;
      r_243__6_ <= r_n_243__6_;
      r_243__5_ <= r_n_243__5_;
      r_243__4_ <= r_n_243__4_;
      r_243__3_ <= r_n_243__3_;
      r_243__2_ <= r_n_243__2_;
      r_243__1_ <= r_n_243__1_;
      r_243__0_ <= r_n_243__0_;
    end 
    if(N3828) begin
      r_244__63_ <= r_n_244__63_;
      r_244__62_ <= r_n_244__62_;
      r_244__61_ <= r_n_244__61_;
      r_244__60_ <= r_n_244__60_;
      r_244__59_ <= r_n_244__59_;
      r_244__58_ <= r_n_244__58_;
      r_244__57_ <= r_n_244__57_;
      r_244__56_ <= r_n_244__56_;
      r_244__55_ <= r_n_244__55_;
      r_244__54_ <= r_n_244__54_;
      r_244__53_ <= r_n_244__53_;
      r_244__52_ <= r_n_244__52_;
      r_244__51_ <= r_n_244__51_;
      r_244__50_ <= r_n_244__50_;
      r_244__49_ <= r_n_244__49_;
      r_244__48_ <= r_n_244__48_;
      r_244__47_ <= r_n_244__47_;
      r_244__46_ <= r_n_244__46_;
      r_244__45_ <= r_n_244__45_;
      r_244__44_ <= r_n_244__44_;
      r_244__43_ <= r_n_244__43_;
      r_244__42_ <= r_n_244__42_;
      r_244__41_ <= r_n_244__41_;
      r_244__40_ <= r_n_244__40_;
      r_244__39_ <= r_n_244__39_;
      r_244__38_ <= r_n_244__38_;
      r_244__37_ <= r_n_244__37_;
      r_244__36_ <= r_n_244__36_;
      r_244__35_ <= r_n_244__35_;
      r_244__34_ <= r_n_244__34_;
      r_244__33_ <= r_n_244__33_;
      r_244__32_ <= r_n_244__32_;
      r_244__31_ <= r_n_244__31_;
      r_244__30_ <= r_n_244__30_;
      r_244__29_ <= r_n_244__29_;
      r_244__28_ <= r_n_244__28_;
      r_244__27_ <= r_n_244__27_;
      r_244__26_ <= r_n_244__26_;
      r_244__25_ <= r_n_244__25_;
      r_244__24_ <= r_n_244__24_;
      r_244__23_ <= r_n_244__23_;
      r_244__22_ <= r_n_244__22_;
      r_244__21_ <= r_n_244__21_;
      r_244__20_ <= r_n_244__20_;
      r_244__19_ <= r_n_244__19_;
      r_244__18_ <= r_n_244__18_;
      r_244__17_ <= r_n_244__17_;
      r_244__16_ <= r_n_244__16_;
      r_244__15_ <= r_n_244__15_;
      r_244__14_ <= r_n_244__14_;
      r_244__13_ <= r_n_244__13_;
      r_244__12_ <= r_n_244__12_;
      r_244__11_ <= r_n_244__11_;
      r_244__10_ <= r_n_244__10_;
      r_244__9_ <= r_n_244__9_;
      r_244__8_ <= r_n_244__8_;
      r_244__7_ <= r_n_244__7_;
      r_244__6_ <= r_n_244__6_;
      r_244__5_ <= r_n_244__5_;
      r_244__4_ <= r_n_244__4_;
      r_244__3_ <= r_n_244__3_;
      r_244__2_ <= r_n_244__2_;
      r_244__1_ <= r_n_244__1_;
      r_244__0_ <= r_n_244__0_;
    end 
    if(N3829) begin
      r_245__63_ <= r_n_245__63_;
      r_245__62_ <= r_n_245__62_;
      r_245__61_ <= r_n_245__61_;
      r_245__60_ <= r_n_245__60_;
      r_245__59_ <= r_n_245__59_;
      r_245__58_ <= r_n_245__58_;
      r_245__57_ <= r_n_245__57_;
      r_245__56_ <= r_n_245__56_;
      r_245__55_ <= r_n_245__55_;
      r_245__54_ <= r_n_245__54_;
      r_245__53_ <= r_n_245__53_;
      r_245__52_ <= r_n_245__52_;
      r_245__51_ <= r_n_245__51_;
      r_245__50_ <= r_n_245__50_;
      r_245__49_ <= r_n_245__49_;
      r_245__48_ <= r_n_245__48_;
      r_245__47_ <= r_n_245__47_;
      r_245__46_ <= r_n_245__46_;
      r_245__45_ <= r_n_245__45_;
      r_245__44_ <= r_n_245__44_;
      r_245__43_ <= r_n_245__43_;
      r_245__42_ <= r_n_245__42_;
      r_245__41_ <= r_n_245__41_;
      r_245__40_ <= r_n_245__40_;
      r_245__39_ <= r_n_245__39_;
      r_245__38_ <= r_n_245__38_;
      r_245__37_ <= r_n_245__37_;
      r_245__36_ <= r_n_245__36_;
      r_245__35_ <= r_n_245__35_;
      r_245__34_ <= r_n_245__34_;
      r_245__33_ <= r_n_245__33_;
      r_245__32_ <= r_n_245__32_;
      r_245__31_ <= r_n_245__31_;
      r_245__30_ <= r_n_245__30_;
      r_245__29_ <= r_n_245__29_;
      r_245__28_ <= r_n_245__28_;
      r_245__27_ <= r_n_245__27_;
      r_245__26_ <= r_n_245__26_;
      r_245__25_ <= r_n_245__25_;
      r_245__24_ <= r_n_245__24_;
      r_245__23_ <= r_n_245__23_;
      r_245__22_ <= r_n_245__22_;
      r_245__21_ <= r_n_245__21_;
      r_245__20_ <= r_n_245__20_;
      r_245__19_ <= r_n_245__19_;
      r_245__18_ <= r_n_245__18_;
      r_245__17_ <= r_n_245__17_;
      r_245__16_ <= r_n_245__16_;
      r_245__15_ <= r_n_245__15_;
      r_245__14_ <= r_n_245__14_;
      r_245__13_ <= r_n_245__13_;
      r_245__12_ <= r_n_245__12_;
      r_245__11_ <= r_n_245__11_;
      r_245__10_ <= r_n_245__10_;
      r_245__9_ <= r_n_245__9_;
      r_245__8_ <= r_n_245__8_;
      r_245__7_ <= r_n_245__7_;
      r_245__6_ <= r_n_245__6_;
      r_245__5_ <= r_n_245__5_;
      r_245__4_ <= r_n_245__4_;
      r_245__3_ <= r_n_245__3_;
      r_245__2_ <= r_n_245__2_;
      r_245__1_ <= r_n_245__1_;
      r_245__0_ <= r_n_245__0_;
    end 
    if(N3830) begin
      r_246__63_ <= r_n_246__63_;
      r_246__62_ <= r_n_246__62_;
      r_246__61_ <= r_n_246__61_;
      r_246__60_ <= r_n_246__60_;
      r_246__59_ <= r_n_246__59_;
      r_246__58_ <= r_n_246__58_;
      r_246__57_ <= r_n_246__57_;
      r_246__56_ <= r_n_246__56_;
      r_246__55_ <= r_n_246__55_;
      r_246__54_ <= r_n_246__54_;
      r_246__53_ <= r_n_246__53_;
      r_246__52_ <= r_n_246__52_;
      r_246__51_ <= r_n_246__51_;
      r_246__50_ <= r_n_246__50_;
      r_246__49_ <= r_n_246__49_;
      r_246__48_ <= r_n_246__48_;
      r_246__47_ <= r_n_246__47_;
      r_246__46_ <= r_n_246__46_;
      r_246__45_ <= r_n_246__45_;
      r_246__44_ <= r_n_246__44_;
      r_246__43_ <= r_n_246__43_;
      r_246__42_ <= r_n_246__42_;
      r_246__41_ <= r_n_246__41_;
      r_246__40_ <= r_n_246__40_;
      r_246__39_ <= r_n_246__39_;
      r_246__38_ <= r_n_246__38_;
      r_246__37_ <= r_n_246__37_;
      r_246__36_ <= r_n_246__36_;
      r_246__35_ <= r_n_246__35_;
      r_246__34_ <= r_n_246__34_;
      r_246__33_ <= r_n_246__33_;
      r_246__32_ <= r_n_246__32_;
      r_246__31_ <= r_n_246__31_;
      r_246__30_ <= r_n_246__30_;
      r_246__29_ <= r_n_246__29_;
      r_246__28_ <= r_n_246__28_;
      r_246__27_ <= r_n_246__27_;
      r_246__26_ <= r_n_246__26_;
      r_246__25_ <= r_n_246__25_;
      r_246__24_ <= r_n_246__24_;
      r_246__23_ <= r_n_246__23_;
      r_246__22_ <= r_n_246__22_;
      r_246__21_ <= r_n_246__21_;
      r_246__20_ <= r_n_246__20_;
      r_246__19_ <= r_n_246__19_;
      r_246__18_ <= r_n_246__18_;
      r_246__17_ <= r_n_246__17_;
      r_246__16_ <= r_n_246__16_;
      r_246__15_ <= r_n_246__15_;
      r_246__14_ <= r_n_246__14_;
      r_246__13_ <= r_n_246__13_;
      r_246__12_ <= r_n_246__12_;
      r_246__11_ <= r_n_246__11_;
      r_246__10_ <= r_n_246__10_;
      r_246__9_ <= r_n_246__9_;
      r_246__8_ <= r_n_246__8_;
      r_246__7_ <= r_n_246__7_;
      r_246__6_ <= r_n_246__6_;
      r_246__5_ <= r_n_246__5_;
      r_246__4_ <= r_n_246__4_;
      r_246__3_ <= r_n_246__3_;
      r_246__2_ <= r_n_246__2_;
      r_246__1_ <= r_n_246__1_;
      r_246__0_ <= r_n_246__0_;
    end 
    if(N3831) begin
      r_247__63_ <= r_n_247__63_;
      r_247__62_ <= r_n_247__62_;
      r_247__61_ <= r_n_247__61_;
      r_247__60_ <= r_n_247__60_;
      r_247__59_ <= r_n_247__59_;
      r_247__58_ <= r_n_247__58_;
      r_247__57_ <= r_n_247__57_;
      r_247__56_ <= r_n_247__56_;
      r_247__55_ <= r_n_247__55_;
      r_247__54_ <= r_n_247__54_;
      r_247__53_ <= r_n_247__53_;
      r_247__52_ <= r_n_247__52_;
      r_247__51_ <= r_n_247__51_;
      r_247__50_ <= r_n_247__50_;
      r_247__49_ <= r_n_247__49_;
      r_247__48_ <= r_n_247__48_;
      r_247__47_ <= r_n_247__47_;
      r_247__46_ <= r_n_247__46_;
      r_247__45_ <= r_n_247__45_;
      r_247__44_ <= r_n_247__44_;
      r_247__43_ <= r_n_247__43_;
      r_247__42_ <= r_n_247__42_;
      r_247__41_ <= r_n_247__41_;
      r_247__40_ <= r_n_247__40_;
      r_247__39_ <= r_n_247__39_;
      r_247__38_ <= r_n_247__38_;
      r_247__37_ <= r_n_247__37_;
      r_247__36_ <= r_n_247__36_;
      r_247__35_ <= r_n_247__35_;
      r_247__34_ <= r_n_247__34_;
      r_247__33_ <= r_n_247__33_;
      r_247__32_ <= r_n_247__32_;
      r_247__31_ <= r_n_247__31_;
      r_247__30_ <= r_n_247__30_;
      r_247__29_ <= r_n_247__29_;
      r_247__28_ <= r_n_247__28_;
      r_247__27_ <= r_n_247__27_;
      r_247__26_ <= r_n_247__26_;
      r_247__25_ <= r_n_247__25_;
      r_247__24_ <= r_n_247__24_;
      r_247__23_ <= r_n_247__23_;
      r_247__22_ <= r_n_247__22_;
      r_247__21_ <= r_n_247__21_;
      r_247__20_ <= r_n_247__20_;
      r_247__19_ <= r_n_247__19_;
      r_247__18_ <= r_n_247__18_;
      r_247__17_ <= r_n_247__17_;
      r_247__16_ <= r_n_247__16_;
      r_247__15_ <= r_n_247__15_;
      r_247__14_ <= r_n_247__14_;
      r_247__13_ <= r_n_247__13_;
      r_247__12_ <= r_n_247__12_;
      r_247__11_ <= r_n_247__11_;
      r_247__10_ <= r_n_247__10_;
      r_247__9_ <= r_n_247__9_;
      r_247__8_ <= r_n_247__8_;
      r_247__7_ <= r_n_247__7_;
      r_247__6_ <= r_n_247__6_;
      r_247__5_ <= r_n_247__5_;
      r_247__4_ <= r_n_247__4_;
      r_247__3_ <= r_n_247__3_;
      r_247__2_ <= r_n_247__2_;
      r_247__1_ <= r_n_247__1_;
      r_247__0_ <= r_n_247__0_;
    end 
    if(N3832) begin
      r_248__63_ <= r_n_248__63_;
      r_248__62_ <= r_n_248__62_;
      r_248__61_ <= r_n_248__61_;
      r_248__60_ <= r_n_248__60_;
      r_248__59_ <= r_n_248__59_;
      r_248__58_ <= r_n_248__58_;
      r_248__57_ <= r_n_248__57_;
      r_248__56_ <= r_n_248__56_;
      r_248__55_ <= r_n_248__55_;
      r_248__54_ <= r_n_248__54_;
      r_248__53_ <= r_n_248__53_;
      r_248__52_ <= r_n_248__52_;
      r_248__51_ <= r_n_248__51_;
      r_248__50_ <= r_n_248__50_;
      r_248__49_ <= r_n_248__49_;
      r_248__48_ <= r_n_248__48_;
      r_248__47_ <= r_n_248__47_;
      r_248__46_ <= r_n_248__46_;
      r_248__45_ <= r_n_248__45_;
      r_248__44_ <= r_n_248__44_;
      r_248__43_ <= r_n_248__43_;
      r_248__42_ <= r_n_248__42_;
      r_248__41_ <= r_n_248__41_;
      r_248__40_ <= r_n_248__40_;
      r_248__39_ <= r_n_248__39_;
      r_248__38_ <= r_n_248__38_;
      r_248__37_ <= r_n_248__37_;
      r_248__36_ <= r_n_248__36_;
      r_248__35_ <= r_n_248__35_;
      r_248__34_ <= r_n_248__34_;
      r_248__33_ <= r_n_248__33_;
      r_248__32_ <= r_n_248__32_;
      r_248__31_ <= r_n_248__31_;
      r_248__30_ <= r_n_248__30_;
      r_248__29_ <= r_n_248__29_;
      r_248__28_ <= r_n_248__28_;
      r_248__27_ <= r_n_248__27_;
      r_248__26_ <= r_n_248__26_;
      r_248__25_ <= r_n_248__25_;
      r_248__24_ <= r_n_248__24_;
      r_248__23_ <= r_n_248__23_;
      r_248__22_ <= r_n_248__22_;
      r_248__21_ <= r_n_248__21_;
      r_248__20_ <= r_n_248__20_;
      r_248__19_ <= r_n_248__19_;
      r_248__18_ <= r_n_248__18_;
      r_248__17_ <= r_n_248__17_;
      r_248__16_ <= r_n_248__16_;
      r_248__15_ <= r_n_248__15_;
      r_248__14_ <= r_n_248__14_;
      r_248__13_ <= r_n_248__13_;
      r_248__12_ <= r_n_248__12_;
      r_248__11_ <= r_n_248__11_;
      r_248__10_ <= r_n_248__10_;
      r_248__9_ <= r_n_248__9_;
      r_248__8_ <= r_n_248__8_;
      r_248__7_ <= r_n_248__7_;
      r_248__6_ <= r_n_248__6_;
      r_248__5_ <= r_n_248__5_;
      r_248__4_ <= r_n_248__4_;
      r_248__3_ <= r_n_248__3_;
      r_248__2_ <= r_n_248__2_;
      r_248__1_ <= r_n_248__1_;
      r_248__0_ <= r_n_248__0_;
    end 
    if(N3833) begin
      r_249__63_ <= r_n_249__63_;
      r_249__62_ <= r_n_249__62_;
      r_249__61_ <= r_n_249__61_;
      r_249__60_ <= r_n_249__60_;
      r_249__59_ <= r_n_249__59_;
      r_249__58_ <= r_n_249__58_;
      r_249__57_ <= r_n_249__57_;
      r_249__56_ <= r_n_249__56_;
      r_249__55_ <= r_n_249__55_;
      r_249__54_ <= r_n_249__54_;
      r_249__53_ <= r_n_249__53_;
      r_249__52_ <= r_n_249__52_;
      r_249__51_ <= r_n_249__51_;
      r_249__50_ <= r_n_249__50_;
      r_249__49_ <= r_n_249__49_;
      r_249__48_ <= r_n_249__48_;
      r_249__47_ <= r_n_249__47_;
      r_249__46_ <= r_n_249__46_;
      r_249__45_ <= r_n_249__45_;
      r_249__44_ <= r_n_249__44_;
      r_249__43_ <= r_n_249__43_;
      r_249__42_ <= r_n_249__42_;
      r_249__41_ <= r_n_249__41_;
      r_249__40_ <= r_n_249__40_;
      r_249__39_ <= r_n_249__39_;
      r_249__38_ <= r_n_249__38_;
      r_249__37_ <= r_n_249__37_;
      r_249__36_ <= r_n_249__36_;
      r_249__35_ <= r_n_249__35_;
      r_249__34_ <= r_n_249__34_;
      r_249__33_ <= r_n_249__33_;
      r_249__32_ <= r_n_249__32_;
      r_249__31_ <= r_n_249__31_;
      r_249__30_ <= r_n_249__30_;
      r_249__29_ <= r_n_249__29_;
      r_249__28_ <= r_n_249__28_;
      r_249__27_ <= r_n_249__27_;
      r_249__26_ <= r_n_249__26_;
      r_249__25_ <= r_n_249__25_;
      r_249__24_ <= r_n_249__24_;
      r_249__23_ <= r_n_249__23_;
      r_249__22_ <= r_n_249__22_;
      r_249__21_ <= r_n_249__21_;
      r_249__20_ <= r_n_249__20_;
      r_249__19_ <= r_n_249__19_;
      r_249__18_ <= r_n_249__18_;
      r_249__17_ <= r_n_249__17_;
      r_249__16_ <= r_n_249__16_;
      r_249__15_ <= r_n_249__15_;
      r_249__14_ <= r_n_249__14_;
      r_249__13_ <= r_n_249__13_;
      r_249__12_ <= r_n_249__12_;
      r_249__11_ <= r_n_249__11_;
      r_249__10_ <= r_n_249__10_;
      r_249__9_ <= r_n_249__9_;
      r_249__8_ <= r_n_249__8_;
      r_249__7_ <= r_n_249__7_;
      r_249__6_ <= r_n_249__6_;
      r_249__5_ <= r_n_249__5_;
      r_249__4_ <= r_n_249__4_;
      r_249__3_ <= r_n_249__3_;
      r_249__2_ <= r_n_249__2_;
      r_249__1_ <= r_n_249__1_;
      r_249__0_ <= r_n_249__0_;
    end 
    if(N3834) begin
      r_250__63_ <= r_n_250__63_;
      r_250__62_ <= r_n_250__62_;
      r_250__61_ <= r_n_250__61_;
      r_250__60_ <= r_n_250__60_;
      r_250__59_ <= r_n_250__59_;
      r_250__58_ <= r_n_250__58_;
      r_250__57_ <= r_n_250__57_;
      r_250__56_ <= r_n_250__56_;
      r_250__55_ <= r_n_250__55_;
      r_250__54_ <= r_n_250__54_;
      r_250__53_ <= r_n_250__53_;
      r_250__52_ <= r_n_250__52_;
      r_250__51_ <= r_n_250__51_;
      r_250__50_ <= r_n_250__50_;
      r_250__49_ <= r_n_250__49_;
      r_250__48_ <= r_n_250__48_;
      r_250__47_ <= r_n_250__47_;
      r_250__46_ <= r_n_250__46_;
      r_250__45_ <= r_n_250__45_;
      r_250__44_ <= r_n_250__44_;
      r_250__43_ <= r_n_250__43_;
      r_250__42_ <= r_n_250__42_;
      r_250__41_ <= r_n_250__41_;
      r_250__40_ <= r_n_250__40_;
      r_250__39_ <= r_n_250__39_;
      r_250__38_ <= r_n_250__38_;
      r_250__37_ <= r_n_250__37_;
      r_250__36_ <= r_n_250__36_;
      r_250__35_ <= r_n_250__35_;
      r_250__34_ <= r_n_250__34_;
      r_250__33_ <= r_n_250__33_;
      r_250__32_ <= r_n_250__32_;
      r_250__31_ <= r_n_250__31_;
      r_250__30_ <= r_n_250__30_;
      r_250__29_ <= r_n_250__29_;
      r_250__28_ <= r_n_250__28_;
      r_250__27_ <= r_n_250__27_;
      r_250__26_ <= r_n_250__26_;
      r_250__25_ <= r_n_250__25_;
      r_250__24_ <= r_n_250__24_;
      r_250__23_ <= r_n_250__23_;
      r_250__22_ <= r_n_250__22_;
      r_250__21_ <= r_n_250__21_;
      r_250__20_ <= r_n_250__20_;
      r_250__19_ <= r_n_250__19_;
      r_250__18_ <= r_n_250__18_;
      r_250__17_ <= r_n_250__17_;
      r_250__16_ <= r_n_250__16_;
      r_250__15_ <= r_n_250__15_;
      r_250__14_ <= r_n_250__14_;
      r_250__13_ <= r_n_250__13_;
      r_250__12_ <= r_n_250__12_;
      r_250__11_ <= r_n_250__11_;
      r_250__10_ <= r_n_250__10_;
      r_250__9_ <= r_n_250__9_;
      r_250__8_ <= r_n_250__8_;
      r_250__7_ <= r_n_250__7_;
      r_250__6_ <= r_n_250__6_;
      r_250__5_ <= r_n_250__5_;
      r_250__4_ <= r_n_250__4_;
      r_250__3_ <= r_n_250__3_;
      r_250__2_ <= r_n_250__2_;
      r_250__1_ <= r_n_250__1_;
      r_250__0_ <= r_n_250__0_;
    end 
    if(N3835) begin
      r_251__63_ <= r_n_251__63_;
      r_251__62_ <= r_n_251__62_;
      r_251__61_ <= r_n_251__61_;
      r_251__60_ <= r_n_251__60_;
      r_251__59_ <= r_n_251__59_;
      r_251__58_ <= r_n_251__58_;
      r_251__57_ <= r_n_251__57_;
      r_251__56_ <= r_n_251__56_;
      r_251__55_ <= r_n_251__55_;
      r_251__54_ <= r_n_251__54_;
      r_251__53_ <= r_n_251__53_;
      r_251__52_ <= r_n_251__52_;
      r_251__51_ <= r_n_251__51_;
      r_251__50_ <= r_n_251__50_;
      r_251__49_ <= r_n_251__49_;
      r_251__48_ <= r_n_251__48_;
      r_251__47_ <= r_n_251__47_;
      r_251__46_ <= r_n_251__46_;
      r_251__45_ <= r_n_251__45_;
      r_251__44_ <= r_n_251__44_;
      r_251__43_ <= r_n_251__43_;
      r_251__42_ <= r_n_251__42_;
      r_251__41_ <= r_n_251__41_;
      r_251__40_ <= r_n_251__40_;
      r_251__39_ <= r_n_251__39_;
      r_251__38_ <= r_n_251__38_;
      r_251__37_ <= r_n_251__37_;
      r_251__36_ <= r_n_251__36_;
      r_251__35_ <= r_n_251__35_;
      r_251__34_ <= r_n_251__34_;
      r_251__33_ <= r_n_251__33_;
      r_251__32_ <= r_n_251__32_;
      r_251__31_ <= r_n_251__31_;
      r_251__30_ <= r_n_251__30_;
      r_251__29_ <= r_n_251__29_;
      r_251__28_ <= r_n_251__28_;
      r_251__27_ <= r_n_251__27_;
      r_251__26_ <= r_n_251__26_;
      r_251__25_ <= r_n_251__25_;
      r_251__24_ <= r_n_251__24_;
      r_251__23_ <= r_n_251__23_;
      r_251__22_ <= r_n_251__22_;
      r_251__21_ <= r_n_251__21_;
      r_251__20_ <= r_n_251__20_;
      r_251__19_ <= r_n_251__19_;
      r_251__18_ <= r_n_251__18_;
      r_251__17_ <= r_n_251__17_;
      r_251__16_ <= r_n_251__16_;
      r_251__15_ <= r_n_251__15_;
      r_251__14_ <= r_n_251__14_;
      r_251__13_ <= r_n_251__13_;
      r_251__12_ <= r_n_251__12_;
      r_251__11_ <= r_n_251__11_;
      r_251__10_ <= r_n_251__10_;
      r_251__9_ <= r_n_251__9_;
      r_251__8_ <= r_n_251__8_;
      r_251__7_ <= r_n_251__7_;
      r_251__6_ <= r_n_251__6_;
      r_251__5_ <= r_n_251__5_;
      r_251__4_ <= r_n_251__4_;
      r_251__3_ <= r_n_251__3_;
      r_251__2_ <= r_n_251__2_;
      r_251__1_ <= r_n_251__1_;
      r_251__0_ <= r_n_251__0_;
    end 
    if(N3836) begin
      r_252__63_ <= r_n_252__63_;
      r_252__62_ <= r_n_252__62_;
      r_252__61_ <= r_n_252__61_;
      r_252__60_ <= r_n_252__60_;
      r_252__59_ <= r_n_252__59_;
      r_252__58_ <= r_n_252__58_;
      r_252__57_ <= r_n_252__57_;
      r_252__56_ <= r_n_252__56_;
      r_252__55_ <= r_n_252__55_;
      r_252__54_ <= r_n_252__54_;
      r_252__53_ <= r_n_252__53_;
      r_252__52_ <= r_n_252__52_;
      r_252__51_ <= r_n_252__51_;
      r_252__50_ <= r_n_252__50_;
      r_252__49_ <= r_n_252__49_;
      r_252__48_ <= r_n_252__48_;
      r_252__47_ <= r_n_252__47_;
      r_252__46_ <= r_n_252__46_;
      r_252__45_ <= r_n_252__45_;
      r_252__44_ <= r_n_252__44_;
      r_252__43_ <= r_n_252__43_;
      r_252__42_ <= r_n_252__42_;
      r_252__41_ <= r_n_252__41_;
      r_252__40_ <= r_n_252__40_;
      r_252__39_ <= r_n_252__39_;
      r_252__38_ <= r_n_252__38_;
      r_252__37_ <= r_n_252__37_;
      r_252__36_ <= r_n_252__36_;
      r_252__35_ <= r_n_252__35_;
      r_252__34_ <= r_n_252__34_;
      r_252__33_ <= r_n_252__33_;
      r_252__32_ <= r_n_252__32_;
      r_252__31_ <= r_n_252__31_;
      r_252__30_ <= r_n_252__30_;
      r_252__29_ <= r_n_252__29_;
      r_252__28_ <= r_n_252__28_;
      r_252__27_ <= r_n_252__27_;
      r_252__26_ <= r_n_252__26_;
      r_252__25_ <= r_n_252__25_;
      r_252__24_ <= r_n_252__24_;
      r_252__23_ <= r_n_252__23_;
      r_252__22_ <= r_n_252__22_;
      r_252__21_ <= r_n_252__21_;
      r_252__20_ <= r_n_252__20_;
      r_252__19_ <= r_n_252__19_;
      r_252__18_ <= r_n_252__18_;
      r_252__17_ <= r_n_252__17_;
      r_252__16_ <= r_n_252__16_;
      r_252__15_ <= r_n_252__15_;
      r_252__14_ <= r_n_252__14_;
      r_252__13_ <= r_n_252__13_;
      r_252__12_ <= r_n_252__12_;
      r_252__11_ <= r_n_252__11_;
      r_252__10_ <= r_n_252__10_;
      r_252__9_ <= r_n_252__9_;
      r_252__8_ <= r_n_252__8_;
      r_252__7_ <= r_n_252__7_;
      r_252__6_ <= r_n_252__6_;
      r_252__5_ <= r_n_252__5_;
      r_252__4_ <= r_n_252__4_;
      r_252__3_ <= r_n_252__3_;
      r_252__2_ <= r_n_252__2_;
      r_252__1_ <= r_n_252__1_;
      r_252__0_ <= r_n_252__0_;
    end 
    if(N3837) begin
      r_253__63_ <= r_n_253__63_;
      r_253__62_ <= r_n_253__62_;
      r_253__61_ <= r_n_253__61_;
      r_253__60_ <= r_n_253__60_;
      r_253__59_ <= r_n_253__59_;
      r_253__58_ <= r_n_253__58_;
      r_253__57_ <= r_n_253__57_;
      r_253__56_ <= r_n_253__56_;
      r_253__55_ <= r_n_253__55_;
      r_253__54_ <= r_n_253__54_;
      r_253__53_ <= r_n_253__53_;
      r_253__52_ <= r_n_253__52_;
      r_253__51_ <= r_n_253__51_;
      r_253__50_ <= r_n_253__50_;
      r_253__49_ <= r_n_253__49_;
      r_253__48_ <= r_n_253__48_;
      r_253__47_ <= r_n_253__47_;
      r_253__46_ <= r_n_253__46_;
      r_253__45_ <= r_n_253__45_;
      r_253__44_ <= r_n_253__44_;
      r_253__43_ <= r_n_253__43_;
      r_253__42_ <= r_n_253__42_;
      r_253__41_ <= r_n_253__41_;
      r_253__40_ <= r_n_253__40_;
      r_253__39_ <= r_n_253__39_;
      r_253__38_ <= r_n_253__38_;
      r_253__37_ <= r_n_253__37_;
      r_253__36_ <= r_n_253__36_;
      r_253__35_ <= r_n_253__35_;
      r_253__34_ <= r_n_253__34_;
      r_253__33_ <= r_n_253__33_;
      r_253__32_ <= r_n_253__32_;
      r_253__31_ <= r_n_253__31_;
      r_253__30_ <= r_n_253__30_;
      r_253__29_ <= r_n_253__29_;
      r_253__28_ <= r_n_253__28_;
      r_253__27_ <= r_n_253__27_;
      r_253__26_ <= r_n_253__26_;
      r_253__25_ <= r_n_253__25_;
      r_253__24_ <= r_n_253__24_;
      r_253__23_ <= r_n_253__23_;
      r_253__22_ <= r_n_253__22_;
      r_253__21_ <= r_n_253__21_;
      r_253__20_ <= r_n_253__20_;
      r_253__19_ <= r_n_253__19_;
      r_253__18_ <= r_n_253__18_;
      r_253__17_ <= r_n_253__17_;
      r_253__16_ <= r_n_253__16_;
      r_253__15_ <= r_n_253__15_;
      r_253__14_ <= r_n_253__14_;
      r_253__13_ <= r_n_253__13_;
      r_253__12_ <= r_n_253__12_;
      r_253__11_ <= r_n_253__11_;
      r_253__10_ <= r_n_253__10_;
      r_253__9_ <= r_n_253__9_;
      r_253__8_ <= r_n_253__8_;
      r_253__7_ <= r_n_253__7_;
      r_253__6_ <= r_n_253__6_;
      r_253__5_ <= r_n_253__5_;
      r_253__4_ <= r_n_253__4_;
      r_253__3_ <= r_n_253__3_;
      r_253__2_ <= r_n_253__2_;
      r_253__1_ <= r_n_253__1_;
      r_253__0_ <= r_n_253__0_;
    end 
    if(N3838) begin
      r_254__63_ <= r_n_254__63_;
      r_254__62_ <= r_n_254__62_;
      r_254__61_ <= r_n_254__61_;
      r_254__60_ <= r_n_254__60_;
      r_254__59_ <= r_n_254__59_;
      r_254__58_ <= r_n_254__58_;
      r_254__57_ <= r_n_254__57_;
      r_254__56_ <= r_n_254__56_;
      r_254__55_ <= r_n_254__55_;
      r_254__54_ <= r_n_254__54_;
      r_254__53_ <= r_n_254__53_;
      r_254__52_ <= r_n_254__52_;
      r_254__51_ <= r_n_254__51_;
      r_254__50_ <= r_n_254__50_;
      r_254__49_ <= r_n_254__49_;
      r_254__48_ <= r_n_254__48_;
      r_254__47_ <= r_n_254__47_;
      r_254__46_ <= r_n_254__46_;
      r_254__45_ <= r_n_254__45_;
      r_254__44_ <= r_n_254__44_;
      r_254__43_ <= r_n_254__43_;
      r_254__42_ <= r_n_254__42_;
      r_254__41_ <= r_n_254__41_;
      r_254__40_ <= r_n_254__40_;
      r_254__39_ <= r_n_254__39_;
      r_254__38_ <= r_n_254__38_;
      r_254__37_ <= r_n_254__37_;
      r_254__36_ <= r_n_254__36_;
      r_254__35_ <= r_n_254__35_;
      r_254__34_ <= r_n_254__34_;
      r_254__33_ <= r_n_254__33_;
      r_254__32_ <= r_n_254__32_;
      r_254__31_ <= r_n_254__31_;
      r_254__30_ <= r_n_254__30_;
      r_254__29_ <= r_n_254__29_;
      r_254__28_ <= r_n_254__28_;
      r_254__27_ <= r_n_254__27_;
      r_254__26_ <= r_n_254__26_;
      r_254__25_ <= r_n_254__25_;
      r_254__24_ <= r_n_254__24_;
      r_254__23_ <= r_n_254__23_;
      r_254__22_ <= r_n_254__22_;
      r_254__21_ <= r_n_254__21_;
      r_254__20_ <= r_n_254__20_;
      r_254__19_ <= r_n_254__19_;
      r_254__18_ <= r_n_254__18_;
      r_254__17_ <= r_n_254__17_;
      r_254__16_ <= r_n_254__16_;
      r_254__15_ <= r_n_254__15_;
      r_254__14_ <= r_n_254__14_;
      r_254__13_ <= r_n_254__13_;
      r_254__12_ <= r_n_254__12_;
      r_254__11_ <= r_n_254__11_;
      r_254__10_ <= r_n_254__10_;
      r_254__9_ <= r_n_254__9_;
      r_254__8_ <= r_n_254__8_;
      r_254__7_ <= r_n_254__7_;
      r_254__6_ <= r_n_254__6_;
      r_254__5_ <= r_n_254__5_;
      r_254__4_ <= r_n_254__4_;
      r_254__3_ <= r_n_254__3_;
      r_254__2_ <= r_n_254__2_;
      r_254__1_ <= r_n_254__1_;
      r_254__0_ <= r_n_254__0_;
    end 
    if(N3839) begin
      r_255__63_ <= r_n_255__63_;
      r_255__62_ <= r_n_255__62_;
      r_255__61_ <= r_n_255__61_;
      r_255__60_ <= r_n_255__60_;
      r_255__59_ <= r_n_255__59_;
      r_255__58_ <= r_n_255__58_;
      r_255__57_ <= r_n_255__57_;
      r_255__56_ <= r_n_255__56_;
      r_255__55_ <= r_n_255__55_;
      r_255__54_ <= r_n_255__54_;
      r_255__53_ <= r_n_255__53_;
      r_255__52_ <= r_n_255__52_;
      r_255__51_ <= r_n_255__51_;
      r_255__50_ <= r_n_255__50_;
      r_255__49_ <= r_n_255__49_;
      r_255__48_ <= r_n_255__48_;
      r_255__47_ <= r_n_255__47_;
      r_255__46_ <= r_n_255__46_;
      r_255__45_ <= r_n_255__45_;
      r_255__44_ <= r_n_255__44_;
      r_255__43_ <= r_n_255__43_;
      r_255__42_ <= r_n_255__42_;
      r_255__41_ <= r_n_255__41_;
      r_255__40_ <= r_n_255__40_;
      r_255__39_ <= r_n_255__39_;
      r_255__38_ <= r_n_255__38_;
      r_255__37_ <= r_n_255__37_;
      r_255__36_ <= r_n_255__36_;
      r_255__35_ <= r_n_255__35_;
      r_255__34_ <= r_n_255__34_;
      r_255__33_ <= r_n_255__33_;
      r_255__32_ <= r_n_255__32_;
      r_255__31_ <= r_n_255__31_;
      r_255__30_ <= r_n_255__30_;
      r_255__29_ <= r_n_255__29_;
      r_255__28_ <= r_n_255__28_;
      r_255__27_ <= r_n_255__27_;
      r_255__26_ <= r_n_255__26_;
      r_255__25_ <= r_n_255__25_;
      r_255__24_ <= r_n_255__24_;
      r_255__23_ <= r_n_255__23_;
      r_255__22_ <= r_n_255__22_;
      r_255__21_ <= r_n_255__21_;
      r_255__20_ <= r_n_255__20_;
      r_255__19_ <= r_n_255__19_;
      r_255__18_ <= r_n_255__18_;
      r_255__17_ <= r_n_255__17_;
      r_255__16_ <= r_n_255__16_;
      r_255__15_ <= r_n_255__15_;
      r_255__14_ <= r_n_255__14_;
      r_255__13_ <= r_n_255__13_;
      r_255__12_ <= r_n_255__12_;
      r_255__11_ <= r_n_255__11_;
      r_255__10_ <= r_n_255__10_;
      r_255__9_ <= r_n_255__9_;
      r_255__8_ <= r_n_255__8_;
      r_255__7_ <= r_n_255__7_;
      r_255__6_ <= r_n_255__6_;
      r_255__5_ <= r_n_255__5_;
      r_255__4_ <= r_n_255__4_;
      r_255__3_ <= r_n_255__3_;
      r_255__2_ <= r_n_255__2_;
      r_255__1_ <= r_n_255__1_;
      r_255__0_ <= r_n_255__0_;
    end 
    if(N3840) begin
      r_256__63_ <= r_n_256__63_;
      r_256__62_ <= r_n_256__62_;
      r_256__61_ <= r_n_256__61_;
      r_256__60_ <= r_n_256__60_;
      r_256__59_ <= r_n_256__59_;
      r_256__58_ <= r_n_256__58_;
      r_256__57_ <= r_n_256__57_;
      r_256__56_ <= r_n_256__56_;
      r_256__55_ <= r_n_256__55_;
      r_256__54_ <= r_n_256__54_;
      r_256__53_ <= r_n_256__53_;
      r_256__52_ <= r_n_256__52_;
      r_256__51_ <= r_n_256__51_;
      r_256__50_ <= r_n_256__50_;
      r_256__49_ <= r_n_256__49_;
      r_256__48_ <= r_n_256__48_;
      r_256__47_ <= r_n_256__47_;
      r_256__46_ <= r_n_256__46_;
      r_256__45_ <= r_n_256__45_;
      r_256__44_ <= r_n_256__44_;
      r_256__43_ <= r_n_256__43_;
      r_256__42_ <= r_n_256__42_;
      r_256__41_ <= r_n_256__41_;
      r_256__40_ <= r_n_256__40_;
      r_256__39_ <= r_n_256__39_;
      r_256__38_ <= r_n_256__38_;
      r_256__37_ <= r_n_256__37_;
      r_256__36_ <= r_n_256__36_;
      r_256__35_ <= r_n_256__35_;
      r_256__34_ <= r_n_256__34_;
      r_256__33_ <= r_n_256__33_;
      r_256__32_ <= r_n_256__32_;
      r_256__31_ <= r_n_256__31_;
      r_256__30_ <= r_n_256__30_;
      r_256__29_ <= r_n_256__29_;
      r_256__28_ <= r_n_256__28_;
      r_256__27_ <= r_n_256__27_;
      r_256__26_ <= r_n_256__26_;
      r_256__25_ <= r_n_256__25_;
      r_256__24_ <= r_n_256__24_;
      r_256__23_ <= r_n_256__23_;
      r_256__22_ <= r_n_256__22_;
      r_256__21_ <= r_n_256__21_;
      r_256__20_ <= r_n_256__20_;
      r_256__19_ <= r_n_256__19_;
      r_256__18_ <= r_n_256__18_;
      r_256__17_ <= r_n_256__17_;
      r_256__16_ <= r_n_256__16_;
      r_256__15_ <= r_n_256__15_;
      r_256__14_ <= r_n_256__14_;
      r_256__13_ <= r_n_256__13_;
      r_256__12_ <= r_n_256__12_;
      r_256__11_ <= r_n_256__11_;
      r_256__10_ <= r_n_256__10_;
      r_256__9_ <= r_n_256__9_;
      r_256__8_ <= r_n_256__8_;
      r_256__7_ <= r_n_256__7_;
      r_256__6_ <= r_n_256__6_;
      r_256__5_ <= r_n_256__5_;
      r_256__4_ <= r_n_256__4_;
      r_256__3_ <= r_n_256__3_;
      r_256__2_ <= r_n_256__2_;
      r_256__1_ <= r_n_256__1_;
      r_256__0_ <= r_n_256__0_;
    end 
    if(N3841) begin
      r_257__63_ <= r_n_257__63_;
      r_257__62_ <= r_n_257__62_;
      r_257__61_ <= r_n_257__61_;
      r_257__60_ <= r_n_257__60_;
      r_257__59_ <= r_n_257__59_;
      r_257__58_ <= r_n_257__58_;
      r_257__57_ <= r_n_257__57_;
      r_257__56_ <= r_n_257__56_;
      r_257__55_ <= r_n_257__55_;
      r_257__54_ <= r_n_257__54_;
      r_257__53_ <= r_n_257__53_;
      r_257__52_ <= r_n_257__52_;
      r_257__51_ <= r_n_257__51_;
      r_257__50_ <= r_n_257__50_;
      r_257__49_ <= r_n_257__49_;
      r_257__48_ <= r_n_257__48_;
      r_257__47_ <= r_n_257__47_;
      r_257__46_ <= r_n_257__46_;
      r_257__45_ <= r_n_257__45_;
      r_257__44_ <= r_n_257__44_;
      r_257__43_ <= r_n_257__43_;
      r_257__42_ <= r_n_257__42_;
      r_257__41_ <= r_n_257__41_;
      r_257__40_ <= r_n_257__40_;
      r_257__39_ <= r_n_257__39_;
      r_257__38_ <= r_n_257__38_;
      r_257__37_ <= r_n_257__37_;
      r_257__36_ <= r_n_257__36_;
      r_257__35_ <= r_n_257__35_;
      r_257__34_ <= r_n_257__34_;
      r_257__33_ <= r_n_257__33_;
      r_257__32_ <= r_n_257__32_;
      r_257__31_ <= r_n_257__31_;
      r_257__30_ <= r_n_257__30_;
      r_257__29_ <= r_n_257__29_;
      r_257__28_ <= r_n_257__28_;
      r_257__27_ <= r_n_257__27_;
      r_257__26_ <= r_n_257__26_;
      r_257__25_ <= r_n_257__25_;
      r_257__24_ <= r_n_257__24_;
      r_257__23_ <= r_n_257__23_;
      r_257__22_ <= r_n_257__22_;
      r_257__21_ <= r_n_257__21_;
      r_257__20_ <= r_n_257__20_;
      r_257__19_ <= r_n_257__19_;
      r_257__18_ <= r_n_257__18_;
      r_257__17_ <= r_n_257__17_;
      r_257__16_ <= r_n_257__16_;
      r_257__15_ <= r_n_257__15_;
      r_257__14_ <= r_n_257__14_;
      r_257__13_ <= r_n_257__13_;
      r_257__12_ <= r_n_257__12_;
      r_257__11_ <= r_n_257__11_;
      r_257__10_ <= r_n_257__10_;
      r_257__9_ <= r_n_257__9_;
      r_257__8_ <= r_n_257__8_;
      r_257__7_ <= r_n_257__7_;
      r_257__6_ <= r_n_257__6_;
      r_257__5_ <= r_n_257__5_;
      r_257__4_ <= r_n_257__4_;
      r_257__3_ <= r_n_257__3_;
      r_257__2_ <= r_n_257__2_;
      r_257__1_ <= r_n_257__1_;
      r_257__0_ <= r_n_257__0_;
    end 
    if(N3842) begin
      r_258__63_ <= r_n_258__63_;
      r_258__62_ <= r_n_258__62_;
      r_258__61_ <= r_n_258__61_;
      r_258__60_ <= r_n_258__60_;
      r_258__59_ <= r_n_258__59_;
      r_258__58_ <= r_n_258__58_;
      r_258__57_ <= r_n_258__57_;
      r_258__56_ <= r_n_258__56_;
      r_258__55_ <= r_n_258__55_;
      r_258__54_ <= r_n_258__54_;
      r_258__53_ <= r_n_258__53_;
      r_258__52_ <= r_n_258__52_;
      r_258__51_ <= r_n_258__51_;
      r_258__50_ <= r_n_258__50_;
      r_258__49_ <= r_n_258__49_;
      r_258__48_ <= r_n_258__48_;
      r_258__47_ <= r_n_258__47_;
      r_258__46_ <= r_n_258__46_;
      r_258__45_ <= r_n_258__45_;
      r_258__44_ <= r_n_258__44_;
      r_258__43_ <= r_n_258__43_;
      r_258__42_ <= r_n_258__42_;
      r_258__41_ <= r_n_258__41_;
      r_258__40_ <= r_n_258__40_;
      r_258__39_ <= r_n_258__39_;
      r_258__38_ <= r_n_258__38_;
      r_258__37_ <= r_n_258__37_;
      r_258__36_ <= r_n_258__36_;
      r_258__35_ <= r_n_258__35_;
      r_258__34_ <= r_n_258__34_;
      r_258__33_ <= r_n_258__33_;
      r_258__32_ <= r_n_258__32_;
      r_258__31_ <= r_n_258__31_;
      r_258__30_ <= r_n_258__30_;
      r_258__29_ <= r_n_258__29_;
      r_258__28_ <= r_n_258__28_;
      r_258__27_ <= r_n_258__27_;
      r_258__26_ <= r_n_258__26_;
      r_258__25_ <= r_n_258__25_;
      r_258__24_ <= r_n_258__24_;
      r_258__23_ <= r_n_258__23_;
      r_258__22_ <= r_n_258__22_;
      r_258__21_ <= r_n_258__21_;
      r_258__20_ <= r_n_258__20_;
      r_258__19_ <= r_n_258__19_;
      r_258__18_ <= r_n_258__18_;
      r_258__17_ <= r_n_258__17_;
      r_258__16_ <= r_n_258__16_;
      r_258__15_ <= r_n_258__15_;
      r_258__14_ <= r_n_258__14_;
      r_258__13_ <= r_n_258__13_;
      r_258__12_ <= r_n_258__12_;
      r_258__11_ <= r_n_258__11_;
      r_258__10_ <= r_n_258__10_;
      r_258__9_ <= r_n_258__9_;
      r_258__8_ <= r_n_258__8_;
      r_258__7_ <= r_n_258__7_;
      r_258__6_ <= r_n_258__6_;
      r_258__5_ <= r_n_258__5_;
      r_258__4_ <= r_n_258__4_;
      r_258__3_ <= r_n_258__3_;
      r_258__2_ <= r_n_258__2_;
      r_258__1_ <= r_n_258__1_;
      r_258__0_ <= r_n_258__0_;
    end 
    if(N3843) begin
      r_259__63_ <= r_n_259__63_;
      r_259__62_ <= r_n_259__62_;
      r_259__61_ <= r_n_259__61_;
      r_259__60_ <= r_n_259__60_;
      r_259__59_ <= r_n_259__59_;
      r_259__58_ <= r_n_259__58_;
      r_259__57_ <= r_n_259__57_;
      r_259__56_ <= r_n_259__56_;
      r_259__55_ <= r_n_259__55_;
      r_259__54_ <= r_n_259__54_;
      r_259__53_ <= r_n_259__53_;
      r_259__52_ <= r_n_259__52_;
      r_259__51_ <= r_n_259__51_;
      r_259__50_ <= r_n_259__50_;
      r_259__49_ <= r_n_259__49_;
      r_259__48_ <= r_n_259__48_;
      r_259__47_ <= r_n_259__47_;
      r_259__46_ <= r_n_259__46_;
      r_259__45_ <= r_n_259__45_;
      r_259__44_ <= r_n_259__44_;
      r_259__43_ <= r_n_259__43_;
      r_259__42_ <= r_n_259__42_;
      r_259__41_ <= r_n_259__41_;
      r_259__40_ <= r_n_259__40_;
      r_259__39_ <= r_n_259__39_;
      r_259__38_ <= r_n_259__38_;
      r_259__37_ <= r_n_259__37_;
      r_259__36_ <= r_n_259__36_;
      r_259__35_ <= r_n_259__35_;
      r_259__34_ <= r_n_259__34_;
      r_259__33_ <= r_n_259__33_;
      r_259__32_ <= r_n_259__32_;
      r_259__31_ <= r_n_259__31_;
      r_259__30_ <= r_n_259__30_;
      r_259__29_ <= r_n_259__29_;
      r_259__28_ <= r_n_259__28_;
      r_259__27_ <= r_n_259__27_;
      r_259__26_ <= r_n_259__26_;
      r_259__25_ <= r_n_259__25_;
      r_259__24_ <= r_n_259__24_;
      r_259__23_ <= r_n_259__23_;
      r_259__22_ <= r_n_259__22_;
      r_259__21_ <= r_n_259__21_;
      r_259__20_ <= r_n_259__20_;
      r_259__19_ <= r_n_259__19_;
      r_259__18_ <= r_n_259__18_;
      r_259__17_ <= r_n_259__17_;
      r_259__16_ <= r_n_259__16_;
      r_259__15_ <= r_n_259__15_;
      r_259__14_ <= r_n_259__14_;
      r_259__13_ <= r_n_259__13_;
      r_259__12_ <= r_n_259__12_;
      r_259__11_ <= r_n_259__11_;
      r_259__10_ <= r_n_259__10_;
      r_259__9_ <= r_n_259__9_;
      r_259__8_ <= r_n_259__8_;
      r_259__7_ <= r_n_259__7_;
      r_259__6_ <= r_n_259__6_;
      r_259__5_ <= r_n_259__5_;
      r_259__4_ <= r_n_259__4_;
      r_259__3_ <= r_n_259__3_;
      r_259__2_ <= r_n_259__2_;
      r_259__1_ <= r_n_259__1_;
      r_259__0_ <= r_n_259__0_;
    end 
    if(N3844) begin
      r_260__63_ <= r_n_260__63_;
      r_260__62_ <= r_n_260__62_;
      r_260__61_ <= r_n_260__61_;
      r_260__60_ <= r_n_260__60_;
      r_260__59_ <= r_n_260__59_;
      r_260__58_ <= r_n_260__58_;
      r_260__57_ <= r_n_260__57_;
      r_260__56_ <= r_n_260__56_;
      r_260__55_ <= r_n_260__55_;
      r_260__54_ <= r_n_260__54_;
      r_260__53_ <= r_n_260__53_;
      r_260__52_ <= r_n_260__52_;
      r_260__51_ <= r_n_260__51_;
      r_260__50_ <= r_n_260__50_;
      r_260__49_ <= r_n_260__49_;
      r_260__48_ <= r_n_260__48_;
      r_260__47_ <= r_n_260__47_;
      r_260__46_ <= r_n_260__46_;
      r_260__45_ <= r_n_260__45_;
      r_260__44_ <= r_n_260__44_;
      r_260__43_ <= r_n_260__43_;
      r_260__42_ <= r_n_260__42_;
      r_260__41_ <= r_n_260__41_;
      r_260__40_ <= r_n_260__40_;
      r_260__39_ <= r_n_260__39_;
      r_260__38_ <= r_n_260__38_;
      r_260__37_ <= r_n_260__37_;
      r_260__36_ <= r_n_260__36_;
      r_260__35_ <= r_n_260__35_;
      r_260__34_ <= r_n_260__34_;
      r_260__33_ <= r_n_260__33_;
      r_260__32_ <= r_n_260__32_;
      r_260__31_ <= r_n_260__31_;
      r_260__30_ <= r_n_260__30_;
      r_260__29_ <= r_n_260__29_;
      r_260__28_ <= r_n_260__28_;
      r_260__27_ <= r_n_260__27_;
      r_260__26_ <= r_n_260__26_;
      r_260__25_ <= r_n_260__25_;
      r_260__24_ <= r_n_260__24_;
      r_260__23_ <= r_n_260__23_;
      r_260__22_ <= r_n_260__22_;
      r_260__21_ <= r_n_260__21_;
      r_260__20_ <= r_n_260__20_;
      r_260__19_ <= r_n_260__19_;
      r_260__18_ <= r_n_260__18_;
      r_260__17_ <= r_n_260__17_;
      r_260__16_ <= r_n_260__16_;
      r_260__15_ <= r_n_260__15_;
      r_260__14_ <= r_n_260__14_;
      r_260__13_ <= r_n_260__13_;
      r_260__12_ <= r_n_260__12_;
      r_260__11_ <= r_n_260__11_;
      r_260__10_ <= r_n_260__10_;
      r_260__9_ <= r_n_260__9_;
      r_260__8_ <= r_n_260__8_;
      r_260__7_ <= r_n_260__7_;
      r_260__6_ <= r_n_260__6_;
      r_260__5_ <= r_n_260__5_;
      r_260__4_ <= r_n_260__4_;
      r_260__3_ <= r_n_260__3_;
      r_260__2_ <= r_n_260__2_;
      r_260__1_ <= r_n_260__1_;
      r_260__0_ <= r_n_260__0_;
    end 
    if(N3845) begin
      r_261__63_ <= r_n_261__63_;
      r_261__62_ <= r_n_261__62_;
      r_261__61_ <= r_n_261__61_;
      r_261__60_ <= r_n_261__60_;
      r_261__59_ <= r_n_261__59_;
      r_261__58_ <= r_n_261__58_;
      r_261__57_ <= r_n_261__57_;
      r_261__56_ <= r_n_261__56_;
      r_261__55_ <= r_n_261__55_;
      r_261__54_ <= r_n_261__54_;
      r_261__53_ <= r_n_261__53_;
      r_261__52_ <= r_n_261__52_;
      r_261__51_ <= r_n_261__51_;
      r_261__50_ <= r_n_261__50_;
      r_261__49_ <= r_n_261__49_;
      r_261__48_ <= r_n_261__48_;
      r_261__47_ <= r_n_261__47_;
      r_261__46_ <= r_n_261__46_;
      r_261__45_ <= r_n_261__45_;
      r_261__44_ <= r_n_261__44_;
      r_261__43_ <= r_n_261__43_;
      r_261__42_ <= r_n_261__42_;
      r_261__41_ <= r_n_261__41_;
      r_261__40_ <= r_n_261__40_;
      r_261__39_ <= r_n_261__39_;
      r_261__38_ <= r_n_261__38_;
      r_261__37_ <= r_n_261__37_;
      r_261__36_ <= r_n_261__36_;
      r_261__35_ <= r_n_261__35_;
      r_261__34_ <= r_n_261__34_;
      r_261__33_ <= r_n_261__33_;
      r_261__32_ <= r_n_261__32_;
      r_261__31_ <= r_n_261__31_;
      r_261__30_ <= r_n_261__30_;
      r_261__29_ <= r_n_261__29_;
      r_261__28_ <= r_n_261__28_;
      r_261__27_ <= r_n_261__27_;
      r_261__26_ <= r_n_261__26_;
      r_261__25_ <= r_n_261__25_;
      r_261__24_ <= r_n_261__24_;
      r_261__23_ <= r_n_261__23_;
      r_261__22_ <= r_n_261__22_;
      r_261__21_ <= r_n_261__21_;
      r_261__20_ <= r_n_261__20_;
      r_261__19_ <= r_n_261__19_;
      r_261__18_ <= r_n_261__18_;
      r_261__17_ <= r_n_261__17_;
      r_261__16_ <= r_n_261__16_;
      r_261__15_ <= r_n_261__15_;
      r_261__14_ <= r_n_261__14_;
      r_261__13_ <= r_n_261__13_;
      r_261__12_ <= r_n_261__12_;
      r_261__11_ <= r_n_261__11_;
      r_261__10_ <= r_n_261__10_;
      r_261__9_ <= r_n_261__9_;
      r_261__8_ <= r_n_261__8_;
      r_261__7_ <= r_n_261__7_;
      r_261__6_ <= r_n_261__6_;
      r_261__5_ <= r_n_261__5_;
      r_261__4_ <= r_n_261__4_;
      r_261__3_ <= r_n_261__3_;
      r_261__2_ <= r_n_261__2_;
      r_261__1_ <= r_n_261__1_;
      r_261__0_ <= r_n_261__0_;
    end 
    if(N3846) begin
      r_262__63_ <= r_n_262__63_;
      r_262__62_ <= r_n_262__62_;
      r_262__61_ <= r_n_262__61_;
      r_262__60_ <= r_n_262__60_;
      r_262__59_ <= r_n_262__59_;
      r_262__58_ <= r_n_262__58_;
      r_262__57_ <= r_n_262__57_;
      r_262__56_ <= r_n_262__56_;
      r_262__55_ <= r_n_262__55_;
      r_262__54_ <= r_n_262__54_;
      r_262__53_ <= r_n_262__53_;
      r_262__52_ <= r_n_262__52_;
      r_262__51_ <= r_n_262__51_;
      r_262__50_ <= r_n_262__50_;
      r_262__49_ <= r_n_262__49_;
      r_262__48_ <= r_n_262__48_;
      r_262__47_ <= r_n_262__47_;
      r_262__46_ <= r_n_262__46_;
      r_262__45_ <= r_n_262__45_;
      r_262__44_ <= r_n_262__44_;
      r_262__43_ <= r_n_262__43_;
      r_262__42_ <= r_n_262__42_;
      r_262__41_ <= r_n_262__41_;
      r_262__40_ <= r_n_262__40_;
      r_262__39_ <= r_n_262__39_;
      r_262__38_ <= r_n_262__38_;
      r_262__37_ <= r_n_262__37_;
      r_262__36_ <= r_n_262__36_;
      r_262__35_ <= r_n_262__35_;
      r_262__34_ <= r_n_262__34_;
      r_262__33_ <= r_n_262__33_;
      r_262__32_ <= r_n_262__32_;
      r_262__31_ <= r_n_262__31_;
      r_262__30_ <= r_n_262__30_;
      r_262__29_ <= r_n_262__29_;
      r_262__28_ <= r_n_262__28_;
      r_262__27_ <= r_n_262__27_;
      r_262__26_ <= r_n_262__26_;
      r_262__25_ <= r_n_262__25_;
      r_262__24_ <= r_n_262__24_;
      r_262__23_ <= r_n_262__23_;
      r_262__22_ <= r_n_262__22_;
      r_262__21_ <= r_n_262__21_;
      r_262__20_ <= r_n_262__20_;
      r_262__19_ <= r_n_262__19_;
      r_262__18_ <= r_n_262__18_;
      r_262__17_ <= r_n_262__17_;
      r_262__16_ <= r_n_262__16_;
      r_262__15_ <= r_n_262__15_;
      r_262__14_ <= r_n_262__14_;
      r_262__13_ <= r_n_262__13_;
      r_262__12_ <= r_n_262__12_;
      r_262__11_ <= r_n_262__11_;
      r_262__10_ <= r_n_262__10_;
      r_262__9_ <= r_n_262__9_;
      r_262__8_ <= r_n_262__8_;
      r_262__7_ <= r_n_262__7_;
      r_262__6_ <= r_n_262__6_;
      r_262__5_ <= r_n_262__5_;
      r_262__4_ <= r_n_262__4_;
      r_262__3_ <= r_n_262__3_;
      r_262__2_ <= r_n_262__2_;
      r_262__1_ <= r_n_262__1_;
      r_262__0_ <= r_n_262__0_;
    end 
    if(N3847) begin
      r_263__63_ <= r_n_263__63_;
      r_263__62_ <= r_n_263__62_;
      r_263__61_ <= r_n_263__61_;
      r_263__60_ <= r_n_263__60_;
      r_263__59_ <= r_n_263__59_;
      r_263__58_ <= r_n_263__58_;
      r_263__57_ <= r_n_263__57_;
      r_263__56_ <= r_n_263__56_;
      r_263__55_ <= r_n_263__55_;
      r_263__54_ <= r_n_263__54_;
      r_263__53_ <= r_n_263__53_;
      r_263__52_ <= r_n_263__52_;
      r_263__51_ <= r_n_263__51_;
      r_263__50_ <= r_n_263__50_;
      r_263__49_ <= r_n_263__49_;
      r_263__48_ <= r_n_263__48_;
      r_263__47_ <= r_n_263__47_;
      r_263__46_ <= r_n_263__46_;
      r_263__45_ <= r_n_263__45_;
      r_263__44_ <= r_n_263__44_;
      r_263__43_ <= r_n_263__43_;
      r_263__42_ <= r_n_263__42_;
      r_263__41_ <= r_n_263__41_;
      r_263__40_ <= r_n_263__40_;
      r_263__39_ <= r_n_263__39_;
      r_263__38_ <= r_n_263__38_;
      r_263__37_ <= r_n_263__37_;
      r_263__36_ <= r_n_263__36_;
      r_263__35_ <= r_n_263__35_;
      r_263__34_ <= r_n_263__34_;
      r_263__33_ <= r_n_263__33_;
      r_263__32_ <= r_n_263__32_;
      r_263__31_ <= r_n_263__31_;
      r_263__30_ <= r_n_263__30_;
      r_263__29_ <= r_n_263__29_;
      r_263__28_ <= r_n_263__28_;
      r_263__27_ <= r_n_263__27_;
      r_263__26_ <= r_n_263__26_;
      r_263__25_ <= r_n_263__25_;
      r_263__24_ <= r_n_263__24_;
      r_263__23_ <= r_n_263__23_;
      r_263__22_ <= r_n_263__22_;
      r_263__21_ <= r_n_263__21_;
      r_263__20_ <= r_n_263__20_;
      r_263__19_ <= r_n_263__19_;
      r_263__18_ <= r_n_263__18_;
      r_263__17_ <= r_n_263__17_;
      r_263__16_ <= r_n_263__16_;
      r_263__15_ <= r_n_263__15_;
      r_263__14_ <= r_n_263__14_;
      r_263__13_ <= r_n_263__13_;
      r_263__12_ <= r_n_263__12_;
      r_263__11_ <= r_n_263__11_;
      r_263__10_ <= r_n_263__10_;
      r_263__9_ <= r_n_263__9_;
      r_263__8_ <= r_n_263__8_;
      r_263__7_ <= r_n_263__7_;
      r_263__6_ <= r_n_263__6_;
      r_263__5_ <= r_n_263__5_;
      r_263__4_ <= r_n_263__4_;
      r_263__3_ <= r_n_263__3_;
      r_263__2_ <= r_n_263__2_;
      r_263__1_ <= r_n_263__1_;
      r_263__0_ <= r_n_263__0_;
    end 
    if(N3848) begin
      r_264__63_ <= r_n_264__63_;
      r_264__62_ <= r_n_264__62_;
      r_264__61_ <= r_n_264__61_;
      r_264__60_ <= r_n_264__60_;
      r_264__59_ <= r_n_264__59_;
      r_264__58_ <= r_n_264__58_;
      r_264__57_ <= r_n_264__57_;
      r_264__56_ <= r_n_264__56_;
      r_264__55_ <= r_n_264__55_;
      r_264__54_ <= r_n_264__54_;
      r_264__53_ <= r_n_264__53_;
      r_264__52_ <= r_n_264__52_;
      r_264__51_ <= r_n_264__51_;
      r_264__50_ <= r_n_264__50_;
      r_264__49_ <= r_n_264__49_;
      r_264__48_ <= r_n_264__48_;
      r_264__47_ <= r_n_264__47_;
      r_264__46_ <= r_n_264__46_;
      r_264__45_ <= r_n_264__45_;
      r_264__44_ <= r_n_264__44_;
      r_264__43_ <= r_n_264__43_;
      r_264__42_ <= r_n_264__42_;
      r_264__41_ <= r_n_264__41_;
      r_264__40_ <= r_n_264__40_;
      r_264__39_ <= r_n_264__39_;
      r_264__38_ <= r_n_264__38_;
      r_264__37_ <= r_n_264__37_;
      r_264__36_ <= r_n_264__36_;
      r_264__35_ <= r_n_264__35_;
      r_264__34_ <= r_n_264__34_;
      r_264__33_ <= r_n_264__33_;
      r_264__32_ <= r_n_264__32_;
      r_264__31_ <= r_n_264__31_;
      r_264__30_ <= r_n_264__30_;
      r_264__29_ <= r_n_264__29_;
      r_264__28_ <= r_n_264__28_;
      r_264__27_ <= r_n_264__27_;
      r_264__26_ <= r_n_264__26_;
      r_264__25_ <= r_n_264__25_;
      r_264__24_ <= r_n_264__24_;
      r_264__23_ <= r_n_264__23_;
      r_264__22_ <= r_n_264__22_;
      r_264__21_ <= r_n_264__21_;
      r_264__20_ <= r_n_264__20_;
      r_264__19_ <= r_n_264__19_;
      r_264__18_ <= r_n_264__18_;
      r_264__17_ <= r_n_264__17_;
      r_264__16_ <= r_n_264__16_;
      r_264__15_ <= r_n_264__15_;
      r_264__14_ <= r_n_264__14_;
      r_264__13_ <= r_n_264__13_;
      r_264__12_ <= r_n_264__12_;
      r_264__11_ <= r_n_264__11_;
      r_264__10_ <= r_n_264__10_;
      r_264__9_ <= r_n_264__9_;
      r_264__8_ <= r_n_264__8_;
      r_264__7_ <= r_n_264__7_;
      r_264__6_ <= r_n_264__6_;
      r_264__5_ <= r_n_264__5_;
      r_264__4_ <= r_n_264__4_;
      r_264__3_ <= r_n_264__3_;
      r_264__2_ <= r_n_264__2_;
      r_264__1_ <= r_n_264__1_;
      r_264__0_ <= r_n_264__0_;
    end 
    if(N3849) begin
      r_265__63_ <= r_n_265__63_;
      r_265__62_ <= r_n_265__62_;
      r_265__61_ <= r_n_265__61_;
      r_265__60_ <= r_n_265__60_;
      r_265__59_ <= r_n_265__59_;
      r_265__58_ <= r_n_265__58_;
      r_265__57_ <= r_n_265__57_;
      r_265__56_ <= r_n_265__56_;
      r_265__55_ <= r_n_265__55_;
      r_265__54_ <= r_n_265__54_;
      r_265__53_ <= r_n_265__53_;
      r_265__52_ <= r_n_265__52_;
      r_265__51_ <= r_n_265__51_;
      r_265__50_ <= r_n_265__50_;
      r_265__49_ <= r_n_265__49_;
      r_265__48_ <= r_n_265__48_;
      r_265__47_ <= r_n_265__47_;
      r_265__46_ <= r_n_265__46_;
      r_265__45_ <= r_n_265__45_;
      r_265__44_ <= r_n_265__44_;
      r_265__43_ <= r_n_265__43_;
      r_265__42_ <= r_n_265__42_;
      r_265__41_ <= r_n_265__41_;
      r_265__40_ <= r_n_265__40_;
      r_265__39_ <= r_n_265__39_;
      r_265__38_ <= r_n_265__38_;
      r_265__37_ <= r_n_265__37_;
      r_265__36_ <= r_n_265__36_;
      r_265__35_ <= r_n_265__35_;
      r_265__34_ <= r_n_265__34_;
      r_265__33_ <= r_n_265__33_;
      r_265__32_ <= r_n_265__32_;
      r_265__31_ <= r_n_265__31_;
      r_265__30_ <= r_n_265__30_;
      r_265__29_ <= r_n_265__29_;
      r_265__28_ <= r_n_265__28_;
      r_265__27_ <= r_n_265__27_;
      r_265__26_ <= r_n_265__26_;
      r_265__25_ <= r_n_265__25_;
      r_265__24_ <= r_n_265__24_;
      r_265__23_ <= r_n_265__23_;
      r_265__22_ <= r_n_265__22_;
      r_265__21_ <= r_n_265__21_;
      r_265__20_ <= r_n_265__20_;
      r_265__19_ <= r_n_265__19_;
      r_265__18_ <= r_n_265__18_;
      r_265__17_ <= r_n_265__17_;
      r_265__16_ <= r_n_265__16_;
      r_265__15_ <= r_n_265__15_;
      r_265__14_ <= r_n_265__14_;
      r_265__13_ <= r_n_265__13_;
      r_265__12_ <= r_n_265__12_;
      r_265__11_ <= r_n_265__11_;
      r_265__10_ <= r_n_265__10_;
      r_265__9_ <= r_n_265__9_;
      r_265__8_ <= r_n_265__8_;
      r_265__7_ <= r_n_265__7_;
      r_265__6_ <= r_n_265__6_;
      r_265__5_ <= r_n_265__5_;
      r_265__4_ <= r_n_265__4_;
      r_265__3_ <= r_n_265__3_;
      r_265__2_ <= r_n_265__2_;
      r_265__1_ <= r_n_265__1_;
      r_265__0_ <= r_n_265__0_;
    end 
    if(N3850) begin
      r_266__63_ <= r_n_266__63_;
      r_266__62_ <= r_n_266__62_;
      r_266__61_ <= r_n_266__61_;
      r_266__60_ <= r_n_266__60_;
      r_266__59_ <= r_n_266__59_;
      r_266__58_ <= r_n_266__58_;
      r_266__57_ <= r_n_266__57_;
      r_266__56_ <= r_n_266__56_;
      r_266__55_ <= r_n_266__55_;
      r_266__54_ <= r_n_266__54_;
      r_266__53_ <= r_n_266__53_;
      r_266__52_ <= r_n_266__52_;
      r_266__51_ <= r_n_266__51_;
      r_266__50_ <= r_n_266__50_;
      r_266__49_ <= r_n_266__49_;
      r_266__48_ <= r_n_266__48_;
      r_266__47_ <= r_n_266__47_;
      r_266__46_ <= r_n_266__46_;
      r_266__45_ <= r_n_266__45_;
      r_266__44_ <= r_n_266__44_;
      r_266__43_ <= r_n_266__43_;
      r_266__42_ <= r_n_266__42_;
      r_266__41_ <= r_n_266__41_;
      r_266__40_ <= r_n_266__40_;
      r_266__39_ <= r_n_266__39_;
      r_266__38_ <= r_n_266__38_;
      r_266__37_ <= r_n_266__37_;
      r_266__36_ <= r_n_266__36_;
      r_266__35_ <= r_n_266__35_;
      r_266__34_ <= r_n_266__34_;
      r_266__33_ <= r_n_266__33_;
      r_266__32_ <= r_n_266__32_;
      r_266__31_ <= r_n_266__31_;
      r_266__30_ <= r_n_266__30_;
      r_266__29_ <= r_n_266__29_;
      r_266__28_ <= r_n_266__28_;
      r_266__27_ <= r_n_266__27_;
      r_266__26_ <= r_n_266__26_;
      r_266__25_ <= r_n_266__25_;
      r_266__24_ <= r_n_266__24_;
      r_266__23_ <= r_n_266__23_;
      r_266__22_ <= r_n_266__22_;
      r_266__21_ <= r_n_266__21_;
      r_266__20_ <= r_n_266__20_;
      r_266__19_ <= r_n_266__19_;
      r_266__18_ <= r_n_266__18_;
      r_266__17_ <= r_n_266__17_;
      r_266__16_ <= r_n_266__16_;
      r_266__15_ <= r_n_266__15_;
      r_266__14_ <= r_n_266__14_;
      r_266__13_ <= r_n_266__13_;
      r_266__12_ <= r_n_266__12_;
      r_266__11_ <= r_n_266__11_;
      r_266__10_ <= r_n_266__10_;
      r_266__9_ <= r_n_266__9_;
      r_266__8_ <= r_n_266__8_;
      r_266__7_ <= r_n_266__7_;
      r_266__6_ <= r_n_266__6_;
      r_266__5_ <= r_n_266__5_;
      r_266__4_ <= r_n_266__4_;
      r_266__3_ <= r_n_266__3_;
      r_266__2_ <= r_n_266__2_;
      r_266__1_ <= r_n_266__1_;
      r_266__0_ <= r_n_266__0_;
    end 
    if(N3851) begin
      r_267__63_ <= r_n_267__63_;
      r_267__62_ <= r_n_267__62_;
      r_267__61_ <= r_n_267__61_;
      r_267__60_ <= r_n_267__60_;
      r_267__59_ <= r_n_267__59_;
      r_267__58_ <= r_n_267__58_;
      r_267__57_ <= r_n_267__57_;
      r_267__56_ <= r_n_267__56_;
      r_267__55_ <= r_n_267__55_;
      r_267__54_ <= r_n_267__54_;
      r_267__53_ <= r_n_267__53_;
      r_267__52_ <= r_n_267__52_;
      r_267__51_ <= r_n_267__51_;
      r_267__50_ <= r_n_267__50_;
      r_267__49_ <= r_n_267__49_;
      r_267__48_ <= r_n_267__48_;
      r_267__47_ <= r_n_267__47_;
      r_267__46_ <= r_n_267__46_;
      r_267__45_ <= r_n_267__45_;
      r_267__44_ <= r_n_267__44_;
      r_267__43_ <= r_n_267__43_;
      r_267__42_ <= r_n_267__42_;
      r_267__41_ <= r_n_267__41_;
      r_267__40_ <= r_n_267__40_;
      r_267__39_ <= r_n_267__39_;
      r_267__38_ <= r_n_267__38_;
      r_267__37_ <= r_n_267__37_;
      r_267__36_ <= r_n_267__36_;
      r_267__35_ <= r_n_267__35_;
      r_267__34_ <= r_n_267__34_;
      r_267__33_ <= r_n_267__33_;
      r_267__32_ <= r_n_267__32_;
      r_267__31_ <= r_n_267__31_;
      r_267__30_ <= r_n_267__30_;
      r_267__29_ <= r_n_267__29_;
      r_267__28_ <= r_n_267__28_;
      r_267__27_ <= r_n_267__27_;
      r_267__26_ <= r_n_267__26_;
      r_267__25_ <= r_n_267__25_;
      r_267__24_ <= r_n_267__24_;
      r_267__23_ <= r_n_267__23_;
      r_267__22_ <= r_n_267__22_;
      r_267__21_ <= r_n_267__21_;
      r_267__20_ <= r_n_267__20_;
      r_267__19_ <= r_n_267__19_;
      r_267__18_ <= r_n_267__18_;
      r_267__17_ <= r_n_267__17_;
      r_267__16_ <= r_n_267__16_;
      r_267__15_ <= r_n_267__15_;
      r_267__14_ <= r_n_267__14_;
      r_267__13_ <= r_n_267__13_;
      r_267__12_ <= r_n_267__12_;
      r_267__11_ <= r_n_267__11_;
      r_267__10_ <= r_n_267__10_;
      r_267__9_ <= r_n_267__9_;
      r_267__8_ <= r_n_267__8_;
      r_267__7_ <= r_n_267__7_;
      r_267__6_ <= r_n_267__6_;
      r_267__5_ <= r_n_267__5_;
      r_267__4_ <= r_n_267__4_;
      r_267__3_ <= r_n_267__3_;
      r_267__2_ <= r_n_267__2_;
      r_267__1_ <= r_n_267__1_;
      r_267__0_ <= r_n_267__0_;
    end 
    if(N3852) begin
      r_268__63_ <= r_n_268__63_;
      r_268__62_ <= r_n_268__62_;
      r_268__61_ <= r_n_268__61_;
      r_268__60_ <= r_n_268__60_;
      r_268__59_ <= r_n_268__59_;
      r_268__58_ <= r_n_268__58_;
      r_268__57_ <= r_n_268__57_;
      r_268__56_ <= r_n_268__56_;
      r_268__55_ <= r_n_268__55_;
      r_268__54_ <= r_n_268__54_;
      r_268__53_ <= r_n_268__53_;
      r_268__52_ <= r_n_268__52_;
      r_268__51_ <= r_n_268__51_;
      r_268__50_ <= r_n_268__50_;
      r_268__49_ <= r_n_268__49_;
      r_268__48_ <= r_n_268__48_;
      r_268__47_ <= r_n_268__47_;
      r_268__46_ <= r_n_268__46_;
      r_268__45_ <= r_n_268__45_;
      r_268__44_ <= r_n_268__44_;
      r_268__43_ <= r_n_268__43_;
      r_268__42_ <= r_n_268__42_;
      r_268__41_ <= r_n_268__41_;
      r_268__40_ <= r_n_268__40_;
      r_268__39_ <= r_n_268__39_;
      r_268__38_ <= r_n_268__38_;
      r_268__37_ <= r_n_268__37_;
      r_268__36_ <= r_n_268__36_;
      r_268__35_ <= r_n_268__35_;
      r_268__34_ <= r_n_268__34_;
      r_268__33_ <= r_n_268__33_;
      r_268__32_ <= r_n_268__32_;
      r_268__31_ <= r_n_268__31_;
      r_268__30_ <= r_n_268__30_;
      r_268__29_ <= r_n_268__29_;
      r_268__28_ <= r_n_268__28_;
      r_268__27_ <= r_n_268__27_;
      r_268__26_ <= r_n_268__26_;
      r_268__25_ <= r_n_268__25_;
      r_268__24_ <= r_n_268__24_;
      r_268__23_ <= r_n_268__23_;
      r_268__22_ <= r_n_268__22_;
      r_268__21_ <= r_n_268__21_;
      r_268__20_ <= r_n_268__20_;
      r_268__19_ <= r_n_268__19_;
      r_268__18_ <= r_n_268__18_;
      r_268__17_ <= r_n_268__17_;
      r_268__16_ <= r_n_268__16_;
      r_268__15_ <= r_n_268__15_;
      r_268__14_ <= r_n_268__14_;
      r_268__13_ <= r_n_268__13_;
      r_268__12_ <= r_n_268__12_;
      r_268__11_ <= r_n_268__11_;
      r_268__10_ <= r_n_268__10_;
      r_268__9_ <= r_n_268__9_;
      r_268__8_ <= r_n_268__8_;
      r_268__7_ <= r_n_268__7_;
      r_268__6_ <= r_n_268__6_;
      r_268__5_ <= r_n_268__5_;
      r_268__4_ <= r_n_268__4_;
      r_268__3_ <= r_n_268__3_;
      r_268__2_ <= r_n_268__2_;
      r_268__1_ <= r_n_268__1_;
      r_268__0_ <= r_n_268__0_;
    end 
    if(N3853) begin
      r_269__63_ <= r_n_269__63_;
      r_269__62_ <= r_n_269__62_;
      r_269__61_ <= r_n_269__61_;
      r_269__60_ <= r_n_269__60_;
      r_269__59_ <= r_n_269__59_;
      r_269__58_ <= r_n_269__58_;
      r_269__57_ <= r_n_269__57_;
      r_269__56_ <= r_n_269__56_;
      r_269__55_ <= r_n_269__55_;
      r_269__54_ <= r_n_269__54_;
      r_269__53_ <= r_n_269__53_;
      r_269__52_ <= r_n_269__52_;
      r_269__51_ <= r_n_269__51_;
      r_269__50_ <= r_n_269__50_;
      r_269__49_ <= r_n_269__49_;
      r_269__48_ <= r_n_269__48_;
      r_269__47_ <= r_n_269__47_;
      r_269__46_ <= r_n_269__46_;
      r_269__45_ <= r_n_269__45_;
      r_269__44_ <= r_n_269__44_;
      r_269__43_ <= r_n_269__43_;
      r_269__42_ <= r_n_269__42_;
      r_269__41_ <= r_n_269__41_;
      r_269__40_ <= r_n_269__40_;
      r_269__39_ <= r_n_269__39_;
      r_269__38_ <= r_n_269__38_;
      r_269__37_ <= r_n_269__37_;
      r_269__36_ <= r_n_269__36_;
      r_269__35_ <= r_n_269__35_;
      r_269__34_ <= r_n_269__34_;
      r_269__33_ <= r_n_269__33_;
      r_269__32_ <= r_n_269__32_;
      r_269__31_ <= r_n_269__31_;
      r_269__30_ <= r_n_269__30_;
      r_269__29_ <= r_n_269__29_;
      r_269__28_ <= r_n_269__28_;
      r_269__27_ <= r_n_269__27_;
      r_269__26_ <= r_n_269__26_;
      r_269__25_ <= r_n_269__25_;
      r_269__24_ <= r_n_269__24_;
      r_269__23_ <= r_n_269__23_;
      r_269__22_ <= r_n_269__22_;
      r_269__21_ <= r_n_269__21_;
      r_269__20_ <= r_n_269__20_;
      r_269__19_ <= r_n_269__19_;
      r_269__18_ <= r_n_269__18_;
      r_269__17_ <= r_n_269__17_;
      r_269__16_ <= r_n_269__16_;
      r_269__15_ <= r_n_269__15_;
      r_269__14_ <= r_n_269__14_;
      r_269__13_ <= r_n_269__13_;
      r_269__12_ <= r_n_269__12_;
      r_269__11_ <= r_n_269__11_;
      r_269__10_ <= r_n_269__10_;
      r_269__9_ <= r_n_269__9_;
      r_269__8_ <= r_n_269__8_;
      r_269__7_ <= r_n_269__7_;
      r_269__6_ <= r_n_269__6_;
      r_269__5_ <= r_n_269__5_;
      r_269__4_ <= r_n_269__4_;
      r_269__3_ <= r_n_269__3_;
      r_269__2_ <= r_n_269__2_;
      r_269__1_ <= r_n_269__1_;
      r_269__0_ <= r_n_269__0_;
    end 
    if(N3854) begin
      r_270__63_ <= r_n_270__63_;
      r_270__62_ <= r_n_270__62_;
      r_270__61_ <= r_n_270__61_;
      r_270__60_ <= r_n_270__60_;
      r_270__59_ <= r_n_270__59_;
      r_270__58_ <= r_n_270__58_;
      r_270__57_ <= r_n_270__57_;
      r_270__56_ <= r_n_270__56_;
      r_270__55_ <= r_n_270__55_;
      r_270__54_ <= r_n_270__54_;
      r_270__53_ <= r_n_270__53_;
      r_270__52_ <= r_n_270__52_;
      r_270__51_ <= r_n_270__51_;
      r_270__50_ <= r_n_270__50_;
      r_270__49_ <= r_n_270__49_;
      r_270__48_ <= r_n_270__48_;
      r_270__47_ <= r_n_270__47_;
      r_270__46_ <= r_n_270__46_;
      r_270__45_ <= r_n_270__45_;
      r_270__44_ <= r_n_270__44_;
      r_270__43_ <= r_n_270__43_;
      r_270__42_ <= r_n_270__42_;
      r_270__41_ <= r_n_270__41_;
      r_270__40_ <= r_n_270__40_;
      r_270__39_ <= r_n_270__39_;
      r_270__38_ <= r_n_270__38_;
      r_270__37_ <= r_n_270__37_;
      r_270__36_ <= r_n_270__36_;
      r_270__35_ <= r_n_270__35_;
      r_270__34_ <= r_n_270__34_;
      r_270__33_ <= r_n_270__33_;
      r_270__32_ <= r_n_270__32_;
      r_270__31_ <= r_n_270__31_;
      r_270__30_ <= r_n_270__30_;
      r_270__29_ <= r_n_270__29_;
      r_270__28_ <= r_n_270__28_;
      r_270__27_ <= r_n_270__27_;
      r_270__26_ <= r_n_270__26_;
      r_270__25_ <= r_n_270__25_;
      r_270__24_ <= r_n_270__24_;
      r_270__23_ <= r_n_270__23_;
      r_270__22_ <= r_n_270__22_;
      r_270__21_ <= r_n_270__21_;
      r_270__20_ <= r_n_270__20_;
      r_270__19_ <= r_n_270__19_;
      r_270__18_ <= r_n_270__18_;
      r_270__17_ <= r_n_270__17_;
      r_270__16_ <= r_n_270__16_;
      r_270__15_ <= r_n_270__15_;
      r_270__14_ <= r_n_270__14_;
      r_270__13_ <= r_n_270__13_;
      r_270__12_ <= r_n_270__12_;
      r_270__11_ <= r_n_270__11_;
      r_270__10_ <= r_n_270__10_;
      r_270__9_ <= r_n_270__9_;
      r_270__8_ <= r_n_270__8_;
      r_270__7_ <= r_n_270__7_;
      r_270__6_ <= r_n_270__6_;
      r_270__5_ <= r_n_270__5_;
      r_270__4_ <= r_n_270__4_;
      r_270__3_ <= r_n_270__3_;
      r_270__2_ <= r_n_270__2_;
      r_270__1_ <= r_n_270__1_;
      r_270__0_ <= r_n_270__0_;
    end 
    if(N3855) begin
      r_271__63_ <= r_n_271__63_;
      r_271__62_ <= r_n_271__62_;
      r_271__61_ <= r_n_271__61_;
      r_271__60_ <= r_n_271__60_;
      r_271__59_ <= r_n_271__59_;
      r_271__58_ <= r_n_271__58_;
      r_271__57_ <= r_n_271__57_;
      r_271__56_ <= r_n_271__56_;
      r_271__55_ <= r_n_271__55_;
      r_271__54_ <= r_n_271__54_;
      r_271__53_ <= r_n_271__53_;
      r_271__52_ <= r_n_271__52_;
      r_271__51_ <= r_n_271__51_;
      r_271__50_ <= r_n_271__50_;
      r_271__49_ <= r_n_271__49_;
      r_271__48_ <= r_n_271__48_;
      r_271__47_ <= r_n_271__47_;
      r_271__46_ <= r_n_271__46_;
      r_271__45_ <= r_n_271__45_;
      r_271__44_ <= r_n_271__44_;
      r_271__43_ <= r_n_271__43_;
      r_271__42_ <= r_n_271__42_;
      r_271__41_ <= r_n_271__41_;
      r_271__40_ <= r_n_271__40_;
      r_271__39_ <= r_n_271__39_;
      r_271__38_ <= r_n_271__38_;
      r_271__37_ <= r_n_271__37_;
      r_271__36_ <= r_n_271__36_;
      r_271__35_ <= r_n_271__35_;
      r_271__34_ <= r_n_271__34_;
      r_271__33_ <= r_n_271__33_;
      r_271__32_ <= r_n_271__32_;
      r_271__31_ <= r_n_271__31_;
      r_271__30_ <= r_n_271__30_;
      r_271__29_ <= r_n_271__29_;
      r_271__28_ <= r_n_271__28_;
      r_271__27_ <= r_n_271__27_;
      r_271__26_ <= r_n_271__26_;
      r_271__25_ <= r_n_271__25_;
      r_271__24_ <= r_n_271__24_;
      r_271__23_ <= r_n_271__23_;
      r_271__22_ <= r_n_271__22_;
      r_271__21_ <= r_n_271__21_;
      r_271__20_ <= r_n_271__20_;
      r_271__19_ <= r_n_271__19_;
      r_271__18_ <= r_n_271__18_;
      r_271__17_ <= r_n_271__17_;
      r_271__16_ <= r_n_271__16_;
      r_271__15_ <= r_n_271__15_;
      r_271__14_ <= r_n_271__14_;
      r_271__13_ <= r_n_271__13_;
      r_271__12_ <= r_n_271__12_;
      r_271__11_ <= r_n_271__11_;
      r_271__10_ <= r_n_271__10_;
      r_271__9_ <= r_n_271__9_;
      r_271__8_ <= r_n_271__8_;
      r_271__7_ <= r_n_271__7_;
      r_271__6_ <= r_n_271__6_;
      r_271__5_ <= r_n_271__5_;
      r_271__4_ <= r_n_271__4_;
      r_271__3_ <= r_n_271__3_;
      r_271__2_ <= r_n_271__2_;
      r_271__1_ <= r_n_271__1_;
      r_271__0_ <= r_n_271__0_;
    end 
    if(N3856) begin
      r_272__63_ <= r_n_272__63_;
      r_272__62_ <= r_n_272__62_;
      r_272__61_ <= r_n_272__61_;
      r_272__60_ <= r_n_272__60_;
      r_272__59_ <= r_n_272__59_;
      r_272__58_ <= r_n_272__58_;
      r_272__57_ <= r_n_272__57_;
      r_272__56_ <= r_n_272__56_;
      r_272__55_ <= r_n_272__55_;
      r_272__54_ <= r_n_272__54_;
      r_272__53_ <= r_n_272__53_;
      r_272__52_ <= r_n_272__52_;
      r_272__51_ <= r_n_272__51_;
      r_272__50_ <= r_n_272__50_;
      r_272__49_ <= r_n_272__49_;
      r_272__48_ <= r_n_272__48_;
      r_272__47_ <= r_n_272__47_;
      r_272__46_ <= r_n_272__46_;
      r_272__45_ <= r_n_272__45_;
      r_272__44_ <= r_n_272__44_;
      r_272__43_ <= r_n_272__43_;
      r_272__42_ <= r_n_272__42_;
      r_272__41_ <= r_n_272__41_;
      r_272__40_ <= r_n_272__40_;
      r_272__39_ <= r_n_272__39_;
      r_272__38_ <= r_n_272__38_;
      r_272__37_ <= r_n_272__37_;
      r_272__36_ <= r_n_272__36_;
      r_272__35_ <= r_n_272__35_;
      r_272__34_ <= r_n_272__34_;
      r_272__33_ <= r_n_272__33_;
      r_272__32_ <= r_n_272__32_;
      r_272__31_ <= r_n_272__31_;
      r_272__30_ <= r_n_272__30_;
      r_272__29_ <= r_n_272__29_;
      r_272__28_ <= r_n_272__28_;
      r_272__27_ <= r_n_272__27_;
      r_272__26_ <= r_n_272__26_;
      r_272__25_ <= r_n_272__25_;
      r_272__24_ <= r_n_272__24_;
      r_272__23_ <= r_n_272__23_;
      r_272__22_ <= r_n_272__22_;
      r_272__21_ <= r_n_272__21_;
      r_272__20_ <= r_n_272__20_;
      r_272__19_ <= r_n_272__19_;
      r_272__18_ <= r_n_272__18_;
      r_272__17_ <= r_n_272__17_;
      r_272__16_ <= r_n_272__16_;
      r_272__15_ <= r_n_272__15_;
      r_272__14_ <= r_n_272__14_;
      r_272__13_ <= r_n_272__13_;
      r_272__12_ <= r_n_272__12_;
      r_272__11_ <= r_n_272__11_;
      r_272__10_ <= r_n_272__10_;
      r_272__9_ <= r_n_272__9_;
      r_272__8_ <= r_n_272__8_;
      r_272__7_ <= r_n_272__7_;
      r_272__6_ <= r_n_272__6_;
      r_272__5_ <= r_n_272__5_;
      r_272__4_ <= r_n_272__4_;
      r_272__3_ <= r_n_272__3_;
      r_272__2_ <= r_n_272__2_;
      r_272__1_ <= r_n_272__1_;
      r_272__0_ <= r_n_272__0_;
    end 
    if(N3857) begin
      r_273__63_ <= r_n_273__63_;
      r_273__62_ <= r_n_273__62_;
      r_273__61_ <= r_n_273__61_;
      r_273__60_ <= r_n_273__60_;
      r_273__59_ <= r_n_273__59_;
      r_273__58_ <= r_n_273__58_;
      r_273__57_ <= r_n_273__57_;
      r_273__56_ <= r_n_273__56_;
      r_273__55_ <= r_n_273__55_;
      r_273__54_ <= r_n_273__54_;
      r_273__53_ <= r_n_273__53_;
      r_273__52_ <= r_n_273__52_;
      r_273__51_ <= r_n_273__51_;
      r_273__50_ <= r_n_273__50_;
      r_273__49_ <= r_n_273__49_;
      r_273__48_ <= r_n_273__48_;
      r_273__47_ <= r_n_273__47_;
      r_273__46_ <= r_n_273__46_;
      r_273__45_ <= r_n_273__45_;
      r_273__44_ <= r_n_273__44_;
      r_273__43_ <= r_n_273__43_;
      r_273__42_ <= r_n_273__42_;
      r_273__41_ <= r_n_273__41_;
      r_273__40_ <= r_n_273__40_;
      r_273__39_ <= r_n_273__39_;
      r_273__38_ <= r_n_273__38_;
      r_273__37_ <= r_n_273__37_;
      r_273__36_ <= r_n_273__36_;
      r_273__35_ <= r_n_273__35_;
      r_273__34_ <= r_n_273__34_;
      r_273__33_ <= r_n_273__33_;
      r_273__32_ <= r_n_273__32_;
      r_273__31_ <= r_n_273__31_;
      r_273__30_ <= r_n_273__30_;
      r_273__29_ <= r_n_273__29_;
      r_273__28_ <= r_n_273__28_;
      r_273__27_ <= r_n_273__27_;
      r_273__26_ <= r_n_273__26_;
      r_273__25_ <= r_n_273__25_;
      r_273__24_ <= r_n_273__24_;
      r_273__23_ <= r_n_273__23_;
      r_273__22_ <= r_n_273__22_;
      r_273__21_ <= r_n_273__21_;
      r_273__20_ <= r_n_273__20_;
      r_273__19_ <= r_n_273__19_;
      r_273__18_ <= r_n_273__18_;
      r_273__17_ <= r_n_273__17_;
      r_273__16_ <= r_n_273__16_;
      r_273__15_ <= r_n_273__15_;
      r_273__14_ <= r_n_273__14_;
      r_273__13_ <= r_n_273__13_;
      r_273__12_ <= r_n_273__12_;
      r_273__11_ <= r_n_273__11_;
      r_273__10_ <= r_n_273__10_;
      r_273__9_ <= r_n_273__9_;
      r_273__8_ <= r_n_273__8_;
      r_273__7_ <= r_n_273__7_;
      r_273__6_ <= r_n_273__6_;
      r_273__5_ <= r_n_273__5_;
      r_273__4_ <= r_n_273__4_;
      r_273__3_ <= r_n_273__3_;
      r_273__2_ <= r_n_273__2_;
      r_273__1_ <= r_n_273__1_;
      r_273__0_ <= r_n_273__0_;
    end 
    if(N3858) begin
      r_274__63_ <= r_n_274__63_;
      r_274__62_ <= r_n_274__62_;
      r_274__61_ <= r_n_274__61_;
      r_274__60_ <= r_n_274__60_;
      r_274__59_ <= r_n_274__59_;
      r_274__58_ <= r_n_274__58_;
      r_274__57_ <= r_n_274__57_;
      r_274__56_ <= r_n_274__56_;
      r_274__55_ <= r_n_274__55_;
      r_274__54_ <= r_n_274__54_;
      r_274__53_ <= r_n_274__53_;
      r_274__52_ <= r_n_274__52_;
      r_274__51_ <= r_n_274__51_;
      r_274__50_ <= r_n_274__50_;
      r_274__49_ <= r_n_274__49_;
      r_274__48_ <= r_n_274__48_;
      r_274__47_ <= r_n_274__47_;
      r_274__46_ <= r_n_274__46_;
      r_274__45_ <= r_n_274__45_;
      r_274__44_ <= r_n_274__44_;
      r_274__43_ <= r_n_274__43_;
      r_274__42_ <= r_n_274__42_;
      r_274__41_ <= r_n_274__41_;
      r_274__40_ <= r_n_274__40_;
      r_274__39_ <= r_n_274__39_;
      r_274__38_ <= r_n_274__38_;
      r_274__37_ <= r_n_274__37_;
      r_274__36_ <= r_n_274__36_;
      r_274__35_ <= r_n_274__35_;
      r_274__34_ <= r_n_274__34_;
      r_274__33_ <= r_n_274__33_;
      r_274__32_ <= r_n_274__32_;
      r_274__31_ <= r_n_274__31_;
      r_274__30_ <= r_n_274__30_;
      r_274__29_ <= r_n_274__29_;
      r_274__28_ <= r_n_274__28_;
      r_274__27_ <= r_n_274__27_;
      r_274__26_ <= r_n_274__26_;
      r_274__25_ <= r_n_274__25_;
      r_274__24_ <= r_n_274__24_;
      r_274__23_ <= r_n_274__23_;
      r_274__22_ <= r_n_274__22_;
      r_274__21_ <= r_n_274__21_;
      r_274__20_ <= r_n_274__20_;
      r_274__19_ <= r_n_274__19_;
      r_274__18_ <= r_n_274__18_;
      r_274__17_ <= r_n_274__17_;
      r_274__16_ <= r_n_274__16_;
      r_274__15_ <= r_n_274__15_;
      r_274__14_ <= r_n_274__14_;
      r_274__13_ <= r_n_274__13_;
      r_274__12_ <= r_n_274__12_;
      r_274__11_ <= r_n_274__11_;
      r_274__10_ <= r_n_274__10_;
      r_274__9_ <= r_n_274__9_;
      r_274__8_ <= r_n_274__8_;
      r_274__7_ <= r_n_274__7_;
      r_274__6_ <= r_n_274__6_;
      r_274__5_ <= r_n_274__5_;
      r_274__4_ <= r_n_274__4_;
      r_274__3_ <= r_n_274__3_;
      r_274__2_ <= r_n_274__2_;
      r_274__1_ <= r_n_274__1_;
      r_274__0_ <= r_n_274__0_;
    end 
    if(N3859) begin
      r_275__63_ <= r_n_275__63_;
      r_275__62_ <= r_n_275__62_;
      r_275__61_ <= r_n_275__61_;
      r_275__60_ <= r_n_275__60_;
      r_275__59_ <= r_n_275__59_;
      r_275__58_ <= r_n_275__58_;
      r_275__57_ <= r_n_275__57_;
      r_275__56_ <= r_n_275__56_;
      r_275__55_ <= r_n_275__55_;
      r_275__54_ <= r_n_275__54_;
      r_275__53_ <= r_n_275__53_;
      r_275__52_ <= r_n_275__52_;
      r_275__51_ <= r_n_275__51_;
      r_275__50_ <= r_n_275__50_;
      r_275__49_ <= r_n_275__49_;
      r_275__48_ <= r_n_275__48_;
      r_275__47_ <= r_n_275__47_;
      r_275__46_ <= r_n_275__46_;
      r_275__45_ <= r_n_275__45_;
      r_275__44_ <= r_n_275__44_;
      r_275__43_ <= r_n_275__43_;
      r_275__42_ <= r_n_275__42_;
      r_275__41_ <= r_n_275__41_;
      r_275__40_ <= r_n_275__40_;
      r_275__39_ <= r_n_275__39_;
      r_275__38_ <= r_n_275__38_;
      r_275__37_ <= r_n_275__37_;
      r_275__36_ <= r_n_275__36_;
      r_275__35_ <= r_n_275__35_;
      r_275__34_ <= r_n_275__34_;
      r_275__33_ <= r_n_275__33_;
      r_275__32_ <= r_n_275__32_;
      r_275__31_ <= r_n_275__31_;
      r_275__30_ <= r_n_275__30_;
      r_275__29_ <= r_n_275__29_;
      r_275__28_ <= r_n_275__28_;
      r_275__27_ <= r_n_275__27_;
      r_275__26_ <= r_n_275__26_;
      r_275__25_ <= r_n_275__25_;
      r_275__24_ <= r_n_275__24_;
      r_275__23_ <= r_n_275__23_;
      r_275__22_ <= r_n_275__22_;
      r_275__21_ <= r_n_275__21_;
      r_275__20_ <= r_n_275__20_;
      r_275__19_ <= r_n_275__19_;
      r_275__18_ <= r_n_275__18_;
      r_275__17_ <= r_n_275__17_;
      r_275__16_ <= r_n_275__16_;
      r_275__15_ <= r_n_275__15_;
      r_275__14_ <= r_n_275__14_;
      r_275__13_ <= r_n_275__13_;
      r_275__12_ <= r_n_275__12_;
      r_275__11_ <= r_n_275__11_;
      r_275__10_ <= r_n_275__10_;
      r_275__9_ <= r_n_275__9_;
      r_275__8_ <= r_n_275__8_;
      r_275__7_ <= r_n_275__7_;
      r_275__6_ <= r_n_275__6_;
      r_275__5_ <= r_n_275__5_;
      r_275__4_ <= r_n_275__4_;
      r_275__3_ <= r_n_275__3_;
      r_275__2_ <= r_n_275__2_;
      r_275__1_ <= r_n_275__1_;
      r_275__0_ <= r_n_275__0_;
    end 
    if(N3860) begin
      r_276__63_ <= r_n_276__63_;
      r_276__62_ <= r_n_276__62_;
      r_276__61_ <= r_n_276__61_;
      r_276__60_ <= r_n_276__60_;
      r_276__59_ <= r_n_276__59_;
      r_276__58_ <= r_n_276__58_;
      r_276__57_ <= r_n_276__57_;
      r_276__56_ <= r_n_276__56_;
      r_276__55_ <= r_n_276__55_;
      r_276__54_ <= r_n_276__54_;
      r_276__53_ <= r_n_276__53_;
      r_276__52_ <= r_n_276__52_;
      r_276__51_ <= r_n_276__51_;
      r_276__50_ <= r_n_276__50_;
      r_276__49_ <= r_n_276__49_;
      r_276__48_ <= r_n_276__48_;
      r_276__47_ <= r_n_276__47_;
      r_276__46_ <= r_n_276__46_;
      r_276__45_ <= r_n_276__45_;
      r_276__44_ <= r_n_276__44_;
      r_276__43_ <= r_n_276__43_;
      r_276__42_ <= r_n_276__42_;
      r_276__41_ <= r_n_276__41_;
      r_276__40_ <= r_n_276__40_;
      r_276__39_ <= r_n_276__39_;
      r_276__38_ <= r_n_276__38_;
      r_276__37_ <= r_n_276__37_;
      r_276__36_ <= r_n_276__36_;
      r_276__35_ <= r_n_276__35_;
      r_276__34_ <= r_n_276__34_;
      r_276__33_ <= r_n_276__33_;
      r_276__32_ <= r_n_276__32_;
      r_276__31_ <= r_n_276__31_;
      r_276__30_ <= r_n_276__30_;
      r_276__29_ <= r_n_276__29_;
      r_276__28_ <= r_n_276__28_;
      r_276__27_ <= r_n_276__27_;
      r_276__26_ <= r_n_276__26_;
      r_276__25_ <= r_n_276__25_;
      r_276__24_ <= r_n_276__24_;
      r_276__23_ <= r_n_276__23_;
      r_276__22_ <= r_n_276__22_;
      r_276__21_ <= r_n_276__21_;
      r_276__20_ <= r_n_276__20_;
      r_276__19_ <= r_n_276__19_;
      r_276__18_ <= r_n_276__18_;
      r_276__17_ <= r_n_276__17_;
      r_276__16_ <= r_n_276__16_;
      r_276__15_ <= r_n_276__15_;
      r_276__14_ <= r_n_276__14_;
      r_276__13_ <= r_n_276__13_;
      r_276__12_ <= r_n_276__12_;
      r_276__11_ <= r_n_276__11_;
      r_276__10_ <= r_n_276__10_;
      r_276__9_ <= r_n_276__9_;
      r_276__8_ <= r_n_276__8_;
      r_276__7_ <= r_n_276__7_;
      r_276__6_ <= r_n_276__6_;
      r_276__5_ <= r_n_276__5_;
      r_276__4_ <= r_n_276__4_;
      r_276__3_ <= r_n_276__3_;
      r_276__2_ <= r_n_276__2_;
      r_276__1_ <= r_n_276__1_;
      r_276__0_ <= r_n_276__0_;
    end 
    if(N3861) begin
      r_277__63_ <= r_n_277__63_;
      r_277__62_ <= r_n_277__62_;
      r_277__61_ <= r_n_277__61_;
      r_277__60_ <= r_n_277__60_;
      r_277__59_ <= r_n_277__59_;
      r_277__58_ <= r_n_277__58_;
      r_277__57_ <= r_n_277__57_;
      r_277__56_ <= r_n_277__56_;
      r_277__55_ <= r_n_277__55_;
      r_277__54_ <= r_n_277__54_;
      r_277__53_ <= r_n_277__53_;
      r_277__52_ <= r_n_277__52_;
      r_277__51_ <= r_n_277__51_;
      r_277__50_ <= r_n_277__50_;
      r_277__49_ <= r_n_277__49_;
      r_277__48_ <= r_n_277__48_;
      r_277__47_ <= r_n_277__47_;
      r_277__46_ <= r_n_277__46_;
      r_277__45_ <= r_n_277__45_;
      r_277__44_ <= r_n_277__44_;
      r_277__43_ <= r_n_277__43_;
      r_277__42_ <= r_n_277__42_;
      r_277__41_ <= r_n_277__41_;
      r_277__40_ <= r_n_277__40_;
      r_277__39_ <= r_n_277__39_;
      r_277__38_ <= r_n_277__38_;
      r_277__37_ <= r_n_277__37_;
      r_277__36_ <= r_n_277__36_;
      r_277__35_ <= r_n_277__35_;
      r_277__34_ <= r_n_277__34_;
      r_277__33_ <= r_n_277__33_;
      r_277__32_ <= r_n_277__32_;
      r_277__31_ <= r_n_277__31_;
      r_277__30_ <= r_n_277__30_;
      r_277__29_ <= r_n_277__29_;
      r_277__28_ <= r_n_277__28_;
      r_277__27_ <= r_n_277__27_;
      r_277__26_ <= r_n_277__26_;
      r_277__25_ <= r_n_277__25_;
      r_277__24_ <= r_n_277__24_;
      r_277__23_ <= r_n_277__23_;
      r_277__22_ <= r_n_277__22_;
      r_277__21_ <= r_n_277__21_;
      r_277__20_ <= r_n_277__20_;
      r_277__19_ <= r_n_277__19_;
      r_277__18_ <= r_n_277__18_;
      r_277__17_ <= r_n_277__17_;
      r_277__16_ <= r_n_277__16_;
      r_277__15_ <= r_n_277__15_;
      r_277__14_ <= r_n_277__14_;
      r_277__13_ <= r_n_277__13_;
      r_277__12_ <= r_n_277__12_;
      r_277__11_ <= r_n_277__11_;
      r_277__10_ <= r_n_277__10_;
      r_277__9_ <= r_n_277__9_;
      r_277__8_ <= r_n_277__8_;
      r_277__7_ <= r_n_277__7_;
      r_277__6_ <= r_n_277__6_;
      r_277__5_ <= r_n_277__5_;
      r_277__4_ <= r_n_277__4_;
      r_277__3_ <= r_n_277__3_;
      r_277__2_ <= r_n_277__2_;
      r_277__1_ <= r_n_277__1_;
      r_277__0_ <= r_n_277__0_;
    end 
    if(N3862) begin
      r_278__63_ <= r_n_278__63_;
      r_278__62_ <= r_n_278__62_;
      r_278__61_ <= r_n_278__61_;
      r_278__60_ <= r_n_278__60_;
      r_278__59_ <= r_n_278__59_;
      r_278__58_ <= r_n_278__58_;
      r_278__57_ <= r_n_278__57_;
      r_278__56_ <= r_n_278__56_;
      r_278__55_ <= r_n_278__55_;
      r_278__54_ <= r_n_278__54_;
      r_278__53_ <= r_n_278__53_;
      r_278__52_ <= r_n_278__52_;
      r_278__51_ <= r_n_278__51_;
      r_278__50_ <= r_n_278__50_;
      r_278__49_ <= r_n_278__49_;
      r_278__48_ <= r_n_278__48_;
      r_278__47_ <= r_n_278__47_;
      r_278__46_ <= r_n_278__46_;
      r_278__45_ <= r_n_278__45_;
      r_278__44_ <= r_n_278__44_;
      r_278__43_ <= r_n_278__43_;
      r_278__42_ <= r_n_278__42_;
      r_278__41_ <= r_n_278__41_;
      r_278__40_ <= r_n_278__40_;
      r_278__39_ <= r_n_278__39_;
      r_278__38_ <= r_n_278__38_;
      r_278__37_ <= r_n_278__37_;
      r_278__36_ <= r_n_278__36_;
      r_278__35_ <= r_n_278__35_;
      r_278__34_ <= r_n_278__34_;
      r_278__33_ <= r_n_278__33_;
      r_278__32_ <= r_n_278__32_;
      r_278__31_ <= r_n_278__31_;
      r_278__30_ <= r_n_278__30_;
      r_278__29_ <= r_n_278__29_;
      r_278__28_ <= r_n_278__28_;
      r_278__27_ <= r_n_278__27_;
      r_278__26_ <= r_n_278__26_;
      r_278__25_ <= r_n_278__25_;
      r_278__24_ <= r_n_278__24_;
      r_278__23_ <= r_n_278__23_;
      r_278__22_ <= r_n_278__22_;
      r_278__21_ <= r_n_278__21_;
      r_278__20_ <= r_n_278__20_;
      r_278__19_ <= r_n_278__19_;
      r_278__18_ <= r_n_278__18_;
      r_278__17_ <= r_n_278__17_;
      r_278__16_ <= r_n_278__16_;
      r_278__15_ <= r_n_278__15_;
      r_278__14_ <= r_n_278__14_;
      r_278__13_ <= r_n_278__13_;
      r_278__12_ <= r_n_278__12_;
      r_278__11_ <= r_n_278__11_;
      r_278__10_ <= r_n_278__10_;
      r_278__9_ <= r_n_278__9_;
      r_278__8_ <= r_n_278__8_;
      r_278__7_ <= r_n_278__7_;
      r_278__6_ <= r_n_278__6_;
      r_278__5_ <= r_n_278__5_;
      r_278__4_ <= r_n_278__4_;
      r_278__3_ <= r_n_278__3_;
      r_278__2_ <= r_n_278__2_;
      r_278__1_ <= r_n_278__1_;
      r_278__0_ <= r_n_278__0_;
    end 
    if(N3863) begin
      r_279__63_ <= r_n_279__63_;
      r_279__62_ <= r_n_279__62_;
      r_279__61_ <= r_n_279__61_;
      r_279__60_ <= r_n_279__60_;
      r_279__59_ <= r_n_279__59_;
      r_279__58_ <= r_n_279__58_;
      r_279__57_ <= r_n_279__57_;
      r_279__56_ <= r_n_279__56_;
      r_279__55_ <= r_n_279__55_;
      r_279__54_ <= r_n_279__54_;
      r_279__53_ <= r_n_279__53_;
      r_279__52_ <= r_n_279__52_;
      r_279__51_ <= r_n_279__51_;
      r_279__50_ <= r_n_279__50_;
      r_279__49_ <= r_n_279__49_;
      r_279__48_ <= r_n_279__48_;
      r_279__47_ <= r_n_279__47_;
      r_279__46_ <= r_n_279__46_;
      r_279__45_ <= r_n_279__45_;
      r_279__44_ <= r_n_279__44_;
      r_279__43_ <= r_n_279__43_;
      r_279__42_ <= r_n_279__42_;
      r_279__41_ <= r_n_279__41_;
      r_279__40_ <= r_n_279__40_;
      r_279__39_ <= r_n_279__39_;
      r_279__38_ <= r_n_279__38_;
      r_279__37_ <= r_n_279__37_;
      r_279__36_ <= r_n_279__36_;
      r_279__35_ <= r_n_279__35_;
      r_279__34_ <= r_n_279__34_;
      r_279__33_ <= r_n_279__33_;
      r_279__32_ <= r_n_279__32_;
      r_279__31_ <= r_n_279__31_;
      r_279__30_ <= r_n_279__30_;
      r_279__29_ <= r_n_279__29_;
      r_279__28_ <= r_n_279__28_;
      r_279__27_ <= r_n_279__27_;
      r_279__26_ <= r_n_279__26_;
      r_279__25_ <= r_n_279__25_;
      r_279__24_ <= r_n_279__24_;
      r_279__23_ <= r_n_279__23_;
      r_279__22_ <= r_n_279__22_;
      r_279__21_ <= r_n_279__21_;
      r_279__20_ <= r_n_279__20_;
      r_279__19_ <= r_n_279__19_;
      r_279__18_ <= r_n_279__18_;
      r_279__17_ <= r_n_279__17_;
      r_279__16_ <= r_n_279__16_;
      r_279__15_ <= r_n_279__15_;
      r_279__14_ <= r_n_279__14_;
      r_279__13_ <= r_n_279__13_;
      r_279__12_ <= r_n_279__12_;
      r_279__11_ <= r_n_279__11_;
      r_279__10_ <= r_n_279__10_;
      r_279__9_ <= r_n_279__9_;
      r_279__8_ <= r_n_279__8_;
      r_279__7_ <= r_n_279__7_;
      r_279__6_ <= r_n_279__6_;
      r_279__5_ <= r_n_279__5_;
      r_279__4_ <= r_n_279__4_;
      r_279__3_ <= r_n_279__3_;
      r_279__2_ <= r_n_279__2_;
      r_279__1_ <= r_n_279__1_;
      r_279__0_ <= r_n_279__0_;
    end 
    if(N3864) begin
      r_280__63_ <= r_n_280__63_;
      r_280__62_ <= r_n_280__62_;
      r_280__61_ <= r_n_280__61_;
      r_280__60_ <= r_n_280__60_;
      r_280__59_ <= r_n_280__59_;
      r_280__58_ <= r_n_280__58_;
      r_280__57_ <= r_n_280__57_;
      r_280__56_ <= r_n_280__56_;
      r_280__55_ <= r_n_280__55_;
      r_280__54_ <= r_n_280__54_;
      r_280__53_ <= r_n_280__53_;
      r_280__52_ <= r_n_280__52_;
      r_280__51_ <= r_n_280__51_;
      r_280__50_ <= r_n_280__50_;
      r_280__49_ <= r_n_280__49_;
      r_280__48_ <= r_n_280__48_;
      r_280__47_ <= r_n_280__47_;
      r_280__46_ <= r_n_280__46_;
      r_280__45_ <= r_n_280__45_;
      r_280__44_ <= r_n_280__44_;
      r_280__43_ <= r_n_280__43_;
      r_280__42_ <= r_n_280__42_;
      r_280__41_ <= r_n_280__41_;
      r_280__40_ <= r_n_280__40_;
      r_280__39_ <= r_n_280__39_;
      r_280__38_ <= r_n_280__38_;
      r_280__37_ <= r_n_280__37_;
      r_280__36_ <= r_n_280__36_;
      r_280__35_ <= r_n_280__35_;
      r_280__34_ <= r_n_280__34_;
      r_280__33_ <= r_n_280__33_;
      r_280__32_ <= r_n_280__32_;
      r_280__31_ <= r_n_280__31_;
      r_280__30_ <= r_n_280__30_;
      r_280__29_ <= r_n_280__29_;
      r_280__28_ <= r_n_280__28_;
      r_280__27_ <= r_n_280__27_;
      r_280__26_ <= r_n_280__26_;
      r_280__25_ <= r_n_280__25_;
      r_280__24_ <= r_n_280__24_;
      r_280__23_ <= r_n_280__23_;
      r_280__22_ <= r_n_280__22_;
      r_280__21_ <= r_n_280__21_;
      r_280__20_ <= r_n_280__20_;
      r_280__19_ <= r_n_280__19_;
      r_280__18_ <= r_n_280__18_;
      r_280__17_ <= r_n_280__17_;
      r_280__16_ <= r_n_280__16_;
      r_280__15_ <= r_n_280__15_;
      r_280__14_ <= r_n_280__14_;
      r_280__13_ <= r_n_280__13_;
      r_280__12_ <= r_n_280__12_;
      r_280__11_ <= r_n_280__11_;
      r_280__10_ <= r_n_280__10_;
      r_280__9_ <= r_n_280__9_;
      r_280__8_ <= r_n_280__8_;
      r_280__7_ <= r_n_280__7_;
      r_280__6_ <= r_n_280__6_;
      r_280__5_ <= r_n_280__5_;
      r_280__4_ <= r_n_280__4_;
      r_280__3_ <= r_n_280__3_;
      r_280__2_ <= r_n_280__2_;
      r_280__1_ <= r_n_280__1_;
      r_280__0_ <= r_n_280__0_;
    end 
    if(N3865) begin
      r_281__63_ <= r_n_281__63_;
      r_281__62_ <= r_n_281__62_;
      r_281__61_ <= r_n_281__61_;
      r_281__60_ <= r_n_281__60_;
      r_281__59_ <= r_n_281__59_;
      r_281__58_ <= r_n_281__58_;
      r_281__57_ <= r_n_281__57_;
      r_281__56_ <= r_n_281__56_;
      r_281__55_ <= r_n_281__55_;
      r_281__54_ <= r_n_281__54_;
      r_281__53_ <= r_n_281__53_;
      r_281__52_ <= r_n_281__52_;
      r_281__51_ <= r_n_281__51_;
      r_281__50_ <= r_n_281__50_;
      r_281__49_ <= r_n_281__49_;
      r_281__48_ <= r_n_281__48_;
      r_281__47_ <= r_n_281__47_;
      r_281__46_ <= r_n_281__46_;
      r_281__45_ <= r_n_281__45_;
      r_281__44_ <= r_n_281__44_;
      r_281__43_ <= r_n_281__43_;
      r_281__42_ <= r_n_281__42_;
      r_281__41_ <= r_n_281__41_;
      r_281__40_ <= r_n_281__40_;
      r_281__39_ <= r_n_281__39_;
      r_281__38_ <= r_n_281__38_;
      r_281__37_ <= r_n_281__37_;
      r_281__36_ <= r_n_281__36_;
      r_281__35_ <= r_n_281__35_;
      r_281__34_ <= r_n_281__34_;
      r_281__33_ <= r_n_281__33_;
      r_281__32_ <= r_n_281__32_;
      r_281__31_ <= r_n_281__31_;
      r_281__30_ <= r_n_281__30_;
      r_281__29_ <= r_n_281__29_;
      r_281__28_ <= r_n_281__28_;
      r_281__27_ <= r_n_281__27_;
      r_281__26_ <= r_n_281__26_;
      r_281__25_ <= r_n_281__25_;
      r_281__24_ <= r_n_281__24_;
      r_281__23_ <= r_n_281__23_;
      r_281__22_ <= r_n_281__22_;
      r_281__21_ <= r_n_281__21_;
      r_281__20_ <= r_n_281__20_;
      r_281__19_ <= r_n_281__19_;
      r_281__18_ <= r_n_281__18_;
      r_281__17_ <= r_n_281__17_;
      r_281__16_ <= r_n_281__16_;
      r_281__15_ <= r_n_281__15_;
      r_281__14_ <= r_n_281__14_;
      r_281__13_ <= r_n_281__13_;
      r_281__12_ <= r_n_281__12_;
      r_281__11_ <= r_n_281__11_;
      r_281__10_ <= r_n_281__10_;
      r_281__9_ <= r_n_281__9_;
      r_281__8_ <= r_n_281__8_;
      r_281__7_ <= r_n_281__7_;
      r_281__6_ <= r_n_281__6_;
      r_281__5_ <= r_n_281__5_;
      r_281__4_ <= r_n_281__4_;
      r_281__3_ <= r_n_281__3_;
      r_281__2_ <= r_n_281__2_;
      r_281__1_ <= r_n_281__1_;
      r_281__0_ <= r_n_281__0_;
    end 
    if(N3866) begin
      r_282__63_ <= r_n_282__63_;
      r_282__62_ <= r_n_282__62_;
      r_282__61_ <= r_n_282__61_;
      r_282__60_ <= r_n_282__60_;
      r_282__59_ <= r_n_282__59_;
      r_282__58_ <= r_n_282__58_;
      r_282__57_ <= r_n_282__57_;
      r_282__56_ <= r_n_282__56_;
      r_282__55_ <= r_n_282__55_;
      r_282__54_ <= r_n_282__54_;
      r_282__53_ <= r_n_282__53_;
      r_282__52_ <= r_n_282__52_;
      r_282__51_ <= r_n_282__51_;
      r_282__50_ <= r_n_282__50_;
      r_282__49_ <= r_n_282__49_;
      r_282__48_ <= r_n_282__48_;
      r_282__47_ <= r_n_282__47_;
      r_282__46_ <= r_n_282__46_;
      r_282__45_ <= r_n_282__45_;
      r_282__44_ <= r_n_282__44_;
      r_282__43_ <= r_n_282__43_;
      r_282__42_ <= r_n_282__42_;
      r_282__41_ <= r_n_282__41_;
      r_282__40_ <= r_n_282__40_;
      r_282__39_ <= r_n_282__39_;
      r_282__38_ <= r_n_282__38_;
      r_282__37_ <= r_n_282__37_;
      r_282__36_ <= r_n_282__36_;
      r_282__35_ <= r_n_282__35_;
      r_282__34_ <= r_n_282__34_;
      r_282__33_ <= r_n_282__33_;
      r_282__32_ <= r_n_282__32_;
      r_282__31_ <= r_n_282__31_;
      r_282__30_ <= r_n_282__30_;
      r_282__29_ <= r_n_282__29_;
      r_282__28_ <= r_n_282__28_;
      r_282__27_ <= r_n_282__27_;
      r_282__26_ <= r_n_282__26_;
      r_282__25_ <= r_n_282__25_;
      r_282__24_ <= r_n_282__24_;
      r_282__23_ <= r_n_282__23_;
      r_282__22_ <= r_n_282__22_;
      r_282__21_ <= r_n_282__21_;
      r_282__20_ <= r_n_282__20_;
      r_282__19_ <= r_n_282__19_;
      r_282__18_ <= r_n_282__18_;
      r_282__17_ <= r_n_282__17_;
      r_282__16_ <= r_n_282__16_;
      r_282__15_ <= r_n_282__15_;
      r_282__14_ <= r_n_282__14_;
      r_282__13_ <= r_n_282__13_;
      r_282__12_ <= r_n_282__12_;
      r_282__11_ <= r_n_282__11_;
      r_282__10_ <= r_n_282__10_;
      r_282__9_ <= r_n_282__9_;
      r_282__8_ <= r_n_282__8_;
      r_282__7_ <= r_n_282__7_;
      r_282__6_ <= r_n_282__6_;
      r_282__5_ <= r_n_282__5_;
      r_282__4_ <= r_n_282__4_;
      r_282__3_ <= r_n_282__3_;
      r_282__2_ <= r_n_282__2_;
      r_282__1_ <= r_n_282__1_;
      r_282__0_ <= r_n_282__0_;
    end 
    if(N3867) begin
      r_283__63_ <= r_n_283__63_;
      r_283__62_ <= r_n_283__62_;
      r_283__61_ <= r_n_283__61_;
      r_283__60_ <= r_n_283__60_;
      r_283__59_ <= r_n_283__59_;
      r_283__58_ <= r_n_283__58_;
      r_283__57_ <= r_n_283__57_;
      r_283__56_ <= r_n_283__56_;
      r_283__55_ <= r_n_283__55_;
      r_283__54_ <= r_n_283__54_;
      r_283__53_ <= r_n_283__53_;
      r_283__52_ <= r_n_283__52_;
      r_283__51_ <= r_n_283__51_;
      r_283__50_ <= r_n_283__50_;
      r_283__49_ <= r_n_283__49_;
      r_283__48_ <= r_n_283__48_;
      r_283__47_ <= r_n_283__47_;
      r_283__46_ <= r_n_283__46_;
      r_283__45_ <= r_n_283__45_;
      r_283__44_ <= r_n_283__44_;
      r_283__43_ <= r_n_283__43_;
      r_283__42_ <= r_n_283__42_;
      r_283__41_ <= r_n_283__41_;
      r_283__40_ <= r_n_283__40_;
      r_283__39_ <= r_n_283__39_;
      r_283__38_ <= r_n_283__38_;
      r_283__37_ <= r_n_283__37_;
      r_283__36_ <= r_n_283__36_;
      r_283__35_ <= r_n_283__35_;
      r_283__34_ <= r_n_283__34_;
      r_283__33_ <= r_n_283__33_;
      r_283__32_ <= r_n_283__32_;
      r_283__31_ <= r_n_283__31_;
      r_283__30_ <= r_n_283__30_;
      r_283__29_ <= r_n_283__29_;
      r_283__28_ <= r_n_283__28_;
      r_283__27_ <= r_n_283__27_;
      r_283__26_ <= r_n_283__26_;
      r_283__25_ <= r_n_283__25_;
      r_283__24_ <= r_n_283__24_;
      r_283__23_ <= r_n_283__23_;
      r_283__22_ <= r_n_283__22_;
      r_283__21_ <= r_n_283__21_;
      r_283__20_ <= r_n_283__20_;
      r_283__19_ <= r_n_283__19_;
      r_283__18_ <= r_n_283__18_;
      r_283__17_ <= r_n_283__17_;
      r_283__16_ <= r_n_283__16_;
      r_283__15_ <= r_n_283__15_;
      r_283__14_ <= r_n_283__14_;
      r_283__13_ <= r_n_283__13_;
      r_283__12_ <= r_n_283__12_;
      r_283__11_ <= r_n_283__11_;
      r_283__10_ <= r_n_283__10_;
      r_283__9_ <= r_n_283__9_;
      r_283__8_ <= r_n_283__8_;
      r_283__7_ <= r_n_283__7_;
      r_283__6_ <= r_n_283__6_;
      r_283__5_ <= r_n_283__5_;
      r_283__4_ <= r_n_283__4_;
      r_283__3_ <= r_n_283__3_;
      r_283__2_ <= r_n_283__2_;
      r_283__1_ <= r_n_283__1_;
      r_283__0_ <= r_n_283__0_;
    end 
    if(N3868) begin
      r_284__63_ <= r_n_284__63_;
      r_284__62_ <= r_n_284__62_;
      r_284__61_ <= r_n_284__61_;
      r_284__60_ <= r_n_284__60_;
      r_284__59_ <= r_n_284__59_;
      r_284__58_ <= r_n_284__58_;
      r_284__57_ <= r_n_284__57_;
      r_284__56_ <= r_n_284__56_;
      r_284__55_ <= r_n_284__55_;
      r_284__54_ <= r_n_284__54_;
      r_284__53_ <= r_n_284__53_;
      r_284__52_ <= r_n_284__52_;
      r_284__51_ <= r_n_284__51_;
      r_284__50_ <= r_n_284__50_;
      r_284__49_ <= r_n_284__49_;
      r_284__48_ <= r_n_284__48_;
      r_284__47_ <= r_n_284__47_;
      r_284__46_ <= r_n_284__46_;
      r_284__45_ <= r_n_284__45_;
      r_284__44_ <= r_n_284__44_;
      r_284__43_ <= r_n_284__43_;
      r_284__42_ <= r_n_284__42_;
      r_284__41_ <= r_n_284__41_;
      r_284__40_ <= r_n_284__40_;
      r_284__39_ <= r_n_284__39_;
      r_284__38_ <= r_n_284__38_;
      r_284__37_ <= r_n_284__37_;
      r_284__36_ <= r_n_284__36_;
      r_284__35_ <= r_n_284__35_;
      r_284__34_ <= r_n_284__34_;
      r_284__33_ <= r_n_284__33_;
      r_284__32_ <= r_n_284__32_;
      r_284__31_ <= r_n_284__31_;
      r_284__30_ <= r_n_284__30_;
      r_284__29_ <= r_n_284__29_;
      r_284__28_ <= r_n_284__28_;
      r_284__27_ <= r_n_284__27_;
      r_284__26_ <= r_n_284__26_;
      r_284__25_ <= r_n_284__25_;
      r_284__24_ <= r_n_284__24_;
      r_284__23_ <= r_n_284__23_;
      r_284__22_ <= r_n_284__22_;
      r_284__21_ <= r_n_284__21_;
      r_284__20_ <= r_n_284__20_;
      r_284__19_ <= r_n_284__19_;
      r_284__18_ <= r_n_284__18_;
      r_284__17_ <= r_n_284__17_;
      r_284__16_ <= r_n_284__16_;
      r_284__15_ <= r_n_284__15_;
      r_284__14_ <= r_n_284__14_;
      r_284__13_ <= r_n_284__13_;
      r_284__12_ <= r_n_284__12_;
      r_284__11_ <= r_n_284__11_;
      r_284__10_ <= r_n_284__10_;
      r_284__9_ <= r_n_284__9_;
      r_284__8_ <= r_n_284__8_;
      r_284__7_ <= r_n_284__7_;
      r_284__6_ <= r_n_284__6_;
      r_284__5_ <= r_n_284__5_;
      r_284__4_ <= r_n_284__4_;
      r_284__3_ <= r_n_284__3_;
      r_284__2_ <= r_n_284__2_;
      r_284__1_ <= r_n_284__1_;
      r_284__0_ <= r_n_284__0_;
    end 
    if(N3869) begin
      r_285__63_ <= r_n_285__63_;
      r_285__62_ <= r_n_285__62_;
      r_285__61_ <= r_n_285__61_;
      r_285__60_ <= r_n_285__60_;
      r_285__59_ <= r_n_285__59_;
      r_285__58_ <= r_n_285__58_;
      r_285__57_ <= r_n_285__57_;
      r_285__56_ <= r_n_285__56_;
      r_285__55_ <= r_n_285__55_;
      r_285__54_ <= r_n_285__54_;
      r_285__53_ <= r_n_285__53_;
      r_285__52_ <= r_n_285__52_;
      r_285__51_ <= r_n_285__51_;
      r_285__50_ <= r_n_285__50_;
      r_285__49_ <= r_n_285__49_;
      r_285__48_ <= r_n_285__48_;
      r_285__47_ <= r_n_285__47_;
      r_285__46_ <= r_n_285__46_;
      r_285__45_ <= r_n_285__45_;
      r_285__44_ <= r_n_285__44_;
      r_285__43_ <= r_n_285__43_;
      r_285__42_ <= r_n_285__42_;
      r_285__41_ <= r_n_285__41_;
      r_285__40_ <= r_n_285__40_;
      r_285__39_ <= r_n_285__39_;
      r_285__38_ <= r_n_285__38_;
      r_285__37_ <= r_n_285__37_;
      r_285__36_ <= r_n_285__36_;
      r_285__35_ <= r_n_285__35_;
      r_285__34_ <= r_n_285__34_;
      r_285__33_ <= r_n_285__33_;
      r_285__32_ <= r_n_285__32_;
      r_285__31_ <= r_n_285__31_;
      r_285__30_ <= r_n_285__30_;
      r_285__29_ <= r_n_285__29_;
      r_285__28_ <= r_n_285__28_;
      r_285__27_ <= r_n_285__27_;
      r_285__26_ <= r_n_285__26_;
      r_285__25_ <= r_n_285__25_;
      r_285__24_ <= r_n_285__24_;
      r_285__23_ <= r_n_285__23_;
      r_285__22_ <= r_n_285__22_;
      r_285__21_ <= r_n_285__21_;
      r_285__20_ <= r_n_285__20_;
      r_285__19_ <= r_n_285__19_;
      r_285__18_ <= r_n_285__18_;
      r_285__17_ <= r_n_285__17_;
      r_285__16_ <= r_n_285__16_;
      r_285__15_ <= r_n_285__15_;
      r_285__14_ <= r_n_285__14_;
      r_285__13_ <= r_n_285__13_;
      r_285__12_ <= r_n_285__12_;
      r_285__11_ <= r_n_285__11_;
      r_285__10_ <= r_n_285__10_;
      r_285__9_ <= r_n_285__9_;
      r_285__8_ <= r_n_285__8_;
      r_285__7_ <= r_n_285__7_;
      r_285__6_ <= r_n_285__6_;
      r_285__5_ <= r_n_285__5_;
      r_285__4_ <= r_n_285__4_;
      r_285__3_ <= r_n_285__3_;
      r_285__2_ <= r_n_285__2_;
      r_285__1_ <= r_n_285__1_;
      r_285__0_ <= r_n_285__0_;
    end 
    if(N3870) begin
      r_286__63_ <= r_n_286__63_;
      r_286__62_ <= r_n_286__62_;
      r_286__61_ <= r_n_286__61_;
      r_286__60_ <= r_n_286__60_;
      r_286__59_ <= r_n_286__59_;
      r_286__58_ <= r_n_286__58_;
      r_286__57_ <= r_n_286__57_;
      r_286__56_ <= r_n_286__56_;
      r_286__55_ <= r_n_286__55_;
      r_286__54_ <= r_n_286__54_;
      r_286__53_ <= r_n_286__53_;
      r_286__52_ <= r_n_286__52_;
      r_286__51_ <= r_n_286__51_;
      r_286__50_ <= r_n_286__50_;
      r_286__49_ <= r_n_286__49_;
      r_286__48_ <= r_n_286__48_;
      r_286__47_ <= r_n_286__47_;
      r_286__46_ <= r_n_286__46_;
      r_286__45_ <= r_n_286__45_;
      r_286__44_ <= r_n_286__44_;
      r_286__43_ <= r_n_286__43_;
      r_286__42_ <= r_n_286__42_;
      r_286__41_ <= r_n_286__41_;
      r_286__40_ <= r_n_286__40_;
      r_286__39_ <= r_n_286__39_;
      r_286__38_ <= r_n_286__38_;
      r_286__37_ <= r_n_286__37_;
      r_286__36_ <= r_n_286__36_;
      r_286__35_ <= r_n_286__35_;
      r_286__34_ <= r_n_286__34_;
      r_286__33_ <= r_n_286__33_;
      r_286__32_ <= r_n_286__32_;
      r_286__31_ <= r_n_286__31_;
      r_286__30_ <= r_n_286__30_;
      r_286__29_ <= r_n_286__29_;
      r_286__28_ <= r_n_286__28_;
      r_286__27_ <= r_n_286__27_;
      r_286__26_ <= r_n_286__26_;
      r_286__25_ <= r_n_286__25_;
      r_286__24_ <= r_n_286__24_;
      r_286__23_ <= r_n_286__23_;
      r_286__22_ <= r_n_286__22_;
      r_286__21_ <= r_n_286__21_;
      r_286__20_ <= r_n_286__20_;
      r_286__19_ <= r_n_286__19_;
      r_286__18_ <= r_n_286__18_;
      r_286__17_ <= r_n_286__17_;
      r_286__16_ <= r_n_286__16_;
      r_286__15_ <= r_n_286__15_;
      r_286__14_ <= r_n_286__14_;
      r_286__13_ <= r_n_286__13_;
      r_286__12_ <= r_n_286__12_;
      r_286__11_ <= r_n_286__11_;
      r_286__10_ <= r_n_286__10_;
      r_286__9_ <= r_n_286__9_;
      r_286__8_ <= r_n_286__8_;
      r_286__7_ <= r_n_286__7_;
      r_286__6_ <= r_n_286__6_;
      r_286__5_ <= r_n_286__5_;
      r_286__4_ <= r_n_286__4_;
      r_286__3_ <= r_n_286__3_;
      r_286__2_ <= r_n_286__2_;
      r_286__1_ <= r_n_286__1_;
      r_286__0_ <= r_n_286__0_;
    end 
    if(N3871) begin
      r_287__63_ <= r_n_287__63_;
      r_287__62_ <= r_n_287__62_;
      r_287__61_ <= r_n_287__61_;
      r_287__60_ <= r_n_287__60_;
      r_287__59_ <= r_n_287__59_;
      r_287__58_ <= r_n_287__58_;
      r_287__57_ <= r_n_287__57_;
      r_287__56_ <= r_n_287__56_;
      r_287__55_ <= r_n_287__55_;
      r_287__54_ <= r_n_287__54_;
      r_287__53_ <= r_n_287__53_;
      r_287__52_ <= r_n_287__52_;
      r_287__51_ <= r_n_287__51_;
      r_287__50_ <= r_n_287__50_;
      r_287__49_ <= r_n_287__49_;
      r_287__48_ <= r_n_287__48_;
      r_287__47_ <= r_n_287__47_;
      r_287__46_ <= r_n_287__46_;
      r_287__45_ <= r_n_287__45_;
      r_287__44_ <= r_n_287__44_;
      r_287__43_ <= r_n_287__43_;
      r_287__42_ <= r_n_287__42_;
      r_287__41_ <= r_n_287__41_;
      r_287__40_ <= r_n_287__40_;
      r_287__39_ <= r_n_287__39_;
      r_287__38_ <= r_n_287__38_;
      r_287__37_ <= r_n_287__37_;
      r_287__36_ <= r_n_287__36_;
      r_287__35_ <= r_n_287__35_;
      r_287__34_ <= r_n_287__34_;
      r_287__33_ <= r_n_287__33_;
      r_287__32_ <= r_n_287__32_;
      r_287__31_ <= r_n_287__31_;
      r_287__30_ <= r_n_287__30_;
      r_287__29_ <= r_n_287__29_;
      r_287__28_ <= r_n_287__28_;
      r_287__27_ <= r_n_287__27_;
      r_287__26_ <= r_n_287__26_;
      r_287__25_ <= r_n_287__25_;
      r_287__24_ <= r_n_287__24_;
      r_287__23_ <= r_n_287__23_;
      r_287__22_ <= r_n_287__22_;
      r_287__21_ <= r_n_287__21_;
      r_287__20_ <= r_n_287__20_;
      r_287__19_ <= r_n_287__19_;
      r_287__18_ <= r_n_287__18_;
      r_287__17_ <= r_n_287__17_;
      r_287__16_ <= r_n_287__16_;
      r_287__15_ <= r_n_287__15_;
      r_287__14_ <= r_n_287__14_;
      r_287__13_ <= r_n_287__13_;
      r_287__12_ <= r_n_287__12_;
      r_287__11_ <= r_n_287__11_;
      r_287__10_ <= r_n_287__10_;
      r_287__9_ <= r_n_287__9_;
      r_287__8_ <= r_n_287__8_;
      r_287__7_ <= r_n_287__7_;
      r_287__6_ <= r_n_287__6_;
      r_287__5_ <= r_n_287__5_;
      r_287__4_ <= r_n_287__4_;
      r_287__3_ <= r_n_287__3_;
      r_287__2_ <= r_n_287__2_;
      r_287__1_ <= r_n_287__1_;
      r_287__0_ <= r_n_287__0_;
    end 
    if(N3872) begin
      r_288__63_ <= r_n_288__63_;
      r_288__62_ <= r_n_288__62_;
      r_288__61_ <= r_n_288__61_;
      r_288__60_ <= r_n_288__60_;
      r_288__59_ <= r_n_288__59_;
      r_288__58_ <= r_n_288__58_;
      r_288__57_ <= r_n_288__57_;
      r_288__56_ <= r_n_288__56_;
      r_288__55_ <= r_n_288__55_;
      r_288__54_ <= r_n_288__54_;
      r_288__53_ <= r_n_288__53_;
      r_288__52_ <= r_n_288__52_;
      r_288__51_ <= r_n_288__51_;
      r_288__50_ <= r_n_288__50_;
      r_288__49_ <= r_n_288__49_;
      r_288__48_ <= r_n_288__48_;
      r_288__47_ <= r_n_288__47_;
      r_288__46_ <= r_n_288__46_;
      r_288__45_ <= r_n_288__45_;
      r_288__44_ <= r_n_288__44_;
      r_288__43_ <= r_n_288__43_;
      r_288__42_ <= r_n_288__42_;
      r_288__41_ <= r_n_288__41_;
      r_288__40_ <= r_n_288__40_;
      r_288__39_ <= r_n_288__39_;
      r_288__38_ <= r_n_288__38_;
      r_288__37_ <= r_n_288__37_;
      r_288__36_ <= r_n_288__36_;
      r_288__35_ <= r_n_288__35_;
      r_288__34_ <= r_n_288__34_;
      r_288__33_ <= r_n_288__33_;
      r_288__32_ <= r_n_288__32_;
      r_288__31_ <= r_n_288__31_;
      r_288__30_ <= r_n_288__30_;
      r_288__29_ <= r_n_288__29_;
      r_288__28_ <= r_n_288__28_;
      r_288__27_ <= r_n_288__27_;
      r_288__26_ <= r_n_288__26_;
      r_288__25_ <= r_n_288__25_;
      r_288__24_ <= r_n_288__24_;
      r_288__23_ <= r_n_288__23_;
      r_288__22_ <= r_n_288__22_;
      r_288__21_ <= r_n_288__21_;
      r_288__20_ <= r_n_288__20_;
      r_288__19_ <= r_n_288__19_;
      r_288__18_ <= r_n_288__18_;
      r_288__17_ <= r_n_288__17_;
      r_288__16_ <= r_n_288__16_;
      r_288__15_ <= r_n_288__15_;
      r_288__14_ <= r_n_288__14_;
      r_288__13_ <= r_n_288__13_;
      r_288__12_ <= r_n_288__12_;
      r_288__11_ <= r_n_288__11_;
      r_288__10_ <= r_n_288__10_;
      r_288__9_ <= r_n_288__9_;
      r_288__8_ <= r_n_288__8_;
      r_288__7_ <= r_n_288__7_;
      r_288__6_ <= r_n_288__6_;
      r_288__5_ <= r_n_288__5_;
      r_288__4_ <= r_n_288__4_;
      r_288__3_ <= r_n_288__3_;
      r_288__2_ <= r_n_288__2_;
      r_288__1_ <= r_n_288__1_;
      r_288__0_ <= r_n_288__0_;
    end 
    if(N3873) begin
      r_289__63_ <= r_n_289__63_;
      r_289__62_ <= r_n_289__62_;
      r_289__61_ <= r_n_289__61_;
      r_289__60_ <= r_n_289__60_;
      r_289__59_ <= r_n_289__59_;
      r_289__58_ <= r_n_289__58_;
      r_289__57_ <= r_n_289__57_;
      r_289__56_ <= r_n_289__56_;
      r_289__55_ <= r_n_289__55_;
      r_289__54_ <= r_n_289__54_;
      r_289__53_ <= r_n_289__53_;
      r_289__52_ <= r_n_289__52_;
      r_289__51_ <= r_n_289__51_;
      r_289__50_ <= r_n_289__50_;
      r_289__49_ <= r_n_289__49_;
      r_289__48_ <= r_n_289__48_;
      r_289__47_ <= r_n_289__47_;
      r_289__46_ <= r_n_289__46_;
      r_289__45_ <= r_n_289__45_;
      r_289__44_ <= r_n_289__44_;
      r_289__43_ <= r_n_289__43_;
      r_289__42_ <= r_n_289__42_;
      r_289__41_ <= r_n_289__41_;
      r_289__40_ <= r_n_289__40_;
      r_289__39_ <= r_n_289__39_;
      r_289__38_ <= r_n_289__38_;
      r_289__37_ <= r_n_289__37_;
      r_289__36_ <= r_n_289__36_;
      r_289__35_ <= r_n_289__35_;
      r_289__34_ <= r_n_289__34_;
      r_289__33_ <= r_n_289__33_;
      r_289__32_ <= r_n_289__32_;
      r_289__31_ <= r_n_289__31_;
      r_289__30_ <= r_n_289__30_;
      r_289__29_ <= r_n_289__29_;
      r_289__28_ <= r_n_289__28_;
      r_289__27_ <= r_n_289__27_;
      r_289__26_ <= r_n_289__26_;
      r_289__25_ <= r_n_289__25_;
      r_289__24_ <= r_n_289__24_;
      r_289__23_ <= r_n_289__23_;
      r_289__22_ <= r_n_289__22_;
      r_289__21_ <= r_n_289__21_;
      r_289__20_ <= r_n_289__20_;
      r_289__19_ <= r_n_289__19_;
      r_289__18_ <= r_n_289__18_;
      r_289__17_ <= r_n_289__17_;
      r_289__16_ <= r_n_289__16_;
      r_289__15_ <= r_n_289__15_;
      r_289__14_ <= r_n_289__14_;
      r_289__13_ <= r_n_289__13_;
      r_289__12_ <= r_n_289__12_;
      r_289__11_ <= r_n_289__11_;
      r_289__10_ <= r_n_289__10_;
      r_289__9_ <= r_n_289__9_;
      r_289__8_ <= r_n_289__8_;
      r_289__7_ <= r_n_289__7_;
      r_289__6_ <= r_n_289__6_;
      r_289__5_ <= r_n_289__5_;
      r_289__4_ <= r_n_289__4_;
      r_289__3_ <= r_n_289__3_;
      r_289__2_ <= r_n_289__2_;
      r_289__1_ <= r_n_289__1_;
      r_289__0_ <= r_n_289__0_;
    end 
    if(N3874) begin
      r_290__63_ <= r_n_290__63_;
      r_290__62_ <= r_n_290__62_;
      r_290__61_ <= r_n_290__61_;
      r_290__60_ <= r_n_290__60_;
      r_290__59_ <= r_n_290__59_;
      r_290__58_ <= r_n_290__58_;
      r_290__57_ <= r_n_290__57_;
      r_290__56_ <= r_n_290__56_;
      r_290__55_ <= r_n_290__55_;
      r_290__54_ <= r_n_290__54_;
      r_290__53_ <= r_n_290__53_;
      r_290__52_ <= r_n_290__52_;
      r_290__51_ <= r_n_290__51_;
      r_290__50_ <= r_n_290__50_;
      r_290__49_ <= r_n_290__49_;
      r_290__48_ <= r_n_290__48_;
      r_290__47_ <= r_n_290__47_;
      r_290__46_ <= r_n_290__46_;
      r_290__45_ <= r_n_290__45_;
      r_290__44_ <= r_n_290__44_;
      r_290__43_ <= r_n_290__43_;
      r_290__42_ <= r_n_290__42_;
      r_290__41_ <= r_n_290__41_;
      r_290__40_ <= r_n_290__40_;
      r_290__39_ <= r_n_290__39_;
      r_290__38_ <= r_n_290__38_;
      r_290__37_ <= r_n_290__37_;
      r_290__36_ <= r_n_290__36_;
      r_290__35_ <= r_n_290__35_;
      r_290__34_ <= r_n_290__34_;
      r_290__33_ <= r_n_290__33_;
      r_290__32_ <= r_n_290__32_;
      r_290__31_ <= r_n_290__31_;
      r_290__30_ <= r_n_290__30_;
      r_290__29_ <= r_n_290__29_;
      r_290__28_ <= r_n_290__28_;
      r_290__27_ <= r_n_290__27_;
      r_290__26_ <= r_n_290__26_;
      r_290__25_ <= r_n_290__25_;
      r_290__24_ <= r_n_290__24_;
      r_290__23_ <= r_n_290__23_;
      r_290__22_ <= r_n_290__22_;
      r_290__21_ <= r_n_290__21_;
      r_290__20_ <= r_n_290__20_;
      r_290__19_ <= r_n_290__19_;
      r_290__18_ <= r_n_290__18_;
      r_290__17_ <= r_n_290__17_;
      r_290__16_ <= r_n_290__16_;
      r_290__15_ <= r_n_290__15_;
      r_290__14_ <= r_n_290__14_;
      r_290__13_ <= r_n_290__13_;
      r_290__12_ <= r_n_290__12_;
      r_290__11_ <= r_n_290__11_;
      r_290__10_ <= r_n_290__10_;
      r_290__9_ <= r_n_290__9_;
      r_290__8_ <= r_n_290__8_;
      r_290__7_ <= r_n_290__7_;
      r_290__6_ <= r_n_290__6_;
      r_290__5_ <= r_n_290__5_;
      r_290__4_ <= r_n_290__4_;
      r_290__3_ <= r_n_290__3_;
      r_290__2_ <= r_n_290__2_;
      r_290__1_ <= r_n_290__1_;
      r_290__0_ <= r_n_290__0_;
    end 
    if(N3875) begin
      r_291__63_ <= r_n_291__63_;
      r_291__62_ <= r_n_291__62_;
      r_291__61_ <= r_n_291__61_;
      r_291__60_ <= r_n_291__60_;
      r_291__59_ <= r_n_291__59_;
      r_291__58_ <= r_n_291__58_;
      r_291__57_ <= r_n_291__57_;
      r_291__56_ <= r_n_291__56_;
      r_291__55_ <= r_n_291__55_;
      r_291__54_ <= r_n_291__54_;
      r_291__53_ <= r_n_291__53_;
      r_291__52_ <= r_n_291__52_;
      r_291__51_ <= r_n_291__51_;
      r_291__50_ <= r_n_291__50_;
      r_291__49_ <= r_n_291__49_;
      r_291__48_ <= r_n_291__48_;
      r_291__47_ <= r_n_291__47_;
      r_291__46_ <= r_n_291__46_;
      r_291__45_ <= r_n_291__45_;
      r_291__44_ <= r_n_291__44_;
      r_291__43_ <= r_n_291__43_;
      r_291__42_ <= r_n_291__42_;
      r_291__41_ <= r_n_291__41_;
      r_291__40_ <= r_n_291__40_;
      r_291__39_ <= r_n_291__39_;
      r_291__38_ <= r_n_291__38_;
      r_291__37_ <= r_n_291__37_;
      r_291__36_ <= r_n_291__36_;
      r_291__35_ <= r_n_291__35_;
      r_291__34_ <= r_n_291__34_;
      r_291__33_ <= r_n_291__33_;
      r_291__32_ <= r_n_291__32_;
      r_291__31_ <= r_n_291__31_;
      r_291__30_ <= r_n_291__30_;
      r_291__29_ <= r_n_291__29_;
      r_291__28_ <= r_n_291__28_;
      r_291__27_ <= r_n_291__27_;
      r_291__26_ <= r_n_291__26_;
      r_291__25_ <= r_n_291__25_;
      r_291__24_ <= r_n_291__24_;
      r_291__23_ <= r_n_291__23_;
      r_291__22_ <= r_n_291__22_;
      r_291__21_ <= r_n_291__21_;
      r_291__20_ <= r_n_291__20_;
      r_291__19_ <= r_n_291__19_;
      r_291__18_ <= r_n_291__18_;
      r_291__17_ <= r_n_291__17_;
      r_291__16_ <= r_n_291__16_;
      r_291__15_ <= r_n_291__15_;
      r_291__14_ <= r_n_291__14_;
      r_291__13_ <= r_n_291__13_;
      r_291__12_ <= r_n_291__12_;
      r_291__11_ <= r_n_291__11_;
      r_291__10_ <= r_n_291__10_;
      r_291__9_ <= r_n_291__9_;
      r_291__8_ <= r_n_291__8_;
      r_291__7_ <= r_n_291__7_;
      r_291__6_ <= r_n_291__6_;
      r_291__5_ <= r_n_291__5_;
      r_291__4_ <= r_n_291__4_;
      r_291__3_ <= r_n_291__3_;
      r_291__2_ <= r_n_291__2_;
      r_291__1_ <= r_n_291__1_;
      r_291__0_ <= r_n_291__0_;
    end 
    if(N3876) begin
      r_292__63_ <= r_n_292__63_;
      r_292__62_ <= r_n_292__62_;
      r_292__61_ <= r_n_292__61_;
      r_292__60_ <= r_n_292__60_;
      r_292__59_ <= r_n_292__59_;
      r_292__58_ <= r_n_292__58_;
      r_292__57_ <= r_n_292__57_;
      r_292__56_ <= r_n_292__56_;
      r_292__55_ <= r_n_292__55_;
      r_292__54_ <= r_n_292__54_;
      r_292__53_ <= r_n_292__53_;
      r_292__52_ <= r_n_292__52_;
      r_292__51_ <= r_n_292__51_;
      r_292__50_ <= r_n_292__50_;
      r_292__49_ <= r_n_292__49_;
      r_292__48_ <= r_n_292__48_;
      r_292__47_ <= r_n_292__47_;
      r_292__46_ <= r_n_292__46_;
      r_292__45_ <= r_n_292__45_;
      r_292__44_ <= r_n_292__44_;
      r_292__43_ <= r_n_292__43_;
      r_292__42_ <= r_n_292__42_;
      r_292__41_ <= r_n_292__41_;
      r_292__40_ <= r_n_292__40_;
      r_292__39_ <= r_n_292__39_;
      r_292__38_ <= r_n_292__38_;
      r_292__37_ <= r_n_292__37_;
      r_292__36_ <= r_n_292__36_;
      r_292__35_ <= r_n_292__35_;
      r_292__34_ <= r_n_292__34_;
      r_292__33_ <= r_n_292__33_;
      r_292__32_ <= r_n_292__32_;
      r_292__31_ <= r_n_292__31_;
      r_292__30_ <= r_n_292__30_;
      r_292__29_ <= r_n_292__29_;
      r_292__28_ <= r_n_292__28_;
      r_292__27_ <= r_n_292__27_;
      r_292__26_ <= r_n_292__26_;
      r_292__25_ <= r_n_292__25_;
      r_292__24_ <= r_n_292__24_;
      r_292__23_ <= r_n_292__23_;
      r_292__22_ <= r_n_292__22_;
      r_292__21_ <= r_n_292__21_;
      r_292__20_ <= r_n_292__20_;
      r_292__19_ <= r_n_292__19_;
      r_292__18_ <= r_n_292__18_;
      r_292__17_ <= r_n_292__17_;
      r_292__16_ <= r_n_292__16_;
      r_292__15_ <= r_n_292__15_;
      r_292__14_ <= r_n_292__14_;
      r_292__13_ <= r_n_292__13_;
      r_292__12_ <= r_n_292__12_;
      r_292__11_ <= r_n_292__11_;
      r_292__10_ <= r_n_292__10_;
      r_292__9_ <= r_n_292__9_;
      r_292__8_ <= r_n_292__8_;
      r_292__7_ <= r_n_292__7_;
      r_292__6_ <= r_n_292__6_;
      r_292__5_ <= r_n_292__5_;
      r_292__4_ <= r_n_292__4_;
      r_292__3_ <= r_n_292__3_;
      r_292__2_ <= r_n_292__2_;
      r_292__1_ <= r_n_292__1_;
      r_292__0_ <= r_n_292__0_;
    end 
    if(N3877) begin
      r_293__63_ <= r_n_293__63_;
      r_293__62_ <= r_n_293__62_;
      r_293__61_ <= r_n_293__61_;
      r_293__60_ <= r_n_293__60_;
      r_293__59_ <= r_n_293__59_;
      r_293__58_ <= r_n_293__58_;
      r_293__57_ <= r_n_293__57_;
      r_293__56_ <= r_n_293__56_;
      r_293__55_ <= r_n_293__55_;
      r_293__54_ <= r_n_293__54_;
      r_293__53_ <= r_n_293__53_;
      r_293__52_ <= r_n_293__52_;
      r_293__51_ <= r_n_293__51_;
      r_293__50_ <= r_n_293__50_;
      r_293__49_ <= r_n_293__49_;
      r_293__48_ <= r_n_293__48_;
      r_293__47_ <= r_n_293__47_;
      r_293__46_ <= r_n_293__46_;
      r_293__45_ <= r_n_293__45_;
      r_293__44_ <= r_n_293__44_;
      r_293__43_ <= r_n_293__43_;
      r_293__42_ <= r_n_293__42_;
      r_293__41_ <= r_n_293__41_;
      r_293__40_ <= r_n_293__40_;
      r_293__39_ <= r_n_293__39_;
      r_293__38_ <= r_n_293__38_;
      r_293__37_ <= r_n_293__37_;
      r_293__36_ <= r_n_293__36_;
      r_293__35_ <= r_n_293__35_;
      r_293__34_ <= r_n_293__34_;
      r_293__33_ <= r_n_293__33_;
      r_293__32_ <= r_n_293__32_;
      r_293__31_ <= r_n_293__31_;
      r_293__30_ <= r_n_293__30_;
      r_293__29_ <= r_n_293__29_;
      r_293__28_ <= r_n_293__28_;
      r_293__27_ <= r_n_293__27_;
      r_293__26_ <= r_n_293__26_;
      r_293__25_ <= r_n_293__25_;
      r_293__24_ <= r_n_293__24_;
      r_293__23_ <= r_n_293__23_;
      r_293__22_ <= r_n_293__22_;
      r_293__21_ <= r_n_293__21_;
      r_293__20_ <= r_n_293__20_;
      r_293__19_ <= r_n_293__19_;
      r_293__18_ <= r_n_293__18_;
      r_293__17_ <= r_n_293__17_;
      r_293__16_ <= r_n_293__16_;
      r_293__15_ <= r_n_293__15_;
      r_293__14_ <= r_n_293__14_;
      r_293__13_ <= r_n_293__13_;
      r_293__12_ <= r_n_293__12_;
      r_293__11_ <= r_n_293__11_;
      r_293__10_ <= r_n_293__10_;
      r_293__9_ <= r_n_293__9_;
      r_293__8_ <= r_n_293__8_;
      r_293__7_ <= r_n_293__7_;
      r_293__6_ <= r_n_293__6_;
      r_293__5_ <= r_n_293__5_;
      r_293__4_ <= r_n_293__4_;
      r_293__3_ <= r_n_293__3_;
      r_293__2_ <= r_n_293__2_;
      r_293__1_ <= r_n_293__1_;
      r_293__0_ <= r_n_293__0_;
    end 
    if(N3878) begin
      r_294__63_ <= r_n_294__63_;
      r_294__62_ <= r_n_294__62_;
      r_294__61_ <= r_n_294__61_;
      r_294__60_ <= r_n_294__60_;
      r_294__59_ <= r_n_294__59_;
      r_294__58_ <= r_n_294__58_;
      r_294__57_ <= r_n_294__57_;
      r_294__56_ <= r_n_294__56_;
      r_294__55_ <= r_n_294__55_;
      r_294__54_ <= r_n_294__54_;
      r_294__53_ <= r_n_294__53_;
      r_294__52_ <= r_n_294__52_;
      r_294__51_ <= r_n_294__51_;
      r_294__50_ <= r_n_294__50_;
      r_294__49_ <= r_n_294__49_;
      r_294__48_ <= r_n_294__48_;
      r_294__47_ <= r_n_294__47_;
      r_294__46_ <= r_n_294__46_;
      r_294__45_ <= r_n_294__45_;
      r_294__44_ <= r_n_294__44_;
      r_294__43_ <= r_n_294__43_;
      r_294__42_ <= r_n_294__42_;
      r_294__41_ <= r_n_294__41_;
      r_294__40_ <= r_n_294__40_;
      r_294__39_ <= r_n_294__39_;
      r_294__38_ <= r_n_294__38_;
      r_294__37_ <= r_n_294__37_;
      r_294__36_ <= r_n_294__36_;
      r_294__35_ <= r_n_294__35_;
      r_294__34_ <= r_n_294__34_;
      r_294__33_ <= r_n_294__33_;
      r_294__32_ <= r_n_294__32_;
      r_294__31_ <= r_n_294__31_;
      r_294__30_ <= r_n_294__30_;
      r_294__29_ <= r_n_294__29_;
      r_294__28_ <= r_n_294__28_;
      r_294__27_ <= r_n_294__27_;
      r_294__26_ <= r_n_294__26_;
      r_294__25_ <= r_n_294__25_;
      r_294__24_ <= r_n_294__24_;
      r_294__23_ <= r_n_294__23_;
      r_294__22_ <= r_n_294__22_;
      r_294__21_ <= r_n_294__21_;
      r_294__20_ <= r_n_294__20_;
      r_294__19_ <= r_n_294__19_;
      r_294__18_ <= r_n_294__18_;
      r_294__17_ <= r_n_294__17_;
      r_294__16_ <= r_n_294__16_;
      r_294__15_ <= r_n_294__15_;
      r_294__14_ <= r_n_294__14_;
      r_294__13_ <= r_n_294__13_;
      r_294__12_ <= r_n_294__12_;
      r_294__11_ <= r_n_294__11_;
      r_294__10_ <= r_n_294__10_;
      r_294__9_ <= r_n_294__9_;
      r_294__8_ <= r_n_294__8_;
      r_294__7_ <= r_n_294__7_;
      r_294__6_ <= r_n_294__6_;
      r_294__5_ <= r_n_294__5_;
      r_294__4_ <= r_n_294__4_;
      r_294__3_ <= r_n_294__3_;
      r_294__2_ <= r_n_294__2_;
      r_294__1_ <= r_n_294__1_;
      r_294__0_ <= r_n_294__0_;
    end 
    if(N3879) begin
      r_295__63_ <= r_n_295__63_;
      r_295__62_ <= r_n_295__62_;
      r_295__61_ <= r_n_295__61_;
      r_295__60_ <= r_n_295__60_;
      r_295__59_ <= r_n_295__59_;
      r_295__58_ <= r_n_295__58_;
      r_295__57_ <= r_n_295__57_;
      r_295__56_ <= r_n_295__56_;
      r_295__55_ <= r_n_295__55_;
      r_295__54_ <= r_n_295__54_;
      r_295__53_ <= r_n_295__53_;
      r_295__52_ <= r_n_295__52_;
      r_295__51_ <= r_n_295__51_;
      r_295__50_ <= r_n_295__50_;
      r_295__49_ <= r_n_295__49_;
      r_295__48_ <= r_n_295__48_;
      r_295__47_ <= r_n_295__47_;
      r_295__46_ <= r_n_295__46_;
      r_295__45_ <= r_n_295__45_;
      r_295__44_ <= r_n_295__44_;
      r_295__43_ <= r_n_295__43_;
      r_295__42_ <= r_n_295__42_;
      r_295__41_ <= r_n_295__41_;
      r_295__40_ <= r_n_295__40_;
      r_295__39_ <= r_n_295__39_;
      r_295__38_ <= r_n_295__38_;
      r_295__37_ <= r_n_295__37_;
      r_295__36_ <= r_n_295__36_;
      r_295__35_ <= r_n_295__35_;
      r_295__34_ <= r_n_295__34_;
      r_295__33_ <= r_n_295__33_;
      r_295__32_ <= r_n_295__32_;
      r_295__31_ <= r_n_295__31_;
      r_295__30_ <= r_n_295__30_;
      r_295__29_ <= r_n_295__29_;
      r_295__28_ <= r_n_295__28_;
      r_295__27_ <= r_n_295__27_;
      r_295__26_ <= r_n_295__26_;
      r_295__25_ <= r_n_295__25_;
      r_295__24_ <= r_n_295__24_;
      r_295__23_ <= r_n_295__23_;
      r_295__22_ <= r_n_295__22_;
      r_295__21_ <= r_n_295__21_;
      r_295__20_ <= r_n_295__20_;
      r_295__19_ <= r_n_295__19_;
      r_295__18_ <= r_n_295__18_;
      r_295__17_ <= r_n_295__17_;
      r_295__16_ <= r_n_295__16_;
      r_295__15_ <= r_n_295__15_;
      r_295__14_ <= r_n_295__14_;
      r_295__13_ <= r_n_295__13_;
      r_295__12_ <= r_n_295__12_;
      r_295__11_ <= r_n_295__11_;
      r_295__10_ <= r_n_295__10_;
      r_295__9_ <= r_n_295__9_;
      r_295__8_ <= r_n_295__8_;
      r_295__7_ <= r_n_295__7_;
      r_295__6_ <= r_n_295__6_;
      r_295__5_ <= r_n_295__5_;
      r_295__4_ <= r_n_295__4_;
      r_295__3_ <= r_n_295__3_;
      r_295__2_ <= r_n_295__2_;
      r_295__1_ <= r_n_295__1_;
      r_295__0_ <= r_n_295__0_;
    end 
    if(N3880) begin
      r_296__63_ <= r_n_296__63_;
      r_296__62_ <= r_n_296__62_;
      r_296__61_ <= r_n_296__61_;
      r_296__60_ <= r_n_296__60_;
      r_296__59_ <= r_n_296__59_;
      r_296__58_ <= r_n_296__58_;
      r_296__57_ <= r_n_296__57_;
      r_296__56_ <= r_n_296__56_;
      r_296__55_ <= r_n_296__55_;
      r_296__54_ <= r_n_296__54_;
      r_296__53_ <= r_n_296__53_;
      r_296__52_ <= r_n_296__52_;
      r_296__51_ <= r_n_296__51_;
      r_296__50_ <= r_n_296__50_;
      r_296__49_ <= r_n_296__49_;
      r_296__48_ <= r_n_296__48_;
      r_296__47_ <= r_n_296__47_;
      r_296__46_ <= r_n_296__46_;
      r_296__45_ <= r_n_296__45_;
      r_296__44_ <= r_n_296__44_;
      r_296__43_ <= r_n_296__43_;
      r_296__42_ <= r_n_296__42_;
      r_296__41_ <= r_n_296__41_;
      r_296__40_ <= r_n_296__40_;
      r_296__39_ <= r_n_296__39_;
      r_296__38_ <= r_n_296__38_;
      r_296__37_ <= r_n_296__37_;
      r_296__36_ <= r_n_296__36_;
      r_296__35_ <= r_n_296__35_;
      r_296__34_ <= r_n_296__34_;
      r_296__33_ <= r_n_296__33_;
      r_296__32_ <= r_n_296__32_;
      r_296__31_ <= r_n_296__31_;
      r_296__30_ <= r_n_296__30_;
      r_296__29_ <= r_n_296__29_;
      r_296__28_ <= r_n_296__28_;
      r_296__27_ <= r_n_296__27_;
      r_296__26_ <= r_n_296__26_;
      r_296__25_ <= r_n_296__25_;
      r_296__24_ <= r_n_296__24_;
      r_296__23_ <= r_n_296__23_;
      r_296__22_ <= r_n_296__22_;
      r_296__21_ <= r_n_296__21_;
      r_296__20_ <= r_n_296__20_;
      r_296__19_ <= r_n_296__19_;
      r_296__18_ <= r_n_296__18_;
      r_296__17_ <= r_n_296__17_;
      r_296__16_ <= r_n_296__16_;
      r_296__15_ <= r_n_296__15_;
      r_296__14_ <= r_n_296__14_;
      r_296__13_ <= r_n_296__13_;
      r_296__12_ <= r_n_296__12_;
      r_296__11_ <= r_n_296__11_;
      r_296__10_ <= r_n_296__10_;
      r_296__9_ <= r_n_296__9_;
      r_296__8_ <= r_n_296__8_;
      r_296__7_ <= r_n_296__7_;
      r_296__6_ <= r_n_296__6_;
      r_296__5_ <= r_n_296__5_;
      r_296__4_ <= r_n_296__4_;
      r_296__3_ <= r_n_296__3_;
      r_296__2_ <= r_n_296__2_;
      r_296__1_ <= r_n_296__1_;
      r_296__0_ <= r_n_296__0_;
    end 
    if(N3881) begin
      r_297__63_ <= r_n_297__63_;
      r_297__62_ <= r_n_297__62_;
      r_297__61_ <= r_n_297__61_;
      r_297__60_ <= r_n_297__60_;
      r_297__59_ <= r_n_297__59_;
      r_297__58_ <= r_n_297__58_;
      r_297__57_ <= r_n_297__57_;
      r_297__56_ <= r_n_297__56_;
      r_297__55_ <= r_n_297__55_;
      r_297__54_ <= r_n_297__54_;
      r_297__53_ <= r_n_297__53_;
      r_297__52_ <= r_n_297__52_;
      r_297__51_ <= r_n_297__51_;
      r_297__50_ <= r_n_297__50_;
      r_297__49_ <= r_n_297__49_;
      r_297__48_ <= r_n_297__48_;
      r_297__47_ <= r_n_297__47_;
      r_297__46_ <= r_n_297__46_;
      r_297__45_ <= r_n_297__45_;
      r_297__44_ <= r_n_297__44_;
      r_297__43_ <= r_n_297__43_;
      r_297__42_ <= r_n_297__42_;
      r_297__41_ <= r_n_297__41_;
      r_297__40_ <= r_n_297__40_;
      r_297__39_ <= r_n_297__39_;
      r_297__38_ <= r_n_297__38_;
      r_297__37_ <= r_n_297__37_;
      r_297__36_ <= r_n_297__36_;
      r_297__35_ <= r_n_297__35_;
      r_297__34_ <= r_n_297__34_;
      r_297__33_ <= r_n_297__33_;
      r_297__32_ <= r_n_297__32_;
      r_297__31_ <= r_n_297__31_;
      r_297__30_ <= r_n_297__30_;
      r_297__29_ <= r_n_297__29_;
      r_297__28_ <= r_n_297__28_;
      r_297__27_ <= r_n_297__27_;
      r_297__26_ <= r_n_297__26_;
      r_297__25_ <= r_n_297__25_;
      r_297__24_ <= r_n_297__24_;
      r_297__23_ <= r_n_297__23_;
      r_297__22_ <= r_n_297__22_;
      r_297__21_ <= r_n_297__21_;
      r_297__20_ <= r_n_297__20_;
      r_297__19_ <= r_n_297__19_;
      r_297__18_ <= r_n_297__18_;
      r_297__17_ <= r_n_297__17_;
      r_297__16_ <= r_n_297__16_;
      r_297__15_ <= r_n_297__15_;
      r_297__14_ <= r_n_297__14_;
      r_297__13_ <= r_n_297__13_;
      r_297__12_ <= r_n_297__12_;
      r_297__11_ <= r_n_297__11_;
      r_297__10_ <= r_n_297__10_;
      r_297__9_ <= r_n_297__9_;
      r_297__8_ <= r_n_297__8_;
      r_297__7_ <= r_n_297__7_;
      r_297__6_ <= r_n_297__6_;
      r_297__5_ <= r_n_297__5_;
      r_297__4_ <= r_n_297__4_;
      r_297__3_ <= r_n_297__3_;
      r_297__2_ <= r_n_297__2_;
      r_297__1_ <= r_n_297__1_;
      r_297__0_ <= r_n_297__0_;
    end 
    if(N3882) begin
      r_298__63_ <= r_n_298__63_;
      r_298__62_ <= r_n_298__62_;
      r_298__61_ <= r_n_298__61_;
      r_298__60_ <= r_n_298__60_;
      r_298__59_ <= r_n_298__59_;
      r_298__58_ <= r_n_298__58_;
      r_298__57_ <= r_n_298__57_;
      r_298__56_ <= r_n_298__56_;
      r_298__55_ <= r_n_298__55_;
      r_298__54_ <= r_n_298__54_;
      r_298__53_ <= r_n_298__53_;
      r_298__52_ <= r_n_298__52_;
      r_298__51_ <= r_n_298__51_;
      r_298__50_ <= r_n_298__50_;
      r_298__49_ <= r_n_298__49_;
      r_298__48_ <= r_n_298__48_;
      r_298__47_ <= r_n_298__47_;
      r_298__46_ <= r_n_298__46_;
      r_298__45_ <= r_n_298__45_;
      r_298__44_ <= r_n_298__44_;
      r_298__43_ <= r_n_298__43_;
      r_298__42_ <= r_n_298__42_;
      r_298__41_ <= r_n_298__41_;
      r_298__40_ <= r_n_298__40_;
      r_298__39_ <= r_n_298__39_;
      r_298__38_ <= r_n_298__38_;
      r_298__37_ <= r_n_298__37_;
      r_298__36_ <= r_n_298__36_;
      r_298__35_ <= r_n_298__35_;
      r_298__34_ <= r_n_298__34_;
      r_298__33_ <= r_n_298__33_;
      r_298__32_ <= r_n_298__32_;
      r_298__31_ <= r_n_298__31_;
      r_298__30_ <= r_n_298__30_;
      r_298__29_ <= r_n_298__29_;
      r_298__28_ <= r_n_298__28_;
      r_298__27_ <= r_n_298__27_;
      r_298__26_ <= r_n_298__26_;
      r_298__25_ <= r_n_298__25_;
      r_298__24_ <= r_n_298__24_;
      r_298__23_ <= r_n_298__23_;
      r_298__22_ <= r_n_298__22_;
      r_298__21_ <= r_n_298__21_;
      r_298__20_ <= r_n_298__20_;
      r_298__19_ <= r_n_298__19_;
      r_298__18_ <= r_n_298__18_;
      r_298__17_ <= r_n_298__17_;
      r_298__16_ <= r_n_298__16_;
      r_298__15_ <= r_n_298__15_;
      r_298__14_ <= r_n_298__14_;
      r_298__13_ <= r_n_298__13_;
      r_298__12_ <= r_n_298__12_;
      r_298__11_ <= r_n_298__11_;
      r_298__10_ <= r_n_298__10_;
      r_298__9_ <= r_n_298__9_;
      r_298__8_ <= r_n_298__8_;
      r_298__7_ <= r_n_298__7_;
      r_298__6_ <= r_n_298__6_;
      r_298__5_ <= r_n_298__5_;
      r_298__4_ <= r_n_298__4_;
      r_298__3_ <= r_n_298__3_;
      r_298__2_ <= r_n_298__2_;
      r_298__1_ <= r_n_298__1_;
      r_298__0_ <= r_n_298__0_;
    end 
    if(N3883) begin
      r_299__63_ <= r_n_299__63_;
      r_299__62_ <= r_n_299__62_;
      r_299__61_ <= r_n_299__61_;
      r_299__60_ <= r_n_299__60_;
      r_299__59_ <= r_n_299__59_;
      r_299__58_ <= r_n_299__58_;
      r_299__57_ <= r_n_299__57_;
      r_299__56_ <= r_n_299__56_;
      r_299__55_ <= r_n_299__55_;
      r_299__54_ <= r_n_299__54_;
      r_299__53_ <= r_n_299__53_;
      r_299__52_ <= r_n_299__52_;
      r_299__51_ <= r_n_299__51_;
      r_299__50_ <= r_n_299__50_;
      r_299__49_ <= r_n_299__49_;
      r_299__48_ <= r_n_299__48_;
      r_299__47_ <= r_n_299__47_;
      r_299__46_ <= r_n_299__46_;
      r_299__45_ <= r_n_299__45_;
      r_299__44_ <= r_n_299__44_;
      r_299__43_ <= r_n_299__43_;
      r_299__42_ <= r_n_299__42_;
      r_299__41_ <= r_n_299__41_;
      r_299__40_ <= r_n_299__40_;
      r_299__39_ <= r_n_299__39_;
      r_299__38_ <= r_n_299__38_;
      r_299__37_ <= r_n_299__37_;
      r_299__36_ <= r_n_299__36_;
      r_299__35_ <= r_n_299__35_;
      r_299__34_ <= r_n_299__34_;
      r_299__33_ <= r_n_299__33_;
      r_299__32_ <= r_n_299__32_;
      r_299__31_ <= r_n_299__31_;
      r_299__30_ <= r_n_299__30_;
      r_299__29_ <= r_n_299__29_;
      r_299__28_ <= r_n_299__28_;
      r_299__27_ <= r_n_299__27_;
      r_299__26_ <= r_n_299__26_;
      r_299__25_ <= r_n_299__25_;
      r_299__24_ <= r_n_299__24_;
      r_299__23_ <= r_n_299__23_;
      r_299__22_ <= r_n_299__22_;
      r_299__21_ <= r_n_299__21_;
      r_299__20_ <= r_n_299__20_;
      r_299__19_ <= r_n_299__19_;
      r_299__18_ <= r_n_299__18_;
      r_299__17_ <= r_n_299__17_;
      r_299__16_ <= r_n_299__16_;
      r_299__15_ <= r_n_299__15_;
      r_299__14_ <= r_n_299__14_;
      r_299__13_ <= r_n_299__13_;
      r_299__12_ <= r_n_299__12_;
      r_299__11_ <= r_n_299__11_;
      r_299__10_ <= r_n_299__10_;
      r_299__9_ <= r_n_299__9_;
      r_299__8_ <= r_n_299__8_;
      r_299__7_ <= r_n_299__7_;
      r_299__6_ <= r_n_299__6_;
      r_299__5_ <= r_n_299__5_;
      r_299__4_ <= r_n_299__4_;
      r_299__3_ <= r_n_299__3_;
      r_299__2_ <= r_n_299__2_;
      r_299__1_ <= r_n_299__1_;
      r_299__0_ <= r_n_299__0_;
    end 
    if(N3884) begin
      r_300__63_ <= r_n_300__63_;
      r_300__62_ <= r_n_300__62_;
      r_300__61_ <= r_n_300__61_;
      r_300__60_ <= r_n_300__60_;
      r_300__59_ <= r_n_300__59_;
      r_300__58_ <= r_n_300__58_;
      r_300__57_ <= r_n_300__57_;
      r_300__56_ <= r_n_300__56_;
      r_300__55_ <= r_n_300__55_;
      r_300__54_ <= r_n_300__54_;
      r_300__53_ <= r_n_300__53_;
      r_300__52_ <= r_n_300__52_;
      r_300__51_ <= r_n_300__51_;
      r_300__50_ <= r_n_300__50_;
      r_300__49_ <= r_n_300__49_;
      r_300__48_ <= r_n_300__48_;
      r_300__47_ <= r_n_300__47_;
      r_300__46_ <= r_n_300__46_;
      r_300__45_ <= r_n_300__45_;
      r_300__44_ <= r_n_300__44_;
      r_300__43_ <= r_n_300__43_;
      r_300__42_ <= r_n_300__42_;
      r_300__41_ <= r_n_300__41_;
      r_300__40_ <= r_n_300__40_;
      r_300__39_ <= r_n_300__39_;
      r_300__38_ <= r_n_300__38_;
      r_300__37_ <= r_n_300__37_;
      r_300__36_ <= r_n_300__36_;
      r_300__35_ <= r_n_300__35_;
      r_300__34_ <= r_n_300__34_;
      r_300__33_ <= r_n_300__33_;
      r_300__32_ <= r_n_300__32_;
      r_300__31_ <= r_n_300__31_;
      r_300__30_ <= r_n_300__30_;
      r_300__29_ <= r_n_300__29_;
      r_300__28_ <= r_n_300__28_;
      r_300__27_ <= r_n_300__27_;
      r_300__26_ <= r_n_300__26_;
      r_300__25_ <= r_n_300__25_;
      r_300__24_ <= r_n_300__24_;
      r_300__23_ <= r_n_300__23_;
      r_300__22_ <= r_n_300__22_;
      r_300__21_ <= r_n_300__21_;
      r_300__20_ <= r_n_300__20_;
      r_300__19_ <= r_n_300__19_;
      r_300__18_ <= r_n_300__18_;
      r_300__17_ <= r_n_300__17_;
      r_300__16_ <= r_n_300__16_;
      r_300__15_ <= r_n_300__15_;
      r_300__14_ <= r_n_300__14_;
      r_300__13_ <= r_n_300__13_;
      r_300__12_ <= r_n_300__12_;
      r_300__11_ <= r_n_300__11_;
      r_300__10_ <= r_n_300__10_;
      r_300__9_ <= r_n_300__9_;
      r_300__8_ <= r_n_300__8_;
      r_300__7_ <= r_n_300__7_;
      r_300__6_ <= r_n_300__6_;
      r_300__5_ <= r_n_300__5_;
      r_300__4_ <= r_n_300__4_;
      r_300__3_ <= r_n_300__3_;
      r_300__2_ <= r_n_300__2_;
      r_300__1_ <= r_n_300__1_;
      r_300__0_ <= r_n_300__0_;
    end 
    if(N3885) begin
      r_301__63_ <= r_n_301__63_;
      r_301__62_ <= r_n_301__62_;
      r_301__61_ <= r_n_301__61_;
      r_301__60_ <= r_n_301__60_;
      r_301__59_ <= r_n_301__59_;
      r_301__58_ <= r_n_301__58_;
      r_301__57_ <= r_n_301__57_;
      r_301__56_ <= r_n_301__56_;
      r_301__55_ <= r_n_301__55_;
      r_301__54_ <= r_n_301__54_;
      r_301__53_ <= r_n_301__53_;
      r_301__52_ <= r_n_301__52_;
      r_301__51_ <= r_n_301__51_;
      r_301__50_ <= r_n_301__50_;
      r_301__49_ <= r_n_301__49_;
      r_301__48_ <= r_n_301__48_;
      r_301__47_ <= r_n_301__47_;
      r_301__46_ <= r_n_301__46_;
      r_301__45_ <= r_n_301__45_;
      r_301__44_ <= r_n_301__44_;
      r_301__43_ <= r_n_301__43_;
      r_301__42_ <= r_n_301__42_;
      r_301__41_ <= r_n_301__41_;
      r_301__40_ <= r_n_301__40_;
      r_301__39_ <= r_n_301__39_;
      r_301__38_ <= r_n_301__38_;
      r_301__37_ <= r_n_301__37_;
      r_301__36_ <= r_n_301__36_;
      r_301__35_ <= r_n_301__35_;
      r_301__34_ <= r_n_301__34_;
      r_301__33_ <= r_n_301__33_;
      r_301__32_ <= r_n_301__32_;
      r_301__31_ <= r_n_301__31_;
      r_301__30_ <= r_n_301__30_;
      r_301__29_ <= r_n_301__29_;
      r_301__28_ <= r_n_301__28_;
      r_301__27_ <= r_n_301__27_;
      r_301__26_ <= r_n_301__26_;
      r_301__25_ <= r_n_301__25_;
      r_301__24_ <= r_n_301__24_;
      r_301__23_ <= r_n_301__23_;
      r_301__22_ <= r_n_301__22_;
      r_301__21_ <= r_n_301__21_;
      r_301__20_ <= r_n_301__20_;
      r_301__19_ <= r_n_301__19_;
      r_301__18_ <= r_n_301__18_;
      r_301__17_ <= r_n_301__17_;
      r_301__16_ <= r_n_301__16_;
      r_301__15_ <= r_n_301__15_;
      r_301__14_ <= r_n_301__14_;
      r_301__13_ <= r_n_301__13_;
      r_301__12_ <= r_n_301__12_;
      r_301__11_ <= r_n_301__11_;
      r_301__10_ <= r_n_301__10_;
      r_301__9_ <= r_n_301__9_;
      r_301__8_ <= r_n_301__8_;
      r_301__7_ <= r_n_301__7_;
      r_301__6_ <= r_n_301__6_;
      r_301__5_ <= r_n_301__5_;
      r_301__4_ <= r_n_301__4_;
      r_301__3_ <= r_n_301__3_;
      r_301__2_ <= r_n_301__2_;
      r_301__1_ <= r_n_301__1_;
      r_301__0_ <= r_n_301__0_;
    end 
    if(N3886) begin
      r_302__63_ <= r_n_302__63_;
      r_302__62_ <= r_n_302__62_;
      r_302__61_ <= r_n_302__61_;
      r_302__60_ <= r_n_302__60_;
      r_302__59_ <= r_n_302__59_;
      r_302__58_ <= r_n_302__58_;
      r_302__57_ <= r_n_302__57_;
      r_302__56_ <= r_n_302__56_;
      r_302__55_ <= r_n_302__55_;
      r_302__54_ <= r_n_302__54_;
      r_302__53_ <= r_n_302__53_;
      r_302__52_ <= r_n_302__52_;
      r_302__51_ <= r_n_302__51_;
      r_302__50_ <= r_n_302__50_;
      r_302__49_ <= r_n_302__49_;
      r_302__48_ <= r_n_302__48_;
      r_302__47_ <= r_n_302__47_;
      r_302__46_ <= r_n_302__46_;
      r_302__45_ <= r_n_302__45_;
      r_302__44_ <= r_n_302__44_;
      r_302__43_ <= r_n_302__43_;
      r_302__42_ <= r_n_302__42_;
      r_302__41_ <= r_n_302__41_;
      r_302__40_ <= r_n_302__40_;
      r_302__39_ <= r_n_302__39_;
      r_302__38_ <= r_n_302__38_;
      r_302__37_ <= r_n_302__37_;
      r_302__36_ <= r_n_302__36_;
      r_302__35_ <= r_n_302__35_;
      r_302__34_ <= r_n_302__34_;
      r_302__33_ <= r_n_302__33_;
      r_302__32_ <= r_n_302__32_;
      r_302__31_ <= r_n_302__31_;
      r_302__30_ <= r_n_302__30_;
      r_302__29_ <= r_n_302__29_;
      r_302__28_ <= r_n_302__28_;
      r_302__27_ <= r_n_302__27_;
      r_302__26_ <= r_n_302__26_;
      r_302__25_ <= r_n_302__25_;
      r_302__24_ <= r_n_302__24_;
      r_302__23_ <= r_n_302__23_;
      r_302__22_ <= r_n_302__22_;
      r_302__21_ <= r_n_302__21_;
      r_302__20_ <= r_n_302__20_;
      r_302__19_ <= r_n_302__19_;
      r_302__18_ <= r_n_302__18_;
      r_302__17_ <= r_n_302__17_;
      r_302__16_ <= r_n_302__16_;
      r_302__15_ <= r_n_302__15_;
      r_302__14_ <= r_n_302__14_;
      r_302__13_ <= r_n_302__13_;
      r_302__12_ <= r_n_302__12_;
      r_302__11_ <= r_n_302__11_;
      r_302__10_ <= r_n_302__10_;
      r_302__9_ <= r_n_302__9_;
      r_302__8_ <= r_n_302__8_;
      r_302__7_ <= r_n_302__7_;
      r_302__6_ <= r_n_302__6_;
      r_302__5_ <= r_n_302__5_;
      r_302__4_ <= r_n_302__4_;
      r_302__3_ <= r_n_302__3_;
      r_302__2_ <= r_n_302__2_;
      r_302__1_ <= r_n_302__1_;
      r_302__0_ <= r_n_302__0_;
    end 
    if(N3887) begin
      r_303__63_ <= r_n_303__63_;
      r_303__62_ <= r_n_303__62_;
      r_303__61_ <= r_n_303__61_;
      r_303__60_ <= r_n_303__60_;
      r_303__59_ <= r_n_303__59_;
      r_303__58_ <= r_n_303__58_;
      r_303__57_ <= r_n_303__57_;
      r_303__56_ <= r_n_303__56_;
      r_303__55_ <= r_n_303__55_;
      r_303__54_ <= r_n_303__54_;
      r_303__53_ <= r_n_303__53_;
      r_303__52_ <= r_n_303__52_;
      r_303__51_ <= r_n_303__51_;
      r_303__50_ <= r_n_303__50_;
      r_303__49_ <= r_n_303__49_;
      r_303__48_ <= r_n_303__48_;
      r_303__47_ <= r_n_303__47_;
      r_303__46_ <= r_n_303__46_;
      r_303__45_ <= r_n_303__45_;
      r_303__44_ <= r_n_303__44_;
      r_303__43_ <= r_n_303__43_;
      r_303__42_ <= r_n_303__42_;
      r_303__41_ <= r_n_303__41_;
      r_303__40_ <= r_n_303__40_;
      r_303__39_ <= r_n_303__39_;
      r_303__38_ <= r_n_303__38_;
      r_303__37_ <= r_n_303__37_;
      r_303__36_ <= r_n_303__36_;
      r_303__35_ <= r_n_303__35_;
      r_303__34_ <= r_n_303__34_;
      r_303__33_ <= r_n_303__33_;
      r_303__32_ <= r_n_303__32_;
      r_303__31_ <= r_n_303__31_;
      r_303__30_ <= r_n_303__30_;
      r_303__29_ <= r_n_303__29_;
      r_303__28_ <= r_n_303__28_;
      r_303__27_ <= r_n_303__27_;
      r_303__26_ <= r_n_303__26_;
      r_303__25_ <= r_n_303__25_;
      r_303__24_ <= r_n_303__24_;
      r_303__23_ <= r_n_303__23_;
      r_303__22_ <= r_n_303__22_;
      r_303__21_ <= r_n_303__21_;
      r_303__20_ <= r_n_303__20_;
      r_303__19_ <= r_n_303__19_;
      r_303__18_ <= r_n_303__18_;
      r_303__17_ <= r_n_303__17_;
      r_303__16_ <= r_n_303__16_;
      r_303__15_ <= r_n_303__15_;
      r_303__14_ <= r_n_303__14_;
      r_303__13_ <= r_n_303__13_;
      r_303__12_ <= r_n_303__12_;
      r_303__11_ <= r_n_303__11_;
      r_303__10_ <= r_n_303__10_;
      r_303__9_ <= r_n_303__9_;
      r_303__8_ <= r_n_303__8_;
      r_303__7_ <= r_n_303__7_;
      r_303__6_ <= r_n_303__6_;
      r_303__5_ <= r_n_303__5_;
      r_303__4_ <= r_n_303__4_;
      r_303__3_ <= r_n_303__3_;
      r_303__2_ <= r_n_303__2_;
      r_303__1_ <= r_n_303__1_;
      r_303__0_ <= r_n_303__0_;
    end 
    if(N3888) begin
      r_304__63_ <= r_n_304__63_;
      r_304__62_ <= r_n_304__62_;
      r_304__61_ <= r_n_304__61_;
      r_304__60_ <= r_n_304__60_;
      r_304__59_ <= r_n_304__59_;
      r_304__58_ <= r_n_304__58_;
      r_304__57_ <= r_n_304__57_;
      r_304__56_ <= r_n_304__56_;
      r_304__55_ <= r_n_304__55_;
      r_304__54_ <= r_n_304__54_;
      r_304__53_ <= r_n_304__53_;
      r_304__52_ <= r_n_304__52_;
      r_304__51_ <= r_n_304__51_;
      r_304__50_ <= r_n_304__50_;
      r_304__49_ <= r_n_304__49_;
      r_304__48_ <= r_n_304__48_;
      r_304__47_ <= r_n_304__47_;
      r_304__46_ <= r_n_304__46_;
      r_304__45_ <= r_n_304__45_;
      r_304__44_ <= r_n_304__44_;
      r_304__43_ <= r_n_304__43_;
      r_304__42_ <= r_n_304__42_;
      r_304__41_ <= r_n_304__41_;
      r_304__40_ <= r_n_304__40_;
      r_304__39_ <= r_n_304__39_;
      r_304__38_ <= r_n_304__38_;
      r_304__37_ <= r_n_304__37_;
      r_304__36_ <= r_n_304__36_;
      r_304__35_ <= r_n_304__35_;
      r_304__34_ <= r_n_304__34_;
      r_304__33_ <= r_n_304__33_;
      r_304__32_ <= r_n_304__32_;
      r_304__31_ <= r_n_304__31_;
      r_304__30_ <= r_n_304__30_;
      r_304__29_ <= r_n_304__29_;
      r_304__28_ <= r_n_304__28_;
      r_304__27_ <= r_n_304__27_;
      r_304__26_ <= r_n_304__26_;
      r_304__25_ <= r_n_304__25_;
      r_304__24_ <= r_n_304__24_;
      r_304__23_ <= r_n_304__23_;
      r_304__22_ <= r_n_304__22_;
      r_304__21_ <= r_n_304__21_;
      r_304__20_ <= r_n_304__20_;
      r_304__19_ <= r_n_304__19_;
      r_304__18_ <= r_n_304__18_;
      r_304__17_ <= r_n_304__17_;
      r_304__16_ <= r_n_304__16_;
      r_304__15_ <= r_n_304__15_;
      r_304__14_ <= r_n_304__14_;
      r_304__13_ <= r_n_304__13_;
      r_304__12_ <= r_n_304__12_;
      r_304__11_ <= r_n_304__11_;
      r_304__10_ <= r_n_304__10_;
      r_304__9_ <= r_n_304__9_;
      r_304__8_ <= r_n_304__8_;
      r_304__7_ <= r_n_304__7_;
      r_304__6_ <= r_n_304__6_;
      r_304__5_ <= r_n_304__5_;
      r_304__4_ <= r_n_304__4_;
      r_304__3_ <= r_n_304__3_;
      r_304__2_ <= r_n_304__2_;
      r_304__1_ <= r_n_304__1_;
      r_304__0_ <= r_n_304__0_;
    end 
    if(N3889) begin
      r_305__63_ <= r_n_305__63_;
      r_305__62_ <= r_n_305__62_;
      r_305__61_ <= r_n_305__61_;
      r_305__60_ <= r_n_305__60_;
      r_305__59_ <= r_n_305__59_;
      r_305__58_ <= r_n_305__58_;
      r_305__57_ <= r_n_305__57_;
      r_305__56_ <= r_n_305__56_;
      r_305__55_ <= r_n_305__55_;
      r_305__54_ <= r_n_305__54_;
      r_305__53_ <= r_n_305__53_;
      r_305__52_ <= r_n_305__52_;
      r_305__51_ <= r_n_305__51_;
      r_305__50_ <= r_n_305__50_;
      r_305__49_ <= r_n_305__49_;
      r_305__48_ <= r_n_305__48_;
      r_305__47_ <= r_n_305__47_;
      r_305__46_ <= r_n_305__46_;
      r_305__45_ <= r_n_305__45_;
      r_305__44_ <= r_n_305__44_;
      r_305__43_ <= r_n_305__43_;
      r_305__42_ <= r_n_305__42_;
      r_305__41_ <= r_n_305__41_;
      r_305__40_ <= r_n_305__40_;
      r_305__39_ <= r_n_305__39_;
      r_305__38_ <= r_n_305__38_;
      r_305__37_ <= r_n_305__37_;
      r_305__36_ <= r_n_305__36_;
      r_305__35_ <= r_n_305__35_;
      r_305__34_ <= r_n_305__34_;
      r_305__33_ <= r_n_305__33_;
      r_305__32_ <= r_n_305__32_;
      r_305__31_ <= r_n_305__31_;
      r_305__30_ <= r_n_305__30_;
      r_305__29_ <= r_n_305__29_;
      r_305__28_ <= r_n_305__28_;
      r_305__27_ <= r_n_305__27_;
      r_305__26_ <= r_n_305__26_;
      r_305__25_ <= r_n_305__25_;
      r_305__24_ <= r_n_305__24_;
      r_305__23_ <= r_n_305__23_;
      r_305__22_ <= r_n_305__22_;
      r_305__21_ <= r_n_305__21_;
      r_305__20_ <= r_n_305__20_;
      r_305__19_ <= r_n_305__19_;
      r_305__18_ <= r_n_305__18_;
      r_305__17_ <= r_n_305__17_;
      r_305__16_ <= r_n_305__16_;
      r_305__15_ <= r_n_305__15_;
      r_305__14_ <= r_n_305__14_;
      r_305__13_ <= r_n_305__13_;
      r_305__12_ <= r_n_305__12_;
      r_305__11_ <= r_n_305__11_;
      r_305__10_ <= r_n_305__10_;
      r_305__9_ <= r_n_305__9_;
      r_305__8_ <= r_n_305__8_;
      r_305__7_ <= r_n_305__7_;
      r_305__6_ <= r_n_305__6_;
      r_305__5_ <= r_n_305__5_;
      r_305__4_ <= r_n_305__4_;
      r_305__3_ <= r_n_305__3_;
      r_305__2_ <= r_n_305__2_;
      r_305__1_ <= r_n_305__1_;
      r_305__0_ <= r_n_305__0_;
    end 
    if(N3890) begin
      r_306__63_ <= r_n_306__63_;
      r_306__62_ <= r_n_306__62_;
      r_306__61_ <= r_n_306__61_;
      r_306__60_ <= r_n_306__60_;
      r_306__59_ <= r_n_306__59_;
      r_306__58_ <= r_n_306__58_;
      r_306__57_ <= r_n_306__57_;
      r_306__56_ <= r_n_306__56_;
      r_306__55_ <= r_n_306__55_;
      r_306__54_ <= r_n_306__54_;
      r_306__53_ <= r_n_306__53_;
      r_306__52_ <= r_n_306__52_;
      r_306__51_ <= r_n_306__51_;
      r_306__50_ <= r_n_306__50_;
      r_306__49_ <= r_n_306__49_;
      r_306__48_ <= r_n_306__48_;
      r_306__47_ <= r_n_306__47_;
      r_306__46_ <= r_n_306__46_;
      r_306__45_ <= r_n_306__45_;
      r_306__44_ <= r_n_306__44_;
      r_306__43_ <= r_n_306__43_;
      r_306__42_ <= r_n_306__42_;
      r_306__41_ <= r_n_306__41_;
      r_306__40_ <= r_n_306__40_;
      r_306__39_ <= r_n_306__39_;
      r_306__38_ <= r_n_306__38_;
      r_306__37_ <= r_n_306__37_;
      r_306__36_ <= r_n_306__36_;
      r_306__35_ <= r_n_306__35_;
      r_306__34_ <= r_n_306__34_;
      r_306__33_ <= r_n_306__33_;
      r_306__32_ <= r_n_306__32_;
      r_306__31_ <= r_n_306__31_;
      r_306__30_ <= r_n_306__30_;
      r_306__29_ <= r_n_306__29_;
      r_306__28_ <= r_n_306__28_;
      r_306__27_ <= r_n_306__27_;
      r_306__26_ <= r_n_306__26_;
      r_306__25_ <= r_n_306__25_;
      r_306__24_ <= r_n_306__24_;
      r_306__23_ <= r_n_306__23_;
      r_306__22_ <= r_n_306__22_;
      r_306__21_ <= r_n_306__21_;
      r_306__20_ <= r_n_306__20_;
      r_306__19_ <= r_n_306__19_;
      r_306__18_ <= r_n_306__18_;
      r_306__17_ <= r_n_306__17_;
      r_306__16_ <= r_n_306__16_;
      r_306__15_ <= r_n_306__15_;
      r_306__14_ <= r_n_306__14_;
      r_306__13_ <= r_n_306__13_;
      r_306__12_ <= r_n_306__12_;
      r_306__11_ <= r_n_306__11_;
      r_306__10_ <= r_n_306__10_;
      r_306__9_ <= r_n_306__9_;
      r_306__8_ <= r_n_306__8_;
      r_306__7_ <= r_n_306__7_;
      r_306__6_ <= r_n_306__6_;
      r_306__5_ <= r_n_306__5_;
      r_306__4_ <= r_n_306__4_;
      r_306__3_ <= r_n_306__3_;
      r_306__2_ <= r_n_306__2_;
      r_306__1_ <= r_n_306__1_;
      r_306__0_ <= r_n_306__0_;
    end 
    if(N3891) begin
      r_307__63_ <= r_n_307__63_;
      r_307__62_ <= r_n_307__62_;
      r_307__61_ <= r_n_307__61_;
      r_307__60_ <= r_n_307__60_;
      r_307__59_ <= r_n_307__59_;
      r_307__58_ <= r_n_307__58_;
      r_307__57_ <= r_n_307__57_;
      r_307__56_ <= r_n_307__56_;
      r_307__55_ <= r_n_307__55_;
      r_307__54_ <= r_n_307__54_;
      r_307__53_ <= r_n_307__53_;
      r_307__52_ <= r_n_307__52_;
      r_307__51_ <= r_n_307__51_;
      r_307__50_ <= r_n_307__50_;
      r_307__49_ <= r_n_307__49_;
      r_307__48_ <= r_n_307__48_;
      r_307__47_ <= r_n_307__47_;
      r_307__46_ <= r_n_307__46_;
      r_307__45_ <= r_n_307__45_;
      r_307__44_ <= r_n_307__44_;
      r_307__43_ <= r_n_307__43_;
      r_307__42_ <= r_n_307__42_;
      r_307__41_ <= r_n_307__41_;
      r_307__40_ <= r_n_307__40_;
      r_307__39_ <= r_n_307__39_;
      r_307__38_ <= r_n_307__38_;
      r_307__37_ <= r_n_307__37_;
      r_307__36_ <= r_n_307__36_;
      r_307__35_ <= r_n_307__35_;
      r_307__34_ <= r_n_307__34_;
      r_307__33_ <= r_n_307__33_;
      r_307__32_ <= r_n_307__32_;
      r_307__31_ <= r_n_307__31_;
      r_307__30_ <= r_n_307__30_;
      r_307__29_ <= r_n_307__29_;
      r_307__28_ <= r_n_307__28_;
      r_307__27_ <= r_n_307__27_;
      r_307__26_ <= r_n_307__26_;
      r_307__25_ <= r_n_307__25_;
      r_307__24_ <= r_n_307__24_;
      r_307__23_ <= r_n_307__23_;
      r_307__22_ <= r_n_307__22_;
      r_307__21_ <= r_n_307__21_;
      r_307__20_ <= r_n_307__20_;
      r_307__19_ <= r_n_307__19_;
      r_307__18_ <= r_n_307__18_;
      r_307__17_ <= r_n_307__17_;
      r_307__16_ <= r_n_307__16_;
      r_307__15_ <= r_n_307__15_;
      r_307__14_ <= r_n_307__14_;
      r_307__13_ <= r_n_307__13_;
      r_307__12_ <= r_n_307__12_;
      r_307__11_ <= r_n_307__11_;
      r_307__10_ <= r_n_307__10_;
      r_307__9_ <= r_n_307__9_;
      r_307__8_ <= r_n_307__8_;
      r_307__7_ <= r_n_307__7_;
      r_307__6_ <= r_n_307__6_;
      r_307__5_ <= r_n_307__5_;
      r_307__4_ <= r_n_307__4_;
      r_307__3_ <= r_n_307__3_;
      r_307__2_ <= r_n_307__2_;
      r_307__1_ <= r_n_307__1_;
      r_307__0_ <= r_n_307__0_;
    end 
    if(N3892) begin
      r_308__63_ <= r_n_308__63_;
      r_308__62_ <= r_n_308__62_;
      r_308__61_ <= r_n_308__61_;
      r_308__60_ <= r_n_308__60_;
      r_308__59_ <= r_n_308__59_;
      r_308__58_ <= r_n_308__58_;
      r_308__57_ <= r_n_308__57_;
      r_308__56_ <= r_n_308__56_;
      r_308__55_ <= r_n_308__55_;
      r_308__54_ <= r_n_308__54_;
      r_308__53_ <= r_n_308__53_;
      r_308__52_ <= r_n_308__52_;
      r_308__51_ <= r_n_308__51_;
      r_308__50_ <= r_n_308__50_;
      r_308__49_ <= r_n_308__49_;
      r_308__48_ <= r_n_308__48_;
      r_308__47_ <= r_n_308__47_;
      r_308__46_ <= r_n_308__46_;
      r_308__45_ <= r_n_308__45_;
      r_308__44_ <= r_n_308__44_;
      r_308__43_ <= r_n_308__43_;
      r_308__42_ <= r_n_308__42_;
      r_308__41_ <= r_n_308__41_;
      r_308__40_ <= r_n_308__40_;
      r_308__39_ <= r_n_308__39_;
      r_308__38_ <= r_n_308__38_;
      r_308__37_ <= r_n_308__37_;
      r_308__36_ <= r_n_308__36_;
      r_308__35_ <= r_n_308__35_;
      r_308__34_ <= r_n_308__34_;
      r_308__33_ <= r_n_308__33_;
      r_308__32_ <= r_n_308__32_;
      r_308__31_ <= r_n_308__31_;
      r_308__30_ <= r_n_308__30_;
      r_308__29_ <= r_n_308__29_;
      r_308__28_ <= r_n_308__28_;
      r_308__27_ <= r_n_308__27_;
      r_308__26_ <= r_n_308__26_;
      r_308__25_ <= r_n_308__25_;
      r_308__24_ <= r_n_308__24_;
      r_308__23_ <= r_n_308__23_;
      r_308__22_ <= r_n_308__22_;
      r_308__21_ <= r_n_308__21_;
      r_308__20_ <= r_n_308__20_;
      r_308__19_ <= r_n_308__19_;
      r_308__18_ <= r_n_308__18_;
      r_308__17_ <= r_n_308__17_;
      r_308__16_ <= r_n_308__16_;
      r_308__15_ <= r_n_308__15_;
      r_308__14_ <= r_n_308__14_;
      r_308__13_ <= r_n_308__13_;
      r_308__12_ <= r_n_308__12_;
      r_308__11_ <= r_n_308__11_;
      r_308__10_ <= r_n_308__10_;
      r_308__9_ <= r_n_308__9_;
      r_308__8_ <= r_n_308__8_;
      r_308__7_ <= r_n_308__7_;
      r_308__6_ <= r_n_308__6_;
      r_308__5_ <= r_n_308__5_;
      r_308__4_ <= r_n_308__4_;
      r_308__3_ <= r_n_308__3_;
      r_308__2_ <= r_n_308__2_;
      r_308__1_ <= r_n_308__1_;
      r_308__0_ <= r_n_308__0_;
    end 
    if(N3893) begin
      r_309__63_ <= r_n_309__63_;
      r_309__62_ <= r_n_309__62_;
      r_309__61_ <= r_n_309__61_;
      r_309__60_ <= r_n_309__60_;
      r_309__59_ <= r_n_309__59_;
      r_309__58_ <= r_n_309__58_;
      r_309__57_ <= r_n_309__57_;
      r_309__56_ <= r_n_309__56_;
      r_309__55_ <= r_n_309__55_;
      r_309__54_ <= r_n_309__54_;
      r_309__53_ <= r_n_309__53_;
      r_309__52_ <= r_n_309__52_;
      r_309__51_ <= r_n_309__51_;
      r_309__50_ <= r_n_309__50_;
      r_309__49_ <= r_n_309__49_;
      r_309__48_ <= r_n_309__48_;
      r_309__47_ <= r_n_309__47_;
      r_309__46_ <= r_n_309__46_;
      r_309__45_ <= r_n_309__45_;
      r_309__44_ <= r_n_309__44_;
      r_309__43_ <= r_n_309__43_;
      r_309__42_ <= r_n_309__42_;
      r_309__41_ <= r_n_309__41_;
      r_309__40_ <= r_n_309__40_;
      r_309__39_ <= r_n_309__39_;
      r_309__38_ <= r_n_309__38_;
      r_309__37_ <= r_n_309__37_;
      r_309__36_ <= r_n_309__36_;
      r_309__35_ <= r_n_309__35_;
      r_309__34_ <= r_n_309__34_;
      r_309__33_ <= r_n_309__33_;
      r_309__32_ <= r_n_309__32_;
      r_309__31_ <= r_n_309__31_;
      r_309__30_ <= r_n_309__30_;
      r_309__29_ <= r_n_309__29_;
      r_309__28_ <= r_n_309__28_;
      r_309__27_ <= r_n_309__27_;
      r_309__26_ <= r_n_309__26_;
      r_309__25_ <= r_n_309__25_;
      r_309__24_ <= r_n_309__24_;
      r_309__23_ <= r_n_309__23_;
      r_309__22_ <= r_n_309__22_;
      r_309__21_ <= r_n_309__21_;
      r_309__20_ <= r_n_309__20_;
      r_309__19_ <= r_n_309__19_;
      r_309__18_ <= r_n_309__18_;
      r_309__17_ <= r_n_309__17_;
      r_309__16_ <= r_n_309__16_;
      r_309__15_ <= r_n_309__15_;
      r_309__14_ <= r_n_309__14_;
      r_309__13_ <= r_n_309__13_;
      r_309__12_ <= r_n_309__12_;
      r_309__11_ <= r_n_309__11_;
      r_309__10_ <= r_n_309__10_;
      r_309__9_ <= r_n_309__9_;
      r_309__8_ <= r_n_309__8_;
      r_309__7_ <= r_n_309__7_;
      r_309__6_ <= r_n_309__6_;
      r_309__5_ <= r_n_309__5_;
      r_309__4_ <= r_n_309__4_;
      r_309__3_ <= r_n_309__3_;
      r_309__2_ <= r_n_309__2_;
      r_309__1_ <= r_n_309__1_;
      r_309__0_ <= r_n_309__0_;
    end 
    if(N3894) begin
      r_310__63_ <= r_n_310__63_;
      r_310__62_ <= r_n_310__62_;
      r_310__61_ <= r_n_310__61_;
      r_310__60_ <= r_n_310__60_;
      r_310__59_ <= r_n_310__59_;
      r_310__58_ <= r_n_310__58_;
      r_310__57_ <= r_n_310__57_;
      r_310__56_ <= r_n_310__56_;
      r_310__55_ <= r_n_310__55_;
      r_310__54_ <= r_n_310__54_;
      r_310__53_ <= r_n_310__53_;
      r_310__52_ <= r_n_310__52_;
      r_310__51_ <= r_n_310__51_;
      r_310__50_ <= r_n_310__50_;
      r_310__49_ <= r_n_310__49_;
      r_310__48_ <= r_n_310__48_;
      r_310__47_ <= r_n_310__47_;
      r_310__46_ <= r_n_310__46_;
      r_310__45_ <= r_n_310__45_;
      r_310__44_ <= r_n_310__44_;
      r_310__43_ <= r_n_310__43_;
      r_310__42_ <= r_n_310__42_;
      r_310__41_ <= r_n_310__41_;
      r_310__40_ <= r_n_310__40_;
      r_310__39_ <= r_n_310__39_;
      r_310__38_ <= r_n_310__38_;
      r_310__37_ <= r_n_310__37_;
      r_310__36_ <= r_n_310__36_;
      r_310__35_ <= r_n_310__35_;
      r_310__34_ <= r_n_310__34_;
      r_310__33_ <= r_n_310__33_;
      r_310__32_ <= r_n_310__32_;
      r_310__31_ <= r_n_310__31_;
      r_310__30_ <= r_n_310__30_;
      r_310__29_ <= r_n_310__29_;
      r_310__28_ <= r_n_310__28_;
      r_310__27_ <= r_n_310__27_;
      r_310__26_ <= r_n_310__26_;
      r_310__25_ <= r_n_310__25_;
      r_310__24_ <= r_n_310__24_;
      r_310__23_ <= r_n_310__23_;
      r_310__22_ <= r_n_310__22_;
      r_310__21_ <= r_n_310__21_;
      r_310__20_ <= r_n_310__20_;
      r_310__19_ <= r_n_310__19_;
      r_310__18_ <= r_n_310__18_;
      r_310__17_ <= r_n_310__17_;
      r_310__16_ <= r_n_310__16_;
      r_310__15_ <= r_n_310__15_;
      r_310__14_ <= r_n_310__14_;
      r_310__13_ <= r_n_310__13_;
      r_310__12_ <= r_n_310__12_;
      r_310__11_ <= r_n_310__11_;
      r_310__10_ <= r_n_310__10_;
      r_310__9_ <= r_n_310__9_;
      r_310__8_ <= r_n_310__8_;
      r_310__7_ <= r_n_310__7_;
      r_310__6_ <= r_n_310__6_;
      r_310__5_ <= r_n_310__5_;
      r_310__4_ <= r_n_310__4_;
      r_310__3_ <= r_n_310__3_;
      r_310__2_ <= r_n_310__2_;
      r_310__1_ <= r_n_310__1_;
      r_310__0_ <= r_n_310__0_;
    end 
    if(N3895) begin
      r_311__63_ <= r_n_311__63_;
      r_311__62_ <= r_n_311__62_;
      r_311__61_ <= r_n_311__61_;
      r_311__60_ <= r_n_311__60_;
      r_311__59_ <= r_n_311__59_;
      r_311__58_ <= r_n_311__58_;
      r_311__57_ <= r_n_311__57_;
      r_311__56_ <= r_n_311__56_;
      r_311__55_ <= r_n_311__55_;
      r_311__54_ <= r_n_311__54_;
      r_311__53_ <= r_n_311__53_;
      r_311__52_ <= r_n_311__52_;
      r_311__51_ <= r_n_311__51_;
      r_311__50_ <= r_n_311__50_;
      r_311__49_ <= r_n_311__49_;
      r_311__48_ <= r_n_311__48_;
      r_311__47_ <= r_n_311__47_;
      r_311__46_ <= r_n_311__46_;
      r_311__45_ <= r_n_311__45_;
      r_311__44_ <= r_n_311__44_;
      r_311__43_ <= r_n_311__43_;
      r_311__42_ <= r_n_311__42_;
      r_311__41_ <= r_n_311__41_;
      r_311__40_ <= r_n_311__40_;
      r_311__39_ <= r_n_311__39_;
      r_311__38_ <= r_n_311__38_;
      r_311__37_ <= r_n_311__37_;
      r_311__36_ <= r_n_311__36_;
      r_311__35_ <= r_n_311__35_;
      r_311__34_ <= r_n_311__34_;
      r_311__33_ <= r_n_311__33_;
      r_311__32_ <= r_n_311__32_;
      r_311__31_ <= r_n_311__31_;
      r_311__30_ <= r_n_311__30_;
      r_311__29_ <= r_n_311__29_;
      r_311__28_ <= r_n_311__28_;
      r_311__27_ <= r_n_311__27_;
      r_311__26_ <= r_n_311__26_;
      r_311__25_ <= r_n_311__25_;
      r_311__24_ <= r_n_311__24_;
      r_311__23_ <= r_n_311__23_;
      r_311__22_ <= r_n_311__22_;
      r_311__21_ <= r_n_311__21_;
      r_311__20_ <= r_n_311__20_;
      r_311__19_ <= r_n_311__19_;
      r_311__18_ <= r_n_311__18_;
      r_311__17_ <= r_n_311__17_;
      r_311__16_ <= r_n_311__16_;
      r_311__15_ <= r_n_311__15_;
      r_311__14_ <= r_n_311__14_;
      r_311__13_ <= r_n_311__13_;
      r_311__12_ <= r_n_311__12_;
      r_311__11_ <= r_n_311__11_;
      r_311__10_ <= r_n_311__10_;
      r_311__9_ <= r_n_311__9_;
      r_311__8_ <= r_n_311__8_;
      r_311__7_ <= r_n_311__7_;
      r_311__6_ <= r_n_311__6_;
      r_311__5_ <= r_n_311__5_;
      r_311__4_ <= r_n_311__4_;
      r_311__3_ <= r_n_311__3_;
      r_311__2_ <= r_n_311__2_;
      r_311__1_ <= r_n_311__1_;
      r_311__0_ <= r_n_311__0_;
    end 
    if(N3896) begin
      r_312__63_ <= r_n_312__63_;
      r_312__62_ <= r_n_312__62_;
      r_312__61_ <= r_n_312__61_;
      r_312__60_ <= r_n_312__60_;
      r_312__59_ <= r_n_312__59_;
      r_312__58_ <= r_n_312__58_;
      r_312__57_ <= r_n_312__57_;
      r_312__56_ <= r_n_312__56_;
      r_312__55_ <= r_n_312__55_;
      r_312__54_ <= r_n_312__54_;
      r_312__53_ <= r_n_312__53_;
      r_312__52_ <= r_n_312__52_;
      r_312__51_ <= r_n_312__51_;
      r_312__50_ <= r_n_312__50_;
      r_312__49_ <= r_n_312__49_;
      r_312__48_ <= r_n_312__48_;
      r_312__47_ <= r_n_312__47_;
      r_312__46_ <= r_n_312__46_;
      r_312__45_ <= r_n_312__45_;
      r_312__44_ <= r_n_312__44_;
      r_312__43_ <= r_n_312__43_;
      r_312__42_ <= r_n_312__42_;
      r_312__41_ <= r_n_312__41_;
      r_312__40_ <= r_n_312__40_;
      r_312__39_ <= r_n_312__39_;
      r_312__38_ <= r_n_312__38_;
      r_312__37_ <= r_n_312__37_;
      r_312__36_ <= r_n_312__36_;
      r_312__35_ <= r_n_312__35_;
      r_312__34_ <= r_n_312__34_;
      r_312__33_ <= r_n_312__33_;
      r_312__32_ <= r_n_312__32_;
      r_312__31_ <= r_n_312__31_;
      r_312__30_ <= r_n_312__30_;
      r_312__29_ <= r_n_312__29_;
      r_312__28_ <= r_n_312__28_;
      r_312__27_ <= r_n_312__27_;
      r_312__26_ <= r_n_312__26_;
      r_312__25_ <= r_n_312__25_;
      r_312__24_ <= r_n_312__24_;
      r_312__23_ <= r_n_312__23_;
      r_312__22_ <= r_n_312__22_;
      r_312__21_ <= r_n_312__21_;
      r_312__20_ <= r_n_312__20_;
      r_312__19_ <= r_n_312__19_;
      r_312__18_ <= r_n_312__18_;
      r_312__17_ <= r_n_312__17_;
      r_312__16_ <= r_n_312__16_;
      r_312__15_ <= r_n_312__15_;
      r_312__14_ <= r_n_312__14_;
      r_312__13_ <= r_n_312__13_;
      r_312__12_ <= r_n_312__12_;
      r_312__11_ <= r_n_312__11_;
      r_312__10_ <= r_n_312__10_;
      r_312__9_ <= r_n_312__9_;
      r_312__8_ <= r_n_312__8_;
      r_312__7_ <= r_n_312__7_;
      r_312__6_ <= r_n_312__6_;
      r_312__5_ <= r_n_312__5_;
      r_312__4_ <= r_n_312__4_;
      r_312__3_ <= r_n_312__3_;
      r_312__2_ <= r_n_312__2_;
      r_312__1_ <= r_n_312__1_;
      r_312__0_ <= r_n_312__0_;
    end 
    if(N3897) begin
      r_313__63_ <= r_n_313__63_;
      r_313__62_ <= r_n_313__62_;
      r_313__61_ <= r_n_313__61_;
      r_313__60_ <= r_n_313__60_;
      r_313__59_ <= r_n_313__59_;
      r_313__58_ <= r_n_313__58_;
      r_313__57_ <= r_n_313__57_;
      r_313__56_ <= r_n_313__56_;
      r_313__55_ <= r_n_313__55_;
      r_313__54_ <= r_n_313__54_;
      r_313__53_ <= r_n_313__53_;
      r_313__52_ <= r_n_313__52_;
      r_313__51_ <= r_n_313__51_;
      r_313__50_ <= r_n_313__50_;
      r_313__49_ <= r_n_313__49_;
      r_313__48_ <= r_n_313__48_;
      r_313__47_ <= r_n_313__47_;
      r_313__46_ <= r_n_313__46_;
      r_313__45_ <= r_n_313__45_;
      r_313__44_ <= r_n_313__44_;
      r_313__43_ <= r_n_313__43_;
      r_313__42_ <= r_n_313__42_;
      r_313__41_ <= r_n_313__41_;
      r_313__40_ <= r_n_313__40_;
      r_313__39_ <= r_n_313__39_;
      r_313__38_ <= r_n_313__38_;
      r_313__37_ <= r_n_313__37_;
      r_313__36_ <= r_n_313__36_;
      r_313__35_ <= r_n_313__35_;
      r_313__34_ <= r_n_313__34_;
      r_313__33_ <= r_n_313__33_;
      r_313__32_ <= r_n_313__32_;
      r_313__31_ <= r_n_313__31_;
      r_313__30_ <= r_n_313__30_;
      r_313__29_ <= r_n_313__29_;
      r_313__28_ <= r_n_313__28_;
      r_313__27_ <= r_n_313__27_;
      r_313__26_ <= r_n_313__26_;
      r_313__25_ <= r_n_313__25_;
      r_313__24_ <= r_n_313__24_;
      r_313__23_ <= r_n_313__23_;
      r_313__22_ <= r_n_313__22_;
      r_313__21_ <= r_n_313__21_;
      r_313__20_ <= r_n_313__20_;
      r_313__19_ <= r_n_313__19_;
      r_313__18_ <= r_n_313__18_;
      r_313__17_ <= r_n_313__17_;
      r_313__16_ <= r_n_313__16_;
      r_313__15_ <= r_n_313__15_;
      r_313__14_ <= r_n_313__14_;
      r_313__13_ <= r_n_313__13_;
      r_313__12_ <= r_n_313__12_;
      r_313__11_ <= r_n_313__11_;
      r_313__10_ <= r_n_313__10_;
      r_313__9_ <= r_n_313__9_;
      r_313__8_ <= r_n_313__8_;
      r_313__7_ <= r_n_313__7_;
      r_313__6_ <= r_n_313__6_;
      r_313__5_ <= r_n_313__5_;
      r_313__4_ <= r_n_313__4_;
      r_313__3_ <= r_n_313__3_;
      r_313__2_ <= r_n_313__2_;
      r_313__1_ <= r_n_313__1_;
      r_313__0_ <= r_n_313__0_;
    end 
    if(N3898) begin
      r_314__63_ <= r_n_314__63_;
      r_314__62_ <= r_n_314__62_;
      r_314__61_ <= r_n_314__61_;
      r_314__60_ <= r_n_314__60_;
      r_314__59_ <= r_n_314__59_;
      r_314__58_ <= r_n_314__58_;
      r_314__57_ <= r_n_314__57_;
      r_314__56_ <= r_n_314__56_;
      r_314__55_ <= r_n_314__55_;
      r_314__54_ <= r_n_314__54_;
      r_314__53_ <= r_n_314__53_;
      r_314__52_ <= r_n_314__52_;
      r_314__51_ <= r_n_314__51_;
      r_314__50_ <= r_n_314__50_;
      r_314__49_ <= r_n_314__49_;
      r_314__48_ <= r_n_314__48_;
      r_314__47_ <= r_n_314__47_;
      r_314__46_ <= r_n_314__46_;
      r_314__45_ <= r_n_314__45_;
      r_314__44_ <= r_n_314__44_;
      r_314__43_ <= r_n_314__43_;
      r_314__42_ <= r_n_314__42_;
      r_314__41_ <= r_n_314__41_;
      r_314__40_ <= r_n_314__40_;
      r_314__39_ <= r_n_314__39_;
      r_314__38_ <= r_n_314__38_;
      r_314__37_ <= r_n_314__37_;
      r_314__36_ <= r_n_314__36_;
      r_314__35_ <= r_n_314__35_;
      r_314__34_ <= r_n_314__34_;
      r_314__33_ <= r_n_314__33_;
      r_314__32_ <= r_n_314__32_;
      r_314__31_ <= r_n_314__31_;
      r_314__30_ <= r_n_314__30_;
      r_314__29_ <= r_n_314__29_;
      r_314__28_ <= r_n_314__28_;
      r_314__27_ <= r_n_314__27_;
      r_314__26_ <= r_n_314__26_;
      r_314__25_ <= r_n_314__25_;
      r_314__24_ <= r_n_314__24_;
      r_314__23_ <= r_n_314__23_;
      r_314__22_ <= r_n_314__22_;
      r_314__21_ <= r_n_314__21_;
      r_314__20_ <= r_n_314__20_;
      r_314__19_ <= r_n_314__19_;
      r_314__18_ <= r_n_314__18_;
      r_314__17_ <= r_n_314__17_;
      r_314__16_ <= r_n_314__16_;
      r_314__15_ <= r_n_314__15_;
      r_314__14_ <= r_n_314__14_;
      r_314__13_ <= r_n_314__13_;
      r_314__12_ <= r_n_314__12_;
      r_314__11_ <= r_n_314__11_;
      r_314__10_ <= r_n_314__10_;
      r_314__9_ <= r_n_314__9_;
      r_314__8_ <= r_n_314__8_;
      r_314__7_ <= r_n_314__7_;
      r_314__6_ <= r_n_314__6_;
      r_314__5_ <= r_n_314__5_;
      r_314__4_ <= r_n_314__4_;
      r_314__3_ <= r_n_314__3_;
      r_314__2_ <= r_n_314__2_;
      r_314__1_ <= r_n_314__1_;
      r_314__0_ <= r_n_314__0_;
    end 
    if(N3899) begin
      r_315__63_ <= r_n_315__63_;
      r_315__62_ <= r_n_315__62_;
      r_315__61_ <= r_n_315__61_;
      r_315__60_ <= r_n_315__60_;
      r_315__59_ <= r_n_315__59_;
      r_315__58_ <= r_n_315__58_;
      r_315__57_ <= r_n_315__57_;
      r_315__56_ <= r_n_315__56_;
      r_315__55_ <= r_n_315__55_;
      r_315__54_ <= r_n_315__54_;
      r_315__53_ <= r_n_315__53_;
      r_315__52_ <= r_n_315__52_;
      r_315__51_ <= r_n_315__51_;
      r_315__50_ <= r_n_315__50_;
      r_315__49_ <= r_n_315__49_;
      r_315__48_ <= r_n_315__48_;
      r_315__47_ <= r_n_315__47_;
      r_315__46_ <= r_n_315__46_;
      r_315__45_ <= r_n_315__45_;
      r_315__44_ <= r_n_315__44_;
      r_315__43_ <= r_n_315__43_;
      r_315__42_ <= r_n_315__42_;
      r_315__41_ <= r_n_315__41_;
      r_315__40_ <= r_n_315__40_;
      r_315__39_ <= r_n_315__39_;
      r_315__38_ <= r_n_315__38_;
      r_315__37_ <= r_n_315__37_;
      r_315__36_ <= r_n_315__36_;
      r_315__35_ <= r_n_315__35_;
      r_315__34_ <= r_n_315__34_;
      r_315__33_ <= r_n_315__33_;
      r_315__32_ <= r_n_315__32_;
      r_315__31_ <= r_n_315__31_;
      r_315__30_ <= r_n_315__30_;
      r_315__29_ <= r_n_315__29_;
      r_315__28_ <= r_n_315__28_;
      r_315__27_ <= r_n_315__27_;
      r_315__26_ <= r_n_315__26_;
      r_315__25_ <= r_n_315__25_;
      r_315__24_ <= r_n_315__24_;
      r_315__23_ <= r_n_315__23_;
      r_315__22_ <= r_n_315__22_;
      r_315__21_ <= r_n_315__21_;
      r_315__20_ <= r_n_315__20_;
      r_315__19_ <= r_n_315__19_;
      r_315__18_ <= r_n_315__18_;
      r_315__17_ <= r_n_315__17_;
      r_315__16_ <= r_n_315__16_;
      r_315__15_ <= r_n_315__15_;
      r_315__14_ <= r_n_315__14_;
      r_315__13_ <= r_n_315__13_;
      r_315__12_ <= r_n_315__12_;
      r_315__11_ <= r_n_315__11_;
      r_315__10_ <= r_n_315__10_;
      r_315__9_ <= r_n_315__9_;
      r_315__8_ <= r_n_315__8_;
      r_315__7_ <= r_n_315__7_;
      r_315__6_ <= r_n_315__6_;
      r_315__5_ <= r_n_315__5_;
      r_315__4_ <= r_n_315__4_;
      r_315__3_ <= r_n_315__3_;
      r_315__2_ <= r_n_315__2_;
      r_315__1_ <= r_n_315__1_;
      r_315__0_ <= r_n_315__0_;
    end 
    if(N3900) begin
      r_316__63_ <= r_n_316__63_;
      r_316__62_ <= r_n_316__62_;
      r_316__61_ <= r_n_316__61_;
      r_316__60_ <= r_n_316__60_;
      r_316__59_ <= r_n_316__59_;
      r_316__58_ <= r_n_316__58_;
      r_316__57_ <= r_n_316__57_;
      r_316__56_ <= r_n_316__56_;
      r_316__55_ <= r_n_316__55_;
      r_316__54_ <= r_n_316__54_;
      r_316__53_ <= r_n_316__53_;
      r_316__52_ <= r_n_316__52_;
      r_316__51_ <= r_n_316__51_;
      r_316__50_ <= r_n_316__50_;
      r_316__49_ <= r_n_316__49_;
      r_316__48_ <= r_n_316__48_;
      r_316__47_ <= r_n_316__47_;
      r_316__46_ <= r_n_316__46_;
      r_316__45_ <= r_n_316__45_;
      r_316__44_ <= r_n_316__44_;
      r_316__43_ <= r_n_316__43_;
      r_316__42_ <= r_n_316__42_;
      r_316__41_ <= r_n_316__41_;
      r_316__40_ <= r_n_316__40_;
      r_316__39_ <= r_n_316__39_;
      r_316__38_ <= r_n_316__38_;
      r_316__37_ <= r_n_316__37_;
      r_316__36_ <= r_n_316__36_;
      r_316__35_ <= r_n_316__35_;
      r_316__34_ <= r_n_316__34_;
      r_316__33_ <= r_n_316__33_;
      r_316__32_ <= r_n_316__32_;
      r_316__31_ <= r_n_316__31_;
      r_316__30_ <= r_n_316__30_;
      r_316__29_ <= r_n_316__29_;
      r_316__28_ <= r_n_316__28_;
      r_316__27_ <= r_n_316__27_;
      r_316__26_ <= r_n_316__26_;
      r_316__25_ <= r_n_316__25_;
      r_316__24_ <= r_n_316__24_;
      r_316__23_ <= r_n_316__23_;
      r_316__22_ <= r_n_316__22_;
      r_316__21_ <= r_n_316__21_;
      r_316__20_ <= r_n_316__20_;
      r_316__19_ <= r_n_316__19_;
      r_316__18_ <= r_n_316__18_;
      r_316__17_ <= r_n_316__17_;
      r_316__16_ <= r_n_316__16_;
      r_316__15_ <= r_n_316__15_;
      r_316__14_ <= r_n_316__14_;
      r_316__13_ <= r_n_316__13_;
      r_316__12_ <= r_n_316__12_;
      r_316__11_ <= r_n_316__11_;
      r_316__10_ <= r_n_316__10_;
      r_316__9_ <= r_n_316__9_;
      r_316__8_ <= r_n_316__8_;
      r_316__7_ <= r_n_316__7_;
      r_316__6_ <= r_n_316__6_;
      r_316__5_ <= r_n_316__5_;
      r_316__4_ <= r_n_316__4_;
      r_316__3_ <= r_n_316__3_;
      r_316__2_ <= r_n_316__2_;
      r_316__1_ <= r_n_316__1_;
      r_316__0_ <= r_n_316__0_;
    end 
    if(N3901) begin
      r_317__63_ <= r_n_317__63_;
      r_317__62_ <= r_n_317__62_;
      r_317__61_ <= r_n_317__61_;
      r_317__60_ <= r_n_317__60_;
      r_317__59_ <= r_n_317__59_;
      r_317__58_ <= r_n_317__58_;
      r_317__57_ <= r_n_317__57_;
      r_317__56_ <= r_n_317__56_;
      r_317__55_ <= r_n_317__55_;
      r_317__54_ <= r_n_317__54_;
      r_317__53_ <= r_n_317__53_;
      r_317__52_ <= r_n_317__52_;
      r_317__51_ <= r_n_317__51_;
      r_317__50_ <= r_n_317__50_;
      r_317__49_ <= r_n_317__49_;
      r_317__48_ <= r_n_317__48_;
      r_317__47_ <= r_n_317__47_;
      r_317__46_ <= r_n_317__46_;
      r_317__45_ <= r_n_317__45_;
      r_317__44_ <= r_n_317__44_;
      r_317__43_ <= r_n_317__43_;
      r_317__42_ <= r_n_317__42_;
      r_317__41_ <= r_n_317__41_;
      r_317__40_ <= r_n_317__40_;
      r_317__39_ <= r_n_317__39_;
      r_317__38_ <= r_n_317__38_;
      r_317__37_ <= r_n_317__37_;
      r_317__36_ <= r_n_317__36_;
      r_317__35_ <= r_n_317__35_;
      r_317__34_ <= r_n_317__34_;
      r_317__33_ <= r_n_317__33_;
      r_317__32_ <= r_n_317__32_;
      r_317__31_ <= r_n_317__31_;
      r_317__30_ <= r_n_317__30_;
      r_317__29_ <= r_n_317__29_;
      r_317__28_ <= r_n_317__28_;
      r_317__27_ <= r_n_317__27_;
      r_317__26_ <= r_n_317__26_;
      r_317__25_ <= r_n_317__25_;
      r_317__24_ <= r_n_317__24_;
      r_317__23_ <= r_n_317__23_;
      r_317__22_ <= r_n_317__22_;
      r_317__21_ <= r_n_317__21_;
      r_317__20_ <= r_n_317__20_;
      r_317__19_ <= r_n_317__19_;
      r_317__18_ <= r_n_317__18_;
      r_317__17_ <= r_n_317__17_;
      r_317__16_ <= r_n_317__16_;
      r_317__15_ <= r_n_317__15_;
      r_317__14_ <= r_n_317__14_;
      r_317__13_ <= r_n_317__13_;
      r_317__12_ <= r_n_317__12_;
      r_317__11_ <= r_n_317__11_;
      r_317__10_ <= r_n_317__10_;
      r_317__9_ <= r_n_317__9_;
      r_317__8_ <= r_n_317__8_;
      r_317__7_ <= r_n_317__7_;
      r_317__6_ <= r_n_317__6_;
      r_317__5_ <= r_n_317__5_;
      r_317__4_ <= r_n_317__4_;
      r_317__3_ <= r_n_317__3_;
      r_317__2_ <= r_n_317__2_;
      r_317__1_ <= r_n_317__1_;
      r_317__0_ <= r_n_317__0_;
    end 
    if(N3902) begin
      r_318__63_ <= r_n_318__63_;
      r_318__62_ <= r_n_318__62_;
      r_318__61_ <= r_n_318__61_;
      r_318__60_ <= r_n_318__60_;
      r_318__59_ <= r_n_318__59_;
      r_318__58_ <= r_n_318__58_;
      r_318__57_ <= r_n_318__57_;
      r_318__56_ <= r_n_318__56_;
      r_318__55_ <= r_n_318__55_;
      r_318__54_ <= r_n_318__54_;
      r_318__53_ <= r_n_318__53_;
      r_318__52_ <= r_n_318__52_;
      r_318__51_ <= r_n_318__51_;
      r_318__50_ <= r_n_318__50_;
      r_318__49_ <= r_n_318__49_;
      r_318__48_ <= r_n_318__48_;
      r_318__47_ <= r_n_318__47_;
      r_318__46_ <= r_n_318__46_;
      r_318__45_ <= r_n_318__45_;
      r_318__44_ <= r_n_318__44_;
      r_318__43_ <= r_n_318__43_;
      r_318__42_ <= r_n_318__42_;
      r_318__41_ <= r_n_318__41_;
      r_318__40_ <= r_n_318__40_;
      r_318__39_ <= r_n_318__39_;
      r_318__38_ <= r_n_318__38_;
      r_318__37_ <= r_n_318__37_;
      r_318__36_ <= r_n_318__36_;
      r_318__35_ <= r_n_318__35_;
      r_318__34_ <= r_n_318__34_;
      r_318__33_ <= r_n_318__33_;
      r_318__32_ <= r_n_318__32_;
      r_318__31_ <= r_n_318__31_;
      r_318__30_ <= r_n_318__30_;
      r_318__29_ <= r_n_318__29_;
      r_318__28_ <= r_n_318__28_;
      r_318__27_ <= r_n_318__27_;
      r_318__26_ <= r_n_318__26_;
      r_318__25_ <= r_n_318__25_;
      r_318__24_ <= r_n_318__24_;
      r_318__23_ <= r_n_318__23_;
      r_318__22_ <= r_n_318__22_;
      r_318__21_ <= r_n_318__21_;
      r_318__20_ <= r_n_318__20_;
      r_318__19_ <= r_n_318__19_;
      r_318__18_ <= r_n_318__18_;
      r_318__17_ <= r_n_318__17_;
      r_318__16_ <= r_n_318__16_;
      r_318__15_ <= r_n_318__15_;
      r_318__14_ <= r_n_318__14_;
      r_318__13_ <= r_n_318__13_;
      r_318__12_ <= r_n_318__12_;
      r_318__11_ <= r_n_318__11_;
      r_318__10_ <= r_n_318__10_;
      r_318__9_ <= r_n_318__9_;
      r_318__8_ <= r_n_318__8_;
      r_318__7_ <= r_n_318__7_;
      r_318__6_ <= r_n_318__6_;
      r_318__5_ <= r_n_318__5_;
      r_318__4_ <= r_n_318__4_;
      r_318__3_ <= r_n_318__3_;
      r_318__2_ <= r_n_318__2_;
      r_318__1_ <= r_n_318__1_;
      r_318__0_ <= r_n_318__0_;
    end 
    if(N3903) begin
      r_319__63_ <= r_n_319__63_;
      r_319__62_ <= r_n_319__62_;
      r_319__61_ <= r_n_319__61_;
      r_319__60_ <= r_n_319__60_;
      r_319__59_ <= r_n_319__59_;
      r_319__58_ <= r_n_319__58_;
      r_319__57_ <= r_n_319__57_;
      r_319__56_ <= r_n_319__56_;
      r_319__55_ <= r_n_319__55_;
      r_319__54_ <= r_n_319__54_;
      r_319__53_ <= r_n_319__53_;
      r_319__52_ <= r_n_319__52_;
      r_319__51_ <= r_n_319__51_;
      r_319__50_ <= r_n_319__50_;
      r_319__49_ <= r_n_319__49_;
      r_319__48_ <= r_n_319__48_;
      r_319__47_ <= r_n_319__47_;
      r_319__46_ <= r_n_319__46_;
      r_319__45_ <= r_n_319__45_;
      r_319__44_ <= r_n_319__44_;
      r_319__43_ <= r_n_319__43_;
      r_319__42_ <= r_n_319__42_;
      r_319__41_ <= r_n_319__41_;
      r_319__40_ <= r_n_319__40_;
      r_319__39_ <= r_n_319__39_;
      r_319__38_ <= r_n_319__38_;
      r_319__37_ <= r_n_319__37_;
      r_319__36_ <= r_n_319__36_;
      r_319__35_ <= r_n_319__35_;
      r_319__34_ <= r_n_319__34_;
      r_319__33_ <= r_n_319__33_;
      r_319__32_ <= r_n_319__32_;
      r_319__31_ <= r_n_319__31_;
      r_319__30_ <= r_n_319__30_;
      r_319__29_ <= r_n_319__29_;
      r_319__28_ <= r_n_319__28_;
      r_319__27_ <= r_n_319__27_;
      r_319__26_ <= r_n_319__26_;
      r_319__25_ <= r_n_319__25_;
      r_319__24_ <= r_n_319__24_;
      r_319__23_ <= r_n_319__23_;
      r_319__22_ <= r_n_319__22_;
      r_319__21_ <= r_n_319__21_;
      r_319__20_ <= r_n_319__20_;
      r_319__19_ <= r_n_319__19_;
      r_319__18_ <= r_n_319__18_;
      r_319__17_ <= r_n_319__17_;
      r_319__16_ <= r_n_319__16_;
      r_319__15_ <= r_n_319__15_;
      r_319__14_ <= r_n_319__14_;
      r_319__13_ <= r_n_319__13_;
      r_319__12_ <= r_n_319__12_;
      r_319__11_ <= r_n_319__11_;
      r_319__10_ <= r_n_319__10_;
      r_319__9_ <= r_n_319__9_;
      r_319__8_ <= r_n_319__8_;
      r_319__7_ <= r_n_319__7_;
      r_319__6_ <= r_n_319__6_;
      r_319__5_ <= r_n_319__5_;
      r_319__4_ <= r_n_319__4_;
      r_319__3_ <= r_n_319__3_;
      r_319__2_ <= r_n_319__2_;
      r_319__1_ <= r_n_319__1_;
      r_319__0_ <= r_n_319__0_;
    end 
    if(N3904) begin
      r_320__63_ <= r_n_320__63_;
      r_320__62_ <= r_n_320__62_;
      r_320__61_ <= r_n_320__61_;
      r_320__60_ <= r_n_320__60_;
      r_320__59_ <= r_n_320__59_;
      r_320__58_ <= r_n_320__58_;
      r_320__57_ <= r_n_320__57_;
      r_320__56_ <= r_n_320__56_;
      r_320__55_ <= r_n_320__55_;
      r_320__54_ <= r_n_320__54_;
      r_320__53_ <= r_n_320__53_;
      r_320__52_ <= r_n_320__52_;
      r_320__51_ <= r_n_320__51_;
      r_320__50_ <= r_n_320__50_;
      r_320__49_ <= r_n_320__49_;
      r_320__48_ <= r_n_320__48_;
      r_320__47_ <= r_n_320__47_;
      r_320__46_ <= r_n_320__46_;
      r_320__45_ <= r_n_320__45_;
      r_320__44_ <= r_n_320__44_;
      r_320__43_ <= r_n_320__43_;
      r_320__42_ <= r_n_320__42_;
      r_320__41_ <= r_n_320__41_;
      r_320__40_ <= r_n_320__40_;
      r_320__39_ <= r_n_320__39_;
      r_320__38_ <= r_n_320__38_;
      r_320__37_ <= r_n_320__37_;
      r_320__36_ <= r_n_320__36_;
      r_320__35_ <= r_n_320__35_;
      r_320__34_ <= r_n_320__34_;
      r_320__33_ <= r_n_320__33_;
      r_320__32_ <= r_n_320__32_;
      r_320__31_ <= r_n_320__31_;
      r_320__30_ <= r_n_320__30_;
      r_320__29_ <= r_n_320__29_;
      r_320__28_ <= r_n_320__28_;
      r_320__27_ <= r_n_320__27_;
      r_320__26_ <= r_n_320__26_;
      r_320__25_ <= r_n_320__25_;
      r_320__24_ <= r_n_320__24_;
      r_320__23_ <= r_n_320__23_;
      r_320__22_ <= r_n_320__22_;
      r_320__21_ <= r_n_320__21_;
      r_320__20_ <= r_n_320__20_;
      r_320__19_ <= r_n_320__19_;
      r_320__18_ <= r_n_320__18_;
      r_320__17_ <= r_n_320__17_;
      r_320__16_ <= r_n_320__16_;
      r_320__15_ <= r_n_320__15_;
      r_320__14_ <= r_n_320__14_;
      r_320__13_ <= r_n_320__13_;
      r_320__12_ <= r_n_320__12_;
      r_320__11_ <= r_n_320__11_;
      r_320__10_ <= r_n_320__10_;
      r_320__9_ <= r_n_320__9_;
      r_320__8_ <= r_n_320__8_;
      r_320__7_ <= r_n_320__7_;
      r_320__6_ <= r_n_320__6_;
      r_320__5_ <= r_n_320__5_;
      r_320__4_ <= r_n_320__4_;
      r_320__3_ <= r_n_320__3_;
      r_320__2_ <= r_n_320__2_;
      r_320__1_ <= r_n_320__1_;
      r_320__0_ <= r_n_320__0_;
    end 
    if(N3905) begin
      r_321__63_ <= r_n_321__63_;
      r_321__62_ <= r_n_321__62_;
      r_321__61_ <= r_n_321__61_;
      r_321__60_ <= r_n_321__60_;
      r_321__59_ <= r_n_321__59_;
      r_321__58_ <= r_n_321__58_;
      r_321__57_ <= r_n_321__57_;
      r_321__56_ <= r_n_321__56_;
      r_321__55_ <= r_n_321__55_;
      r_321__54_ <= r_n_321__54_;
      r_321__53_ <= r_n_321__53_;
      r_321__52_ <= r_n_321__52_;
      r_321__51_ <= r_n_321__51_;
      r_321__50_ <= r_n_321__50_;
      r_321__49_ <= r_n_321__49_;
      r_321__48_ <= r_n_321__48_;
      r_321__47_ <= r_n_321__47_;
      r_321__46_ <= r_n_321__46_;
      r_321__45_ <= r_n_321__45_;
      r_321__44_ <= r_n_321__44_;
      r_321__43_ <= r_n_321__43_;
      r_321__42_ <= r_n_321__42_;
      r_321__41_ <= r_n_321__41_;
      r_321__40_ <= r_n_321__40_;
      r_321__39_ <= r_n_321__39_;
      r_321__38_ <= r_n_321__38_;
      r_321__37_ <= r_n_321__37_;
      r_321__36_ <= r_n_321__36_;
      r_321__35_ <= r_n_321__35_;
      r_321__34_ <= r_n_321__34_;
      r_321__33_ <= r_n_321__33_;
      r_321__32_ <= r_n_321__32_;
      r_321__31_ <= r_n_321__31_;
      r_321__30_ <= r_n_321__30_;
      r_321__29_ <= r_n_321__29_;
      r_321__28_ <= r_n_321__28_;
      r_321__27_ <= r_n_321__27_;
      r_321__26_ <= r_n_321__26_;
      r_321__25_ <= r_n_321__25_;
      r_321__24_ <= r_n_321__24_;
      r_321__23_ <= r_n_321__23_;
      r_321__22_ <= r_n_321__22_;
      r_321__21_ <= r_n_321__21_;
      r_321__20_ <= r_n_321__20_;
      r_321__19_ <= r_n_321__19_;
      r_321__18_ <= r_n_321__18_;
      r_321__17_ <= r_n_321__17_;
      r_321__16_ <= r_n_321__16_;
      r_321__15_ <= r_n_321__15_;
      r_321__14_ <= r_n_321__14_;
      r_321__13_ <= r_n_321__13_;
      r_321__12_ <= r_n_321__12_;
      r_321__11_ <= r_n_321__11_;
      r_321__10_ <= r_n_321__10_;
      r_321__9_ <= r_n_321__9_;
      r_321__8_ <= r_n_321__8_;
      r_321__7_ <= r_n_321__7_;
      r_321__6_ <= r_n_321__6_;
      r_321__5_ <= r_n_321__5_;
      r_321__4_ <= r_n_321__4_;
      r_321__3_ <= r_n_321__3_;
      r_321__2_ <= r_n_321__2_;
      r_321__1_ <= r_n_321__1_;
      r_321__0_ <= r_n_321__0_;
    end 
    if(N3906) begin
      r_322__63_ <= r_n_322__63_;
      r_322__62_ <= r_n_322__62_;
      r_322__61_ <= r_n_322__61_;
      r_322__60_ <= r_n_322__60_;
      r_322__59_ <= r_n_322__59_;
      r_322__58_ <= r_n_322__58_;
      r_322__57_ <= r_n_322__57_;
      r_322__56_ <= r_n_322__56_;
      r_322__55_ <= r_n_322__55_;
      r_322__54_ <= r_n_322__54_;
      r_322__53_ <= r_n_322__53_;
      r_322__52_ <= r_n_322__52_;
      r_322__51_ <= r_n_322__51_;
      r_322__50_ <= r_n_322__50_;
      r_322__49_ <= r_n_322__49_;
      r_322__48_ <= r_n_322__48_;
      r_322__47_ <= r_n_322__47_;
      r_322__46_ <= r_n_322__46_;
      r_322__45_ <= r_n_322__45_;
      r_322__44_ <= r_n_322__44_;
      r_322__43_ <= r_n_322__43_;
      r_322__42_ <= r_n_322__42_;
      r_322__41_ <= r_n_322__41_;
      r_322__40_ <= r_n_322__40_;
      r_322__39_ <= r_n_322__39_;
      r_322__38_ <= r_n_322__38_;
      r_322__37_ <= r_n_322__37_;
      r_322__36_ <= r_n_322__36_;
      r_322__35_ <= r_n_322__35_;
      r_322__34_ <= r_n_322__34_;
      r_322__33_ <= r_n_322__33_;
      r_322__32_ <= r_n_322__32_;
      r_322__31_ <= r_n_322__31_;
      r_322__30_ <= r_n_322__30_;
      r_322__29_ <= r_n_322__29_;
      r_322__28_ <= r_n_322__28_;
      r_322__27_ <= r_n_322__27_;
      r_322__26_ <= r_n_322__26_;
      r_322__25_ <= r_n_322__25_;
      r_322__24_ <= r_n_322__24_;
      r_322__23_ <= r_n_322__23_;
      r_322__22_ <= r_n_322__22_;
      r_322__21_ <= r_n_322__21_;
      r_322__20_ <= r_n_322__20_;
      r_322__19_ <= r_n_322__19_;
      r_322__18_ <= r_n_322__18_;
      r_322__17_ <= r_n_322__17_;
      r_322__16_ <= r_n_322__16_;
      r_322__15_ <= r_n_322__15_;
      r_322__14_ <= r_n_322__14_;
      r_322__13_ <= r_n_322__13_;
      r_322__12_ <= r_n_322__12_;
      r_322__11_ <= r_n_322__11_;
      r_322__10_ <= r_n_322__10_;
      r_322__9_ <= r_n_322__9_;
      r_322__8_ <= r_n_322__8_;
      r_322__7_ <= r_n_322__7_;
      r_322__6_ <= r_n_322__6_;
      r_322__5_ <= r_n_322__5_;
      r_322__4_ <= r_n_322__4_;
      r_322__3_ <= r_n_322__3_;
      r_322__2_ <= r_n_322__2_;
      r_322__1_ <= r_n_322__1_;
      r_322__0_ <= r_n_322__0_;
    end 
    if(N3907) begin
      r_323__63_ <= r_n_323__63_;
      r_323__62_ <= r_n_323__62_;
      r_323__61_ <= r_n_323__61_;
      r_323__60_ <= r_n_323__60_;
      r_323__59_ <= r_n_323__59_;
      r_323__58_ <= r_n_323__58_;
      r_323__57_ <= r_n_323__57_;
      r_323__56_ <= r_n_323__56_;
      r_323__55_ <= r_n_323__55_;
      r_323__54_ <= r_n_323__54_;
      r_323__53_ <= r_n_323__53_;
      r_323__52_ <= r_n_323__52_;
      r_323__51_ <= r_n_323__51_;
      r_323__50_ <= r_n_323__50_;
      r_323__49_ <= r_n_323__49_;
      r_323__48_ <= r_n_323__48_;
      r_323__47_ <= r_n_323__47_;
      r_323__46_ <= r_n_323__46_;
      r_323__45_ <= r_n_323__45_;
      r_323__44_ <= r_n_323__44_;
      r_323__43_ <= r_n_323__43_;
      r_323__42_ <= r_n_323__42_;
      r_323__41_ <= r_n_323__41_;
      r_323__40_ <= r_n_323__40_;
      r_323__39_ <= r_n_323__39_;
      r_323__38_ <= r_n_323__38_;
      r_323__37_ <= r_n_323__37_;
      r_323__36_ <= r_n_323__36_;
      r_323__35_ <= r_n_323__35_;
      r_323__34_ <= r_n_323__34_;
      r_323__33_ <= r_n_323__33_;
      r_323__32_ <= r_n_323__32_;
      r_323__31_ <= r_n_323__31_;
      r_323__30_ <= r_n_323__30_;
      r_323__29_ <= r_n_323__29_;
      r_323__28_ <= r_n_323__28_;
      r_323__27_ <= r_n_323__27_;
      r_323__26_ <= r_n_323__26_;
      r_323__25_ <= r_n_323__25_;
      r_323__24_ <= r_n_323__24_;
      r_323__23_ <= r_n_323__23_;
      r_323__22_ <= r_n_323__22_;
      r_323__21_ <= r_n_323__21_;
      r_323__20_ <= r_n_323__20_;
      r_323__19_ <= r_n_323__19_;
      r_323__18_ <= r_n_323__18_;
      r_323__17_ <= r_n_323__17_;
      r_323__16_ <= r_n_323__16_;
      r_323__15_ <= r_n_323__15_;
      r_323__14_ <= r_n_323__14_;
      r_323__13_ <= r_n_323__13_;
      r_323__12_ <= r_n_323__12_;
      r_323__11_ <= r_n_323__11_;
      r_323__10_ <= r_n_323__10_;
      r_323__9_ <= r_n_323__9_;
      r_323__8_ <= r_n_323__8_;
      r_323__7_ <= r_n_323__7_;
      r_323__6_ <= r_n_323__6_;
      r_323__5_ <= r_n_323__5_;
      r_323__4_ <= r_n_323__4_;
      r_323__3_ <= r_n_323__3_;
      r_323__2_ <= r_n_323__2_;
      r_323__1_ <= r_n_323__1_;
      r_323__0_ <= r_n_323__0_;
    end 
    if(N3908) begin
      r_324__63_ <= r_n_324__63_;
      r_324__62_ <= r_n_324__62_;
      r_324__61_ <= r_n_324__61_;
      r_324__60_ <= r_n_324__60_;
      r_324__59_ <= r_n_324__59_;
      r_324__58_ <= r_n_324__58_;
      r_324__57_ <= r_n_324__57_;
      r_324__56_ <= r_n_324__56_;
      r_324__55_ <= r_n_324__55_;
      r_324__54_ <= r_n_324__54_;
      r_324__53_ <= r_n_324__53_;
      r_324__52_ <= r_n_324__52_;
      r_324__51_ <= r_n_324__51_;
      r_324__50_ <= r_n_324__50_;
      r_324__49_ <= r_n_324__49_;
      r_324__48_ <= r_n_324__48_;
      r_324__47_ <= r_n_324__47_;
      r_324__46_ <= r_n_324__46_;
      r_324__45_ <= r_n_324__45_;
      r_324__44_ <= r_n_324__44_;
      r_324__43_ <= r_n_324__43_;
      r_324__42_ <= r_n_324__42_;
      r_324__41_ <= r_n_324__41_;
      r_324__40_ <= r_n_324__40_;
      r_324__39_ <= r_n_324__39_;
      r_324__38_ <= r_n_324__38_;
      r_324__37_ <= r_n_324__37_;
      r_324__36_ <= r_n_324__36_;
      r_324__35_ <= r_n_324__35_;
      r_324__34_ <= r_n_324__34_;
      r_324__33_ <= r_n_324__33_;
      r_324__32_ <= r_n_324__32_;
      r_324__31_ <= r_n_324__31_;
      r_324__30_ <= r_n_324__30_;
      r_324__29_ <= r_n_324__29_;
      r_324__28_ <= r_n_324__28_;
      r_324__27_ <= r_n_324__27_;
      r_324__26_ <= r_n_324__26_;
      r_324__25_ <= r_n_324__25_;
      r_324__24_ <= r_n_324__24_;
      r_324__23_ <= r_n_324__23_;
      r_324__22_ <= r_n_324__22_;
      r_324__21_ <= r_n_324__21_;
      r_324__20_ <= r_n_324__20_;
      r_324__19_ <= r_n_324__19_;
      r_324__18_ <= r_n_324__18_;
      r_324__17_ <= r_n_324__17_;
      r_324__16_ <= r_n_324__16_;
      r_324__15_ <= r_n_324__15_;
      r_324__14_ <= r_n_324__14_;
      r_324__13_ <= r_n_324__13_;
      r_324__12_ <= r_n_324__12_;
      r_324__11_ <= r_n_324__11_;
      r_324__10_ <= r_n_324__10_;
      r_324__9_ <= r_n_324__9_;
      r_324__8_ <= r_n_324__8_;
      r_324__7_ <= r_n_324__7_;
      r_324__6_ <= r_n_324__6_;
      r_324__5_ <= r_n_324__5_;
      r_324__4_ <= r_n_324__4_;
      r_324__3_ <= r_n_324__3_;
      r_324__2_ <= r_n_324__2_;
      r_324__1_ <= r_n_324__1_;
      r_324__0_ <= r_n_324__0_;
    end 
    if(N3909) begin
      r_325__63_ <= r_n_325__63_;
      r_325__62_ <= r_n_325__62_;
      r_325__61_ <= r_n_325__61_;
      r_325__60_ <= r_n_325__60_;
      r_325__59_ <= r_n_325__59_;
      r_325__58_ <= r_n_325__58_;
      r_325__57_ <= r_n_325__57_;
      r_325__56_ <= r_n_325__56_;
      r_325__55_ <= r_n_325__55_;
      r_325__54_ <= r_n_325__54_;
      r_325__53_ <= r_n_325__53_;
      r_325__52_ <= r_n_325__52_;
      r_325__51_ <= r_n_325__51_;
      r_325__50_ <= r_n_325__50_;
      r_325__49_ <= r_n_325__49_;
      r_325__48_ <= r_n_325__48_;
      r_325__47_ <= r_n_325__47_;
      r_325__46_ <= r_n_325__46_;
      r_325__45_ <= r_n_325__45_;
      r_325__44_ <= r_n_325__44_;
      r_325__43_ <= r_n_325__43_;
      r_325__42_ <= r_n_325__42_;
      r_325__41_ <= r_n_325__41_;
      r_325__40_ <= r_n_325__40_;
      r_325__39_ <= r_n_325__39_;
      r_325__38_ <= r_n_325__38_;
      r_325__37_ <= r_n_325__37_;
      r_325__36_ <= r_n_325__36_;
      r_325__35_ <= r_n_325__35_;
      r_325__34_ <= r_n_325__34_;
      r_325__33_ <= r_n_325__33_;
      r_325__32_ <= r_n_325__32_;
      r_325__31_ <= r_n_325__31_;
      r_325__30_ <= r_n_325__30_;
      r_325__29_ <= r_n_325__29_;
      r_325__28_ <= r_n_325__28_;
      r_325__27_ <= r_n_325__27_;
      r_325__26_ <= r_n_325__26_;
      r_325__25_ <= r_n_325__25_;
      r_325__24_ <= r_n_325__24_;
      r_325__23_ <= r_n_325__23_;
      r_325__22_ <= r_n_325__22_;
      r_325__21_ <= r_n_325__21_;
      r_325__20_ <= r_n_325__20_;
      r_325__19_ <= r_n_325__19_;
      r_325__18_ <= r_n_325__18_;
      r_325__17_ <= r_n_325__17_;
      r_325__16_ <= r_n_325__16_;
      r_325__15_ <= r_n_325__15_;
      r_325__14_ <= r_n_325__14_;
      r_325__13_ <= r_n_325__13_;
      r_325__12_ <= r_n_325__12_;
      r_325__11_ <= r_n_325__11_;
      r_325__10_ <= r_n_325__10_;
      r_325__9_ <= r_n_325__9_;
      r_325__8_ <= r_n_325__8_;
      r_325__7_ <= r_n_325__7_;
      r_325__6_ <= r_n_325__6_;
      r_325__5_ <= r_n_325__5_;
      r_325__4_ <= r_n_325__4_;
      r_325__3_ <= r_n_325__3_;
      r_325__2_ <= r_n_325__2_;
      r_325__1_ <= r_n_325__1_;
      r_325__0_ <= r_n_325__0_;
    end 
    if(N3910) begin
      r_326__63_ <= r_n_326__63_;
      r_326__62_ <= r_n_326__62_;
      r_326__61_ <= r_n_326__61_;
      r_326__60_ <= r_n_326__60_;
      r_326__59_ <= r_n_326__59_;
      r_326__58_ <= r_n_326__58_;
      r_326__57_ <= r_n_326__57_;
      r_326__56_ <= r_n_326__56_;
      r_326__55_ <= r_n_326__55_;
      r_326__54_ <= r_n_326__54_;
      r_326__53_ <= r_n_326__53_;
      r_326__52_ <= r_n_326__52_;
      r_326__51_ <= r_n_326__51_;
      r_326__50_ <= r_n_326__50_;
      r_326__49_ <= r_n_326__49_;
      r_326__48_ <= r_n_326__48_;
      r_326__47_ <= r_n_326__47_;
      r_326__46_ <= r_n_326__46_;
      r_326__45_ <= r_n_326__45_;
      r_326__44_ <= r_n_326__44_;
      r_326__43_ <= r_n_326__43_;
      r_326__42_ <= r_n_326__42_;
      r_326__41_ <= r_n_326__41_;
      r_326__40_ <= r_n_326__40_;
      r_326__39_ <= r_n_326__39_;
      r_326__38_ <= r_n_326__38_;
      r_326__37_ <= r_n_326__37_;
      r_326__36_ <= r_n_326__36_;
      r_326__35_ <= r_n_326__35_;
      r_326__34_ <= r_n_326__34_;
      r_326__33_ <= r_n_326__33_;
      r_326__32_ <= r_n_326__32_;
      r_326__31_ <= r_n_326__31_;
      r_326__30_ <= r_n_326__30_;
      r_326__29_ <= r_n_326__29_;
      r_326__28_ <= r_n_326__28_;
      r_326__27_ <= r_n_326__27_;
      r_326__26_ <= r_n_326__26_;
      r_326__25_ <= r_n_326__25_;
      r_326__24_ <= r_n_326__24_;
      r_326__23_ <= r_n_326__23_;
      r_326__22_ <= r_n_326__22_;
      r_326__21_ <= r_n_326__21_;
      r_326__20_ <= r_n_326__20_;
      r_326__19_ <= r_n_326__19_;
      r_326__18_ <= r_n_326__18_;
      r_326__17_ <= r_n_326__17_;
      r_326__16_ <= r_n_326__16_;
      r_326__15_ <= r_n_326__15_;
      r_326__14_ <= r_n_326__14_;
      r_326__13_ <= r_n_326__13_;
      r_326__12_ <= r_n_326__12_;
      r_326__11_ <= r_n_326__11_;
      r_326__10_ <= r_n_326__10_;
      r_326__9_ <= r_n_326__9_;
      r_326__8_ <= r_n_326__8_;
      r_326__7_ <= r_n_326__7_;
      r_326__6_ <= r_n_326__6_;
      r_326__5_ <= r_n_326__5_;
      r_326__4_ <= r_n_326__4_;
      r_326__3_ <= r_n_326__3_;
      r_326__2_ <= r_n_326__2_;
      r_326__1_ <= r_n_326__1_;
      r_326__0_ <= r_n_326__0_;
    end 
    if(N3911) begin
      r_327__63_ <= r_n_327__63_;
      r_327__62_ <= r_n_327__62_;
      r_327__61_ <= r_n_327__61_;
      r_327__60_ <= r_n_327__60_;
      r_327__59_ <= r_n_327__59_;
      r_327__58_ <= r_n_327__58_;
      r_327__57_ <= r_n_327__57_;
      r_327__56_ <= r_n_327__56_;
      r_327__55_ <= r_n_327__55_;
      r_327__54_ <= r_n_327__54_;
      r_327__53_ <= r_n_327__53_;
      r_327__52_ <= r_n_327__52_;
      r_327__51_ <= r_n_327__51_;
      r_327__50_ <= r_n_327__50_;
      r_327__49_ <= r_n_327__49_;
      r_327__48_ <= r_n_327__48_;
      r_327__47_ <= r_n_327__47_;
      r_327__46_ <= r_n_327__46_;
      r_327__45_ <= r_n_327__45_;
      r_327__44_ <= r_n_327__44_;
      r_327__43_ <= r_n_327__43_;
      r_327__42_ <= r_n_327__42_;
      r_327__41_ <= r_n_327__41_;
      r_327__40_ <= r_n_327__40_;
      r_327__39_ <= r_n_327__39_;
      r_327__38_ <= r_n_327__38_;
      r_327__37_ <= r_n_327__37_;
      r_327__36_ <= r_n_327__36_;
      r_327__35_ <= r_n_327__35_;
      r_327__34_ <= r_n_327__34_;
      r_327__33_ <= r_n_327__33_;
      r_327__32_ <= r_n_327__32_;
      r_327__31_ <= r_n_327__31_;
      r_327__30_ <= r_n_327__30_;
      r_327__29_ <= r_n_327__29_;
      r_327__28_ <= r_n_327__28_;
      r_327__27_ <= r_n_327__27_;
      r_327__26_ <= r_n_327__26_;
      r_327__25_ <= r_n_327__25_;
      r_327__24_ <= r_n_327__24_;
      r_327__23_ <= r_n_327__23_;
      r_327__22_ <= r_n_327__22_;
      r_327__21_ <= r_n_327__21_;
      r_327__20_ <= r_n_327__20_;
      r_327__19_ <= r_n_327__19_;
      r_327__18_ <= r_n_327__18_;
      r_327__17_ <= r_n_327__17_;
      r_327__16_ <= r_n_327__16_;
      r_327__15_ <= r_n_327__15_;
      r_327__14_ <= r_n_327__14_;
      r_327__13_ <= r_n_327__13_;
      r_327__12_ <= r_n_327__12_;
      r_327__11_ <= r_n_327__11_;
      r_327__10_ <= r_n_327__10_;
      r_327__9_ <= r_n_327__9_;
      r_327__8_ <= r_n_327__8_;
      r_327__7_ <= r_n_327__7_;
      r_327__6_ <= r_n_327__6_;
      r_327__5_ <= r_n_327__5_;
      r_327__4_ <= r_n_327__4_;
      r_327__3_ <= r_n_327__3_;
      r_327__2_ <= r_n_327__2_;
      r_327__1_ <= r_n_327__1_;
      r_327__0_ <= r_n_327__0_;
    end 
    if(N3912) begin
      r_328__63_ <= r_n_328__63_;
      r_328__62_ <= r_n_328__62_;
      r_328__61_ <= r_n_328__61_;
      r_328__60_ <= r_n_328__60_;
      r_328__59_ <= r_n_328__59_;
      r_328__58_ <= r_n_328__58_;
      r_328__57_ <= r_n_328__57_;
      r_328__56_ <= r_n_328__56_;
      r_328__55_ <= r_n_328__55_;
      r_328__54_ <= r_n_328__54_;
      r_328__53_ <= r_n_328__53_;
      r_328__52_ <= r_n_328__52_;
      r_328__51_ <= r_n_328__51_;
      r_328__50_ <= r_n_328__50_;
      r_328__49_ <= r_n_328__49_;
      r_328__48_ <= r_n_328__48_;
      r_328__47_ <= r_n_328__47_;
      r_328__46_ <= r_n_328__46_;
      r_328__45_ <= r_n_328__45_;
      r_328__44_ <= r_n_328__44_;
      r_328__43_ <= r_n_328__43_;
      r_328__42_ <= r_n_328__42_;
      r_328__41_ <= r_n_328__41_;
      r_328__40_ <= r_n_328__40_;
      r_328__39_ <= r_n_328__39_;
      r_328__38_ <= r_n_328__38_;
      r_328__37_ <= r_n_328__37_;
      r_328__36_ <= r_n_328__36_;
      r_328__35_ <= r_n_328__35_;
      r_328__34_ <= r_n_328__34_;
      r_328__33_ <= r_n_328__33_;
      r_328__32_ <= r_n_328__32_;
      r_328__31_ <= r_n_328__31_;
      r_328__30_ <= r_n_328__30_;
      r_328__29_ <= r_n_328__29_;
      r_328__28_ <= r_n_328__28_;
      r_328__27_ <= r_n_328__27_;
      r_328__26_ <= r_n_328__26_;
      r_328__25_ <= r_n_328__25_;
      r_328__24_ <= r_n_328__24_;
      r_328__23_ <= r_n_328__23_;
      r_328__22_ <= r_n_328__22_;
      r_328__21_ <= r_n_328__21_;
      r_328__20_ <= r_n_328__20_;
      r_328__19_ <= r_n_328__19_;
      r_328__18_ <= r_n_328__18_;
      r_328__17_ <= r_n_328__17_;
      r_328__16_ <= r_n_328__16_;
      r_328__15_ <= r_n_328__15_;
      r_328__14_ <= r_n_328__14_;
      r_328__13_ <= r_n_328__13_;
      r_328__12_ <= r_n_328__12_;
      r_328__11_ <= r_n_328__11_;
      r_328__10_ <= r_n_328__10_;
      r_328__9_ <= r_n_328__9_;
      r_328__8_ <= r_n_328__8_;
      r_328__7_ <= r_n_328__7_;
      r_328__6_ <= r_n_328__6_;
      r_328__5_ <= r_n_328__5_;
      r_328__4_ <= r_n_328__4_;
      r_328__3_ <= r_n_328__3_;
      r_328__2_ <= r_n_328__2_;
      r_328__1_ <= r_n_328__1_;
      r_328__0_ <= r_n_328__0_;
    end 
    if(N3913) begin
      r_329__63_ <= r_n_329__63_;
      r_329__62_ <= r_n_329__62_;
      r_329__61_ <= r_n_329__61_;
      r_329__60_ <= r_n_329__60_;
      r_329__59_ <= r_n_329__59_;
      r_329__58_ <= r_n_329__58_;
      r_329__57_ <= r_n_329__57_;
      r_329__56_ <= r_n_329__56_;
      r_329__55_ <= r_n_329__55_;
      r_329__54_ <= r_n_329__54_;
      r_329__53_ <= r_n_329__53_;
      r_329__52_ <= r_n_329__52_;
      r_329__51_ <= r_n_329__51_;
      r_329__50_ <= r_n_329__50_;
      r_329__49_ <= r_n_329__49_;
      r_329__48_ <= r_n_329__48_;
      r_329__47_ <= r_n_329__47_;
      r_329__46_ <= r_n_329__46_;
      r_329__45_ <= r_n_329__45_;
      r_329__44_ <= r_n_329__44_;
      r_329__43_ <= r_n_329__43_;
      r_329__42_ <= r_n_329__42_;
      r_329__41_ <= r_n_329__41_;
      r_329__40_ <= r_n_329__40_;
      r_329__39_ <= r_n_329__39_;
      r_329__38_ <= r_n_329__38_;
      r_329__37_ <= r_n_329__37_;
      r_329__36_ <= r_n_329__36_;
      r_329__35_ <= r_n_329__35_;
      r_329__34_ <= r_n_329__34_;
      r_329__33_ <= r_n_329__33_;
      r_329__32_ <= r_n_329__32_;
      r_329__31_ <= r_n_329__31_;
      r_329__30_ <= r_n_329__30_;
      r_329__29_ <= r_n_329__29_;
      r_329__28_ <= r_n_329__28_;
      r_329__27_ <= r_n_329__27_;
      r_329__26_ <= r_n_329__26_;
      r_329__25_ <= r_n_329__25_;
      r_329__24_ <= r_n_329__24_;
      r_329__23_ <= r_n_329__23_;
      r_329__22_ <= r_n_329__22_;
      r_329__21_ <= r_n_329__21_;
      r_329__20_ <= r_n_329__20_;
      r_329__19_ <= r_n_329__19_;
      r_329__18_ <= r_n_329__18_;
      r_329__17_ <= r_n_329__17_;
      r_329__16_ <= r_n_329__16_;
      r_329__15_ <= r_n_329__15_;
      r_329__14_ <= r_n_329__14_;
      r_329__13_ <= r_n_329__13_;
      r_329__12_ <= r_n_329__12_;
      r_329__11_ <= r_n_329__11_;
      r_329__10_ <= r_n_329__10_;
      r_329__9_ <= r_n_329__9_;
      r_329__8_ <= r_n_329__8_;
      r_329__7_ <= r_n_329__7_;
      r_329__6_ <= r_n_329__6_;
      r_329__5_ <= r_n_329__5_;
      r_329__4_ <= r_n_329__4_;
      r_329__3_ <= r_n_329__3_;
      r_329__2_ <= r_n_329__2_;
      r_329__1_ <= r_n_329__1_;
      r_329__0_ <= r_n_329__0_;
    end 
    if(N3914) begin
      r_330__63_ <= r_n_330__63_;
      r_330__62_ <= r_n_330__62_;
      r_330__61_ <= r_n_330__61_;
      r_330__60_ <= r_n_330__60_;
      r_330__59_ <= r_n_330__59_;
      r_330__58_ <= r_n_330__58_;
      r_330__57_ <= r_n_330__57_;
      r_330__56_ <= r_n_330__56_;
      r_330__55_ <= r_n_330__55_;
      r_330__54_ <= r_n_330__54_;
      r_330__53_ <= r_n_330__53_;
      r_330__52_ <= r_n_330__52_;
      r_330__51_ <= r_n_330__51_;
      r_330__50_ <= r_n_330__50_;
      r_330__49_ <= r_n_330__49_;
      r_330__48_ <= r_n_330__48_;
      r_330__47_ <= r_n_330__47_;
      r_330__46_ <= r_n_330__46_;
      r_330__45_ <= r_n_330__45_;
      r_330__44_ <= r_n_330__44_;
      r_330__43_ <= r_n_330__43_;
      r_330__42_ <= r_n_330__42_;
      r_330__41_ <= r_n_330__41_;
      r_330__40_ <= r_n_330__40_;
      r_330__39_ <= r_n_330__39_;
      r_330__38_ <= r_n_330__38_;
      r_330__37_ <= r_n_330__37_;
      r_330__36_ <= r_n_330__36_;
      r_330__35_ <= r_n_330__35_;
      r_330__34_ <= r_n_330__34_;
      r_330__33_ <= r_n_330__33_;
      r_330__32_ <= r_n_330__32_;
      r_330__31_ <= r_n_330__31_;
      r_330__30_ <= r_n_330__30_;
      r_330__29_ <= r_n_330__29_;
      r_330__28_ <= r_n_330__28_;
      r_330__27_ <= r_n_330__27_;
      r_330__26_ <= r_n_330__26_;
      r_330__25_ <= r_n_330__25_;
      r_330__24_ <= r_n_330__24_;
      r_330__23_ <= r_n_330__23_;
      r_330__22_ <= r_n_330__22_;
      r_330__21_ <= r_n_330__21_;
      r_330__20_ <= r_n_330__20_;
      r_330__19_ <= r_n_330__19_;
      r_330__18_ <= r_n_330__18_;
      r_330__17_ <= r_n_330__17_;
      r_330__16_ <= r_n_330__16_;
      r_330__15_ <= r_n_330__15_;
      r_330__14_ <= r_n_330__14_;
      r_330__13_ <= r_n_330__13_;
      r_330__12_ <= r_n_330__12_;
      r_330__11_ <= r_n_330__11_;
      r_330__10_ <= r_n_330__10_;
      r_330__9_ <= r_n_330__9_;
      r_330__8_ <= r_n_330__8_;
      r_330__7_ <= r_n_330__7_;
      r_330__6_ <= r_n_330__6_;
      r_330__5_ <= r_n_330__5_;
      r_330__4_ <= r_n_330__4_;
      r_330__3_ <= r_n_330__3_;
      r_330__2_ <= r_n_330__2_;
      r_330__1_ <= r_n_330__1_;
      r_330__0_ <= r_n_330__0_;
    end 
    if(N3915) begin
      r_331__63_ <= r_n_331__63_;
      r_331__62_ <= r_n_331__62_;
      r_331__61_ <= r_n_331__61_;
      r_331__60_ <= r_n_331__60_;
      r_331__59_ <= r_n_331__59_;
      r_331__58_ <= r_n_331__58_;
      r_331__57_ <= r_n_331__57_;
      r_331__56_ <= r_n_331__56_;
      r_331__55_ <= r_n_331__55_;
      r_331__54_ <= r_n_331__54_;
      r_331__53_ <= r_n_331__53_;
      r_331__52_ <= r_n_331__52_;
      r_331__51_ <= r_n_331__51_;
      r_331__50_ <= r_n_331__50_;
      r_331__49_ <= r_n_331__49_;
      r_331__48_ <= r_n_331__48_;
      r_331__47_ <= r_n_331__47_;
      r_331__46_ <= r_n_331__46_;
      r_331__45_ <= r_n_331__45_;
      r_331__44_ <= r_n_331__44_;
      r_331__43_ <= r_n_331__43_;
      r_331__42_ <= r_n_331__42_;
      r_331__41_ <= r_n_331__41_;
      r_331__40_ <= r_n_331__40_;
      r_331__39_ <= r_n_331__39_;
      r_331__38_ <= r_n_331__38_;
      r_331__37_ <= r_n_331__37_;
      r_331__36_ <= r_n_331__36_;
      r_331__35_ <= r_n_331__35_;
      r_331__34_ <= r_n_331__34_;
      r_331__33_ <= r_n_331__33_;
      r_331__32_ <= r_n_331__32_;
      r_331__31_ <= r_n_331__31_;
      r_331__30_ <= r_n_331__30_;
      r_331__29_ <= r_n_331__29_;
      r_331__28_ <= r_n_331__28_;
      r_331__27_ <= r_n_331__27_;
      r_331__26_ <= r_n_331__26_;
      r_331__25_ <= r_n_331__25_;
      r_331__24_ <= r_n_331__24_;
      r_331__23_ <= r_n_331__23_;
      r_331__22_ <= r_n_331__22_;
      r_331__21_ <= r_n_331__21_;
      r_331__20_ <= r_n_331__20_;
      r_331__19_ <= r_n_331__19_;
      r_331__18_ <= r_n_331__18_;
      r_331__17_ <= r_n_331__17_;
      r_331__16_ <= r_n_331__16_;
      r_331__15_ <= r_n_331__15_;
      r_331__14_ <= r_n_331__14_;
      r_331__13_ <= r_n_331__13_;
      r_331__12_ <= r_n_331__12_;
      r_331__11_ <= r_n_331__11_;
      r_331__10_ <= r_n_331__10_;
      r_331__9_ <= r_n_331__9_;
      r_331__8_ <= r_n_331__8_;
      r_331__7_ <= r_n_331__7_;
      r_331__6_ <= r_n_331__6_;
      r_331__5_ <= r_n_331__5_;
      r_331__4_ <= r_n_331__4_;
      r_331__3_ <= r_n_331__3_;
      r_331__2_ <= r_n_331__2_;
      r_331__1_ <= r_n_331__1_;
      r_331__0_ <= r_n_331__0_;
    end 
    if(N3916) begin
      r_332__63_ <= r_n_332__63_;
      r_332__62_ <= r_n_332__62_;
      r_332__61_ <= r_n_332__61_;
      r_332__60_ <= r_n_332__60_;
      r_332__59_ <= r_n_332__59_;
      r_332__58_ <= r_n_332__58_;
      r_332__57_ <= r_n_332__57_;
      r_332__56_ <= r_n_332__56_;
      r_332__55_ <= r_n_332__55_;
      r_332__54_ <= r_n_332__54_;
      r_332__53_ <= r_n_332__53_;
      r_332__52_ <= r_n_332__52_;
      r_332__51_ <= r_n_332__51_;
      r_332__50_ <= r_n_332__50_;
      r_332__49_ <= r_n_332__49_;
      r_332__48_ <= r_n_332__48_;
      r_332__47_ <= r_n_332__47_;
      r_332__46_ <= r_n_332__46_;
      r_332__45_ <= r_n_332__45_;
      r_332__44_ <= r_n_332__44_;
      r_332__43_ <= r_n_332__43_;
      r_332__42_ <= r_n_332__42_;
      r_332__41_ <= r_n_332__41_;
      r_332__40_ <= r_n_332__40_;
      r_332__39_ <= r_n_332__39_;
      r_332__38_ <= r_n_332__38_;
      r_332__37_ <= r_n_332__37_;
      r_332__36_ <= r_n_332__36_;
      r_332__35_ <= r_n_332__35_;
      r_332__34_ <= r_n_332__34_;
      r_332__33_ <= r_n_332__33_;
      r_332__32_ <= r_n_332__32_;
      r_332__31_ <= r_n_332__31_;
      r_332__30_ <= r_n_332__30_;
      r_332__29_ <= r_n_332__29_;
      r_332__28_ <= r_n_332__28_;
      r_332__27_ <= r_n_332__27_;
      r_332__26_ <= r_n_332__26_;
      r_332__25_ <= r_n_332__25_;
      r_332__24_ <= r_n_332__24_;
      r_332__23_ <= r_n_332__23_;
      r_332__22_ <= r_n_332__22_;
      r_332__21_ <= r_n_332__21_;
      r_332__20_ <= r_n_332__20_;
      r_332__19_ <= r_n_332__19_;
      r_332__18_ <= r_n_332__18_;
      r_332__17_ <= r_n_332__17_;
      r_332__16_ <= r_n_332__16_;
      r_332__15_ <= r_n_332__15_;
      r_332__14_ <= r_n_332__14_;
      r_332__13_ <= r_n_332__13_;
      r_332__12_ <= r_n_332__12_;
      r_332__11_ <= r_n_332__11_;
      r_332__10_ <= r_n_332__10_;
      r_332__9_ <= r_n_332__9_;
      r_332__8_ <= r_n_332__8_;
      r_332__7_ <= r_n_332__7_;
      r_332__6_ <= r_n_332__6_;
      r_332__5_ <= r_n_332__5_;
      r_332__4_ <= r_n_332__4_;
      r_332__3_ <= r_n_332__3_;
      r_332__2_ <= r_n_332__2_;
      r_332__1_ <= r_n_332__1_;
      r_332__0_ <= r_n_332__0_;
    end 
    if(N3917) begin
      r_333__63_ <= r_n_333__63_;
      r_333__62_ <= r_n_333__62_;
      r_333__61_ <= r_n_333__61_;
      r_333__60_ <= r_n_333__60_;
      r_333__59_ <= r_n_333__59_;
      r_333__58_ <= r_n_333__58_;
      r_333__57_ <= r_n_333__57_;
      r_333__56_ <= r_n_333__56_;
      r_333__55_ <= r_n_333__55_;
      r_333__54_ <= r_n_333__54_;
      r_333__53_ <= r_n_333__53_;
      r_333__52_ <= r_n_333__52_;
      r_333__51_ <= r_n_333__51_;
      r_333__50_ <= r_n_333__50_;
      r_333__49_ <= r_n_333__49_;
      r_333__48_ <= r_n_333__48_;
      r_333__47_ <= r_n_333__47_;
      r_333__46_ <= r_n_333__46_;
      r_333__45_ <= r_n_333__45_;
      r_333__44_ <= r_n_333__44_;
      r_333__43_ <= r_n_333__43_;
      r_333__42_ <= r_n_333__42_;
      r_333__41_ <= r_n_333__41_;
      r_333__40_ <= r_n_333__40_;
      r_333__39_ <= r_n_333__39_;
      r_333__38_ <= r_n_333__38_;
      r_333__37_ <= r_n_333__37_;
      r_333__36_ <= r_n_333__36_;
      r_333__35_ <= r_n_333__35_;
      r_333__34_ <= r_n_333__34_;
      r_333__33_ <= r_n_333__33_;
      r_333__32_ <= r_n_333__32_;
      r_333__31_ <= r_n_333__31_;
      r_333__30_ <= r_n_333__30_;
      r_333__29_ <= r_n_333__29_;
      r_333__28_ <= r_n_333__28_;
      r_333__27_ <= r_n_333__27_;
      r_333__26_ <= r_n_333__26_;
      r_333__25_ <= r_n_333__25_;
      r_333__24_ <= r_n_333__24_;
      r_333__23_ <= r_n_333__23_;
      r_333__22_ <= r_n_333__22_;
      r_333__21_ <= r_n_333__21_;
      r_333__20_ <= r_n_333__20_;
      r_333__19_ <= r_n_333__19_;
      r_333__18_ <= r_n_333__18_;
      r_333__17_ <= r_n_333__17_;
      r_333__16_ <= r_n_333__16_;
      r_333__15_ <= r_n_333__15_;
      r_333__14_ <= r_n_333__14_;
      r_333__13_ <= r_n_333__13_;
      r_333__12_ <= r_n_333__12_;
      r_333__11_ <= r_n_333__11_;
      r_333__10_ <= r_n_333__10_;
      r_333__9_ <= r_n_333__9_;
      r_333__8_ <= r_n_333__8_;
      r_333__7_ <= r_n_333__7_;
      r_333__6_ <= r_n_333__6_;
      r_333__5_ <= r_n_333__5_;
      r_333__4_ <= r_n_333__4_;
      r_333__3_ <= r_n_333__3_;
      r_333__2_ <= r_n_333__2_;
      r_333__1_ <= r_n_333__1_;
      r_333__0_ <= r_n_333__0_;
    end 
    if(N3918) begin
      r_334__63_ <= r_n_334__63_;
      r_334__62_ <= r_n_334__62_;
      r_334__61_ <= r_n_334__61_;
      r_334__60_ <= r_n_334__60_;
      r_334__59_ <= r_n_334__59_;
      r_334__58_ <= r_n_334__58_;
      r_334__57_ <= r_n_334__57_;
      r_334__56_ <= r_n_334__56_;
      r_334__55_ <= r_n_334__55_;
      r_334__54_ <= r_n_334__54_;
      r_334__53_ <= r_n_334__53_;
      r_334__52_ <= r_n_334__52_;
      r_334__51_ <= r_n_334__51_;
      r_334__50_ <= r_n_334__50_;
      r_334__49_ <= r_n_334__49_;
      r_334__48_ <= r_n_334__48_;
      r_334__47_ <= r_n_334__47_;
      r_334__46_ <= r_n_334__46_;
      r_334__45_ <= r_n_334__45_;
      r_334__44_ <= r_n_334__44_;
      r_334__43_ <= r_n_334__43_;
      r_334__42_ <= r_n_334__42_;
      r_334__41_ <= r_n_334__41_;
      r_334__40_ <= r_n_334__40_;
      r_334__39_ <= r_n_334__39_;
      r_334__38_ <= r_n_334__38_;
      r_334__37_ <= r_n_334__37_;
      r_334__36_ <= r_n_334__36_;
      r_334__35_ <= r_n_334__35_;
      r_334__34_ <= r_n_334__34_;
      r_334__33_ <= r_n_334__33_;
      r_334__32_ <= r_n_334__32_;
      r_334__31_ <= r_n_334__31_;
      r_334__30_ <= r_n_334__30_;
      r_334__29_ <= r_n_334__29_;
      r_334__28_ <= r_n_334__28_;
      r_334__27_ <= r_n_334__27_;
      r_334__26_ <= r_n_334__26_;
      r_334__25_ <= r_n_334__25_;
      r_334__24_ <= r_n_334__24_;
      r_334__23_ <= r_n_334__23_;
      r_334__22_ <= r_n_334__22_;
      r_334__21_ <= r_n_334__21_;
      r_334__20_ <= r_n_334__20_;
      r_334__19_ <= r_n_334__19_;
      r_334__18_ <= r_n_334__18_;
      r_334__17_ <= r_n_334__17_;
      r_334__16_ <= r_n_334__16_;
      r_334__15_ <= r_n_334__15_;
      r_334__14_ <= r_n_334__14_;
      r_334__13_ <= r_n_334__13_;
      r_334__12_ <= r_n_334__12_;
      r_334__11_ <= r_n_334__11_;
      r_334__10_ <= r_n_334__10_;
      r_334__9_ <= r_n_334__9_;
      r_334__8_ <= r_n_334__8_;
      r_334__7_ <= r_n_334__7_;
      r_334__6_ <= r_n_334__6_;
      r_334__5_ <= r_n_334__5_;
      r_334__4_ <= r_n_334__4_;
      r_334__3_ <= r_n_334__3_;
      r_334__2_ <= r_n_334__2_;
      r_334__1_ <= r_n_334__1_;
      r_334__0_ <= r_n_334__0_;
    end 
    if(N3919) begin
      r_335__63_ <= r_n_335__63_;
      r_335__62_ <= r_n_335__62_;
      r_335__61_ <= r_n_335__61_;
      r_335__60_ <= r_n_335__60_;
      r_335__59_ <= r_n_335__59_;
      r_335__58_ <= r_n_335__58_;
      r_335__57_ <= r_n_335__57_;
      r_335__56_ <= r_n_335__56_;
      r_335__55_ <= r_n_335__55_;
      r_335__54_ <= r_n_335__54_;
      r_335__53_ <= r_n_335__53_;
      r_335__52_ <= r_n_335__52_;
      r_335__51_ <= r_n_335__51_;
      r_335__50_ <= r_n_335__50_;
      r_335__49_ <= r_n_335__49_;
      r_335__48_ <= r_n_335__48_;
      r_335__47_ <= r_n_335__47_;
      r_335__46_ <= r_n_335__46_;
      r_335__45_ <= r_n_335__45_;
      r_335__44_ <= r_n_335__44_;
      r_335__43_ <= r_n_335__43_;
      r_335__42_ <= r_n_335__42_;
      r_335__41_ <= r_n_335__41_;
      r_335__40_ <= r_n_335__40_;
      r_335__39_ <= r_n_335__39_;
      r_335__38_ <= r_n_335__38_;
      r_335__37_ <= r_n_335__37_;
      r_335__36_ <= r_n_335__36_;
      r_335__35_ <= r_n_335__35_;
      r_335__34_ <= r_n_335__34_;
      r_335__33_ <= r_n_335__33_;
      r_335__32_ <= r_n_335__32_;
      r_335__31_ <= r_n_335__31_;
      r_335__30_ <= r_n_335__30_;
      r_335__29_ <= r_n_335__29_;
      r_335__28_ <= r_n_335__28_;
      r_335__27_ <= r_n_335__27_;
      r_335__26_ <= r_n_335__26_;
      r_335__25_ <= r_n_335__25_;
      r_335__24_ <= r_n_335__24_;
      r_335__23_ <= r_n_335__23_;
      r_335__22_ <= r_n_335__22_;
      r_335__21_ <= r_n_335__21_;
      r_335__20_ <= r_n_335__20_;
      r_335__19_ <= r_n_335__19_;
      r_335__18_ <= r_n_335__18_;
      r_335__17_ <= r_n_335__17_;
      r_335__16_ <= r_n_335__16_;
      r_335__15_ <= r_n_335__15_;
      r_335__14_ <= r_n_335__14_;
      r_335__13_ <= r_n_335__13_;
      r_335__12_ <= r_n_335__12_;
      r_335__11_ <= r_n_335__11_;
      r_335__10_ <= r_n_335__10_;
      r_335__9_ <= r_n_335__9_;
      r_335__8_ <= r_n_335__8_;
      r_335__7_ <= r_n_335__7_;
      r_335__6_ <= r_n_335__6_;
      r_335__5_ <= r_n_335__5_;
      r_335__4_ <= r_n_335__4_;
      r_335__3_ <= r_n_335__3_;
      r_335__2_ <= r_n_335__2_;
      r_335__1_ <= r_n_335__1_;
      r_335__0_ <= r_n_335__0_;
    end 
    if(N3920) begin
      r_336__63_ <= r_n_336__63_;
      r_336__62_ <= r_n_336__62_;
      r_336__61_ <= r_n_336__61_;
      r_336__60_ <= r_n_336__60_;
      r_336__59_ <= r_n_336__59_;
      r_336__58_ <= r_n_336__58_;
      r_336__57_ <= r_n_336__57_;
      r_336__56_ <= r_n_336__56_;
      r_336__55_ <= r_n_336__55_;
      r_336__54_ <= r_n_336__54_;
      r_336__53_ <= r_n_336__53_;
      r_336__52_ <= r_n_336__52_;
      r_336__51_ <= r_n_336__51_;
      r_336__50_ <= r_n_336__50_;
      r_336__49_ <= r_n_336__49_;
      r_336__48_ <= r_n_336__48_;
      r_336__47_ <= r_n_336__47_;
      r_336__46_ <= r_n_336__46_;
      r_336__45_ <= r_n_336__45_;
      r_336__44_ <= r_n_336__44_;
      r_336__43_ <= r_n_336__43_;
      r_336__42_ <= r_n_336__42_;
      r_336__41_ <= r_n_336__41_;
      r_336__40_ <= r_n_336__40_;
      r_336__39_ <= r_n_336__39_;
      r_336__38_ <= r_n_336__38_;
      r_336__37_ <= r_n_336__37_;
      r_336__36_ <= r_n_336__36_;
      r_336__35_ <= r_n_336__35_;
      r_336__34_ <= r_n_336__34_;
      r_336__33_ <= r_n_336__33_;
      r_336__32_ <= r_n_336__32_;
      r_336__31_ <= r_n_336__31_;
      r_336__30_ <= r_n_336__30_;
      r_336__29_ <= r_n_336__29_;
      r_336__28_ <= r_n_336__28_;
      r_336__27_ <= r_n_336__27_;
      r_336__26_ <= r_n_336__26_;
      r_336__25_ <= r_n_336__25_;
      r_336__24_ <= r_n_336__24_;
      r_336__23_ <= r_n_336__23_;
      r_336__22_ <= r_n_336__22_;
      r_336__21_ <= r_n_336__21_;
      r_336__20_ <= r_n_336__20_;
      r_336__19_ <= r_n_336__19_;
      r_336__18_ <= r_n_336__18_;
      r_336__17_ <= r_n_336__17_;
      r_336__16_ <= r_n_336__16_;
      r_336__15_ <= r_n_336__15_;
      r_336__14_ <= r_n_336__14_;
      r_336__13_ <= r_n_336__13_;
      r_336__12_ <= r_n_336__12_;
      r_336__11_ <= r_n_336__11_;
      r_336__10_ <= r_n_336__10_;
      r_336__9_ <= r_n_336__9_;
      r_336__8_ <= r_n_336__8_;
      r_336__7_ <= r_n_336__7_;
      r_336__6_ <= r_n_336__6_;
      r_336__5_ <= r_n_336__5_;
      r_336__4_ <= r_n_336__4_;
      r_336__3_ <= r_n_336__3_;
      r_336__2_ <= r_n_336__2_;
      r_336__1_ <= r_n_336__1_;
      r_336__0_ <= r_n_336__0_;
    end 
    if(N3921) begin
      r_337__63_ <= r_n_337__63_;
      r_337__62_ <= r_n_337__62_;
      r_337__61_ <= r_n_337__61_;
      r_337__60_ <= r_n_337__60_;
      r_337__59_ <= r_n_337__59_;
      r_337__58_ <= r_n_337__58_;
      r_337__57_ <= r_n_337__57_;
      r_337__56_ <= r_n_337__56_;
      r_337__55_ <= r_n_337__55_;
      r_337__54_ <= r_n_337__54_;
      r_337__53_ <= r_n_337__53_;
      r_337__52_ <= r_n_337__52_;
      r_337__51_ <= r_n_337__51_;
      r_337__50_ <= r_n_337__50_;
      r_337__49_ <= r_n_337__49_;
      r_337__48_ <= r_n_337__48_;
      r_337__47_ <= r_n_337__47_;
      r_337__46_ <= r_n_337__46_;
      r_337__45_ <= r_n_337__45_;
      r_337__44_ <= r_n_337__44_;
      r_337__43_ <= r_n_337__43_;
      r_337__42_ <= r_n_337__42_;
      r_337__41_ <= r_n_337__41_;
      r_337__40_ <= r_n_337__40_;
      r_337__39_ <= r_n_337__39_;
      r_337__38_ <= r_n_337__38_;
      r_337__37_ <= r_n_337__37_;
      r_337__36_ <= r_n_337__36_;
      r_337__35_ <= r_n_337__35_;
      r_337__34_ <= r_n_337__34_;
      r_337__33_ <= r_n_337__33_;
      r_337__32_ <= r_n_337__32_;
      r_337__31_ <= r_n_337__31_;
      r_337__30_ <= r_n_337__30_;
      r_337__29_ <= r_n_337__29_;
      r_337__28_ <= r_n_337__28_;
      r_337__27_ <= r_n_337__27_;
      r_337__26_ <= r_n_337__26_;
      r_337__25_ <= r_n_337__25_;
      r_337__24_ <= r_n_337__24_;
      r_337__23_ <= r_n_337__23_;
      r_337__22_ <= r_n_337__22_;
      r_337__21_ <= r_n_337__21_;
      r_337__20_ <= r_n_337__20_;
      r_337__19_ <= r_n_337__19_;
      r_337__18_ <= r_n_337__18_;
      r_337__17_ <= r_n_337__17_;
      r_337__16_ <= r_n_337__16_;
      r_337__15_ <= r_n_337__15_;
      r_337__14_ <= r_n_337__14_;
      r_337__13_ <= r_n_337__13_;
      r_337__12_ <= r_n_337__12_;
      r_337__11_ <= r_n_337__11_;
      r_337__10_ <= r_n_337__10_;
      r_337__9_ <= r_n_337__9_;
      r_337__8_ <= r_n_337__8_;
      r_337__7_ <= r_n_337__7_;
      r_337__6_ <= r_n_337__6_;
      r_337__5_ <= r_n_337__5_;
      r_337__4_ <= r_n_337__4_;
      r_337__3_ <= r_n_337__3_;
      r_337__2_ <= r_n_337__2_;
      r_337__1_ <= r_n_337__1_;
      r_337__0_ <= r_n_337__0_;
    end 
    if(N3922) begin
      r_338__63_ <= r_n_338__63_;
      r_338__62_ <= r_n_338__62_;
      r_338__61_ <= r_n_338__61_;
      r_338__60_ <= r_n_338__60_;
      r_338__59_ <= r_n_338__59_;
      r_338__58_ <= r_n_338__58_;
      r_338__57_ <= r_n_338__57_;
      r_338__56_ <= r_n_338__56_;
      r_338__55_ <= r_n_338__55_;
      r_338__54_ <= r_n_338__54_;
      r_338__53_ <= r_n_338__53_;
      r_338__52_ <= r_n_338__52_;
      r_338__51_ <= r_n_338__51_;
      r_338__50_ <= r_n_338__50_;
      r_338__49_ <= r_n_338__49_;
      r_338__48_ <= r_n_338__48_;
      r_338__47_ <= r_n_338__47_;
      r_338__46_ <= r_n_338__46_;
      r_338__45_ <= r_n_338__45_;
      r_338__44_ <= r_n_338__44_;
      r_338__43_ <= r_n_338__43_;
      r_338__42_ <= r_n_338__42_;
      r_338__41_ <= r_n_338__41_;
      r_338__40_ <= r_n_338__40_;
      r_338__39_ <= r_n_338__39_;
      r_338__38_ <= r_n_338__38_;
      r_338__37_ <= r_n_338__37_;
      r_338__36_ <= r_n_338__36_;
      r_338__35_ <= r_n_338__35_;
      r_338__34_ <= r_n_338__34_;
      r_338__33_ <= r_n_338__33_;
      r_338__32_ <= r_n_338__32_;
      r_338__31_ <= r_n_338__31_;
      r_338__30_ <= r_n_338__30_;
      r_338__29_ <= r_n_338__29_;
      r_338__28_ <= r_n_338__28_;
      r_338__27_ <= r_n_338__27_;
      r_338__26_ <= r_n_338__26_;
      r_338__25_ <= r_n_338__25_;
      r_338__24_ <= r_n_338__24_;
      r_338__23_ <= r_n_338__23_;
      r_338__22_ <= r_n_338__22_;
      r_338__21_ <= r_n_338__21_;
      r_338__20_ <= r_n_338__20_;
      r_338__19_ <= r_n_338__19_;
      r_338__18_ <= r_n_338__18_;
      r_338__17_ <= r_n_338__17_;
      r_338__16_ <= r_n_338__16_;
      r_338__15_ <= r_n_338__15_;
      r_338__14_ <= r_n_338__14_;
      r_338__13_ <= r_n_338__13_;
      r_338__12_ <= r_n_338__12_;
      r_338__11_ <= r_n_338__11_;
      r_338__10_ <= r_n_338__10_;
      r_338__9_ <= r_n_338__9_;
      r_338__8_ <= r_n_338__8_;
      r_338__7_ <= r_n_338__7_;
      r_338__6_ <= r_n_338__6_;
      r_338__5_ <= r_n_338__5_;
      r_338__4_ <= r_n_338__4_;
      r_338__3_ <= r_n_338__3_;
      r_338__2_ <= r_n_338__2_;
      r_338__1_ <= r_n_338__1_;
      r_338__0_ <= r_n_338__0_;
    end 
    if(N3923) begin
      r_339__63_ <= r_n_339__63_;
      r_339__62_ <= r_n_339__62_;
      r_339__61_ <= r_n_339__61_;
      r_339__60_ <= r_n_339__60_;
      r_339__59_ <= r_n_339__59_;
      r_339__58_ <= r_n_339__58_;
      r_339__57_ <= r_n_339__57_;
      r_339__56_ <= r_n_339__56_;
      r_339__55_ <= r_n_339__55_;
      r_339__54_ <= r_n_339__54_;
      r_339__53_ <= r_n_339__53_;
      r_339__52_ <= r_n_339__52_;
      r_339__51_ <= r_n_339__51_;
      r_339__50_ <= r_n_339__50_;
      r_339__49_ <= r_n_339__49_;
      r_339__48_ <= r_n_339__48_;
      r_339__47_ <= r_n_339__47_;
      r_339__46_ <= r_n_339__46_;
      r_339__45_ <= r_n_339__45_;
      r_339__44_ <= r_n_339__44_;
      r_339__43_ <= r_n_339__43_;
      r_339__42_ <= r_n_339__42_;
      r_339__41_ <= r_n_339__41_;
      r_339__40_ <= r_n_339__40_;
      r_339__39_ <= r_n_339__39_;
      r_339__38_ <= r_n_339__38_;
      r_339__37_ <= r_n_339__37_;
      r_339__36_ <= r_n_339__36_;
      r_339__35_ <= r_n_339__35_;
      r_339__34_ <= r_n_339__34_;
      r_339__33_ <= r_n_339__33_;
      r_339__32_ <= r_n_339__32_;
      r_339__31_ <= r_n_339__31_;
      r_339__30_ <= r_n_339__30_;
      r_339__29_ <= r_n_339__29_;
      r_339__28_ <= r_n_339__28_;
      r_339__27_ <= r_n_339__27_;
      r_339__26_ <= r_n_339__26_;
      r_339__25_ <= r_n_339__25_;
      r_339__24_ <= r_n_339__24_;
      r_339__23_ <= r_n_339__23_;
      r_339__22_ <= r_n_339__22_;
      r_339__21_ <= r_n_339__21_;
      r_339__20_ <= r_n_339__20_;
      r_339__19_ <= r_n_339__19_;
      r_339__18_ <= r_n_339__18_;
      r_339__17_ <= r_n_339__17_;
      r_339__16_ <= r_n_339__16_;
      r_339__15_ <= r_n_339__15_;
      r_339__14_ <= r_n_339__14_;
      r_339__13_ <= r_n_339__13_;
      r_339__12_ <= r_n_339__12_;
      r_339__11_ <= r_n_339__11_;
      r_339__10_ <= r_n_339__10_;
      r_339__9_ <= r_n_339__9_;
      r_339__8_ <= r_n_339__8_;
      r_339__7_ <= r_n_339__7_;
      r_339__6_ <= r_n_339__6_;
      r_339__5_ <= r_n_339__5_;
      r_339__4_ <= r_n_339__4_;
      r_339__3_ <= r_n_339__3_;
      r_339__2_ <= r_n_339__2_;
      r_339__1_ <= r_n_339__1_;
      r_339__0_ <= r_n_339__0_;
    end 
    if(N3924) begin
      r_340__63_ <= r_n_340__63_;
      r_340__62_ <= r_n_340__62_;
      r_340__61_ <= r_n_340__61_;
      r_340__60_ <= r_n_340__60_;
      r_340__59_ <= r_n_340__59_;
      r_340__58_ <= r_n_340__58_;
      r_340__57_ <= r_n_340__57_;
      r_340__56_ <= r_n_340__56_;
      r_340__55_ <= r_n_340__55_;
      r_340__54_ <= r_n_340__54_;
      r_340__53_ <= r_n_340__53_;
      r_340__52_ <= r_n_340__52_;
      r_340__51_ <= r_n_340__51_;
      r_340__50_ <= r_n_340__50_;
      r_340__49_ <= r_n_340__49_;
      r_340__48_ <= r_n_340__48_;
      r_340__47_ <= r_n_340__47_;
      r_340__46_ <= r_n_340__46_;
      r_340__45_ <= r_n_340__45_;
      r_340__44_ <= r_n_340__44_;
      r_340__43_ <= r_n_340__43_;
      r_340__42_ <= r_n_340__42_;
      r_340__41_ <= r_n_340__41_;
      r_340__40_ <= r_n_340__40_;
      r_340__39_ <= r_n_340__39_;
      r_340__38_ <= r_n_340__38_;
      r_340__37_ <= r_n_340__37_;
      r_340__36_ <= r_n_340__36_;
      r_340__35_ <= r_n_340__35_;
      r_340__34_ <= r_n_340__34_;
      r_340__33_ <= r_n_340__33_;
      r_340__32_ <= r_n_340__32_;
      r_340__31_ <= r_n_340__31_;
      r_340__30_ <= r_n_340__30_;
      r_340__29_ <= r_n_340__29_;
      r_340__28_ <= r_n_340__28_;
      r_340__27_ <= r_n_340__27_;
      r_340__26_ <= r_n_340__26_;
      r_340__25_ <= r_n_340__25_;
      r_340__24_ <= r_n_340__24_;
      r_340__23_ <= r_n_340__23_;
      r_340__22_ <= r_n_340__22_;
      r_340__21_ <= r_n_340__21_;
      r_340__20_ <= r_n_340__20_;
      r_340__19_ <= r_n_340__19_;
      r_340__18_ <= r_n_340__18_;
      r_340__17_ <= r_n_340__17_;
      r_340__16_ <= r_n_340__16_;
      r_340__15_ <= r_n_340__15_;
      r_340__14_ <= r_n_340__14_;
      r_340__13_ <= r_n_340__13_;
      r_340__12_ <= r_n_340__12_;
      r_340__11_ <= r_n_340__11_;
      r_340__10_ <= r_n_340__10_;
      r_340__9_ <= r_n_340__9_;
      r_340__8_ <= r_n_340__8_;
      r_340__7_ <= r_n_340__7_;
      r_340__6_ <= r_n_340__6_;
      r_340__5_ <= r_n_340__5_;
      r_340__4_ <= r_n_340__4_;
      r_340__3_ <= r_n_340__3_;
      r_340__2_ <= r_n_340__2_;
      r_340__1_ <= r_n_340__1_;
      r_340__0_ <= r_n_340__0_;
    end 
    if(N3925) begin
      r_341__63_ <= r_n_341__63_;
      r_341__62_ <= r_n_341__62_;
      r_341__61_ <= r_n_341__61_;
      r_341__60_ <= r_n_341__60_;
      r_341__59_ <= r_n_341__59_;
      r_341__58_ <= r_n_341__58_;
      r_341__57_ <= r_n_341__57_;
      r_341__56_ <= r_n_341__56_;
      r_341__55_ <= r_n_341__55_;
      r_341__54_ <= r_n_341__54_;
      r_341__53_ <= r_n_341__53_;
      r_341__52_ <= r_n_341__52_;
      r_341__51_ <= r_n_341__51_;
      r_341__50_ <= r_n_341__50_;
      r_341__49_ <= r_n_341__49_;
      r_341__48_ <= r_n_341__48_;
      r_341__47_ <= r_n_341__47_;
      r_341__46_ <= r_n_341__46_;
      r_341__45_ <= r_n_341__45_;
      r_341__44_ <= r_n_341__44_;
      r_341__43_ <= r_n_341__43_;
      r_341__42_ <= r_n_341__42_;
      r_341__41_ <= r_n_341__41_;
      r_341__40_ <= r_n_341__40_;
      r_341__39_ <= r_n_341__39_;
      r_341__38_ <= r_n_341__38_;
      r_341__37_ <= r_n_341__37_;
      r_341__36_ <= r_n_341__36_;
      r_341__35_ <= r_n_341__35_;
      r_341__34_ <= r_n_341__34_;
      r_341__33_ <= r_n_341__33_;
      r_341__32_ <= r_n_341__32_;
      r_341__31_ <= r_n_341__31_;
      r_341__30_ <= r_n_341__30_;
      r_341__29_ <= r_n_341__29_;
      r_341__28_ <= r_n_341__28_;
      r_341__27_ <= r_n_341__27_;
      r_341__26_ <= r_n_341__26_;
      r_341__25_ <= r_n_341__25_;
      r_341__24_ <= r_n_341__24_;
      r_341__23_ <= r_n_341__23_;
      r_341__22_ <= r_n_341__22_;
      r_341__21_ <= r_n_341__21_;
      r_341__20_ <= r_n_341__20_;
      r_341__19_ <= r_n_341__19_;
      r_341__18_ <= r_n_341__18_;
      r_341__17_ <= r_n_341__17_;
      r_341__16_ <= r_n_341__16_;
      r_341__15_ <= r_n_341__15_;
      r_341__14_ <= r_n_341__14_;
      r_341__13_ <= r_n_341__13_;
      r_341__12_ <= r_n_341__12_;
      r_341__11_ <= r_n_341__11_;
      r_341__10_ <= r_n_341__10_;
      r_341__9_ <= r_n_341__9_;
      r_341__8_ <= r_n_341__8_;
      r_341__7_ <= r_n_341__7_;
      r_341__6_ <= r_n_341__6_;
      r_341__5_ <= r_n_341__5_;
      r_341__4_ <= r_n_341__4_;
      r_341__3_ <= r_n_341__3_;
      r_341__2_ <= r_n_341__2_;
      r_341__1_ <= r_n_341__1_;
      r_341__0_ <= r_n_341__0_;
    end 
    if(N3926) begin
      r_342__63_ <= r_n_342__63_;
      r_342__62_ <= r_n_342__62_;
      r_342__61_ <= r_n_342__61_;
      r_342__60_ <= r_n_342__60_;
      r_342__59_ <= r_n_342__59_;
      r_342__58_ <= r_n_342__58_;
      r_342__57_ <= r_n_342__57_;
      r_342__56_ <= r_n_342__56_;
      r_342__55_ <= r_n_342__55_;
      r_342__54_ <= r_n_342__54_;
      r_342__53_ <= r_n_342__53_;
      r_342__52_ <= r_n_342__52_;
      r_342__51_ <= r_n_342__51_;
      r_342__50_ <= r_n_342__50_;
      r_342__49_ <= r_n_342__49_;
      r_342__48_ <= r_n_342__48_;
      r_342__47_ <= r_n_342__47_;
      r_342__46_ <= r_n_342__46_;
      r_342__45_ <= r_n_342__45_;
      r_342__44_ <= r_n_342__44_;
      r_342__43_ <= r_n_342__43_;
      r_342__42_ <= r_n_342__42_;
      r_342__41_ <= r_n_342__41_;
      r_342__40_ <= r_n_342__40_;
      r_342__39_ <= r_n_342__39_;
      r_342__38_ <= r_n_342__38_;
      r_342__37_ <= r_n_342__37_;
      r_342__36_ <= r_n_342__36_;
      r_342__35_ <= r_n_342__35_;
      r_342__34_ <= r_n_342__34_;
      r_342__33_ <= r_n_342__33_;
      r_342__32_ <= r_n_342__32_;
      r_342__31_ <= r_n_342__31_;
      r_342__30_ <= r_n_342__30_;
      r_342__29_ <= r_n_342__29_;
      r_342__28_ <= r_n_342__28_;
      r_342__27_ <= r_n_342__27_;
      r_342__26_ <= r_n_342__26_;
      r_342__25_ <= r_n_342__25_;
      r_342__24_ <= r_n_342__24_;
      r_342__23_ <= r_n_342__23_;
      r_342__22_ <= r_n_342__22_;
      r_342__21_ <= r_n_342__21_;
      r_342__20_ <= r_n_342__20_;
      r_342__19_ <= r_n_342__19_;
      r_342__18_ <= r_n_342__18_;
      r_342__17_ <= r_n_342__17_;
      r_342__16_ <= r_n_342__16_;
      r_342__15_ <= r_n_342__15_;
      r_342__14_ <= r_n_342__14_;
      r_342__13_ <= r_n_342__13_;
      r_342__12_ <= r_n_342__12_;
      r_342__11_ <= r_n_342__11_;
      r_342__10_ <= r_n_342__10_;
      r_342__9_ <= r_n_342__9_;
      r_342__8_ <= r_n_342__8_;
      r_342__7_ <= r_n_342__7_;
      r_342__6_ <= r_n_342__6_;
      r_342__5_ <= r_n_342__5_;
      r_342__4_ <= r_n_342__4_;
      r_342__3_ <= r_n_342__3_;
      r_342__2_ <= r_n_342__2_;
      r_342__1_ <= r_n_342__1_;
      r_342__0_ <= r_n_342__0_;
    end 
    if(N3927) begin
      r_343__63_ <= r_n_343__63_;
      r_343__62_ <= r_n_343__62_;
      r_343__61_ <= r_n_343__61_;
      r_343__60_ <= r_n_343__60_;
      r_343__59_ <= r_n_343__59_;
      r_343__58_ <= r_n_343__58_;
      r_343__57_ <= r_n_343__57_;
      r_343__56_ <= r_n_343__56_;
      r_343__55_ <= r_n_343__55_;
      r_343__54_ <= r_n_343__54_;
      r_343__53_ <= r_n_343__53_;
      r_343__52_ <= r_n_343__52_;
      r_343__51_ <= r_n_343__51_;
      r_343__50_ <= r_n_343__50_;
      r_343__49_ <= r_n_343__49_;
      r_343__48_ <= r_n_343__48_;
      r_343__47_ <= r_n_343__47_;
      r_343__46_ <= r_n_343__46_;
      r_343__45_ <= r_n_343__45_;
      r_343__44_ <= r_n_343__44_;
      r_343__43_ <= r_n_343__43_;
      r_343__42_ <= r_n_343__42_;
      r_343__41_ <= r_n_343__41_;
      r_343__40_ <= r_n_343__40_;
      r_343__39_ <= r_n_343__39_;
      r_343__38_ <= r_n_343__38_;
      r_343__37_ <= r_n_343__37_;
      r_343__36_ <= r_n_343__36_;
      r_343__35_ <= r_n_343__35_;
      r_343__34_ <= r_n_343__34_;
      r_343__33_ <= r_n_343__33_;
      r_343__32_ <= r_n_343__32_;
      r_343__31_ <= r_n_343__31_;
      r_343__30_ <= r_n_343__30_;
      r_343__29_ <= r_n_343__29_;
      r_343__28_ <= r_n_343__28_;
      r_343__27_ <= r_n_343__27_;
      r_343__26_ <= r_n_343__26_;
      r_343__25_ <= r_n_343__25_;
      r_343__24_ <= r_n_343__24_;
      r_343__23_ <= r_n_343__23_;
      r_343__22_ <= r_n_343__22_;
      r_343__21_ <= r_n_343__21_;
      r_343__20_ <= r_n_343__20_;
      r_343__19_ <= r_n_343__19_;
      r_343__18_ <= r_n_343__18_;
      r_343__17_ <= r_n_343__17_;
      r_343__16_ <= r_n_343__16_;
      r_343__15_ <= r_n_343__15_;
      r_343__14_ <= r_n_343__14_;
      r_343__13_ <= r_n_343__13_;
      r_343__12_ <= r_n_343__12_;
      r_343__11_ <= r_n_343__11_;
      r_343__10_ <= r_n_343__10_;
      r_343__9_ <= r_n_343__9_;
      r_343__8_ <= r_n_343__8_;
      r_343__7_ <= r_n_343__7_;
      r_343__6_ <= r_n_343__6_;
      r_343__5_ <= r_n_343__5_;
      r_343__4_ <= r_n_343__4_;
      r_343__3_ <= r_n_343__3_;
      r_343__2_ <= r_n_343__2_;
      r_343__1_ <= r_n_343__1_;
      r_343__0_ <= r_n_343__0_;
    end 
    if(N3928) begin
      r_344__63_ <= r_n_344__63_;
      r_344__62_ <= r_n_344__62_;
      r_344__61_ <= r_n_344__61_;
      r_344__60_ <= r_n_344__60_;
      r_344__59_ <= r_n_344__59_;
      r_344__58_ <= r_n_344__58_;
      r_344__57_ <= r_n_344__57_;
      r_344__56_ <= r_n_344__56_;
      r_344__55_ <= r_n_344__55_;
      r_344__54_ <= r_n_344__54_;
      r_344__53_ <= r_n_344__53_;
      r_344__52_ <= r_n_344__52_;
      r_344__51_ <= r_n_344__51_;
      r_344__50_ <= r_n_344__50_;
      r_344__49_ <= r_n_344__49_;
      r_344__48_ <= r_n_344__48_;
      r_344__47_ <= r_n_344__47_;
      r_344__46_ <= r_n_344__46_;
      r_344__45_ <= r_n_344__45_;
      r_344__44_ <= r_n_344__44_;
      r_344__43_ <= r_n_344__43_;
      r_344__42_ <= r_n_344__42_;
      r_344__41_ <= r_n_344__41_;
      r_344__40_ <= r_n_344__40_;
      r_344__39_ <= r_n_344__39_;
      r_344__38_ <= r_n_344__38_;
      r_344__37_ <= r_n_344__37_;
      r_344__36_ <= r_n_344__36_;
      r_344__35_ <= r_n_344__35_;
      r_344__34_ <= r_n_344__34_;
      r_344__33_ <= r_n_344__33_;
      r_344__32_ <= r_n_344__32_;
      r_344__31_ <= r_n_344__31_;
      r_344__30_ <= r_n_344__30_;
      r_344__29_ <= r_n_344__29_;
      r_344__28_ <= r_n_344__28_;
      r_344__27_ <= r_n_344__27_;
      r_344__26_ <= r_n_344__26_;
      r_344__25_ <= r_n_344__25_;
      r_344__24_ <= r_n_344__24_;
      r_344__23_ <= r_n_344__23_;
      r_344__22_ <= r_n_344__22_;
      r_344__21_ <= r_n_344__21_;
      r_344__20_ <= r_n_344__20_;
      r_344__19_ <= r_n_344__19_;
      r_344__18_ <= r_n_344__18_;
      r_344__17_ <= r_n_344__17_;
      r_344__16_ <= r_n_344__16_;
      r_344__15_ <= r_n_344__15_;
      r_344__14_ <= r_n_344__14_;
      r_344__13_ <= r_n_344__13_;
      r_344__12_ <= r_n_344__12_;
      r_344__11_ <= r_n_344__11_;
      r_344__10_ <= r_n_344__10_;
      r_344__9_ <= r_n_344__9_;
      r_344__8_ <= r_n_344__8_;
      r_344__7_ <= r_n_344__7_;
      r_344__6_ <= r_n_344__6_;
      r_344__5_ <= r_n_344__5_;
      r_344__4_ <= r_n_344__4_;
      r_344__3_ <= r_n_344__3_;
      r_344__2_ <= r_n_344__2_;
      r_344__1_ <= r_n_344__1_;
      r_344__0_ <= r_n_344__0_;
    end 
    if(N3929) begin
      r_345__63_ <= r_n_345__63_;
      r_345__62_ <= r_n_345__62_;
      r_345__61_ <= r_n_345__61_;
      r_345__60_ <= r_n_345__60_;
      r_345__59_ <= r_n_345__59_;
      r_345__58_ <= r_n_345__58_;
      r_345__57_ <= r_n_345__57_;
      r_345__56_ <= r_n_345__56_;
      r_345__55_ <= r_n_345__55_;
      r_345__54_ <= r_n_345__54_;
      r_345__53_ <= r_n_345__53_;
      r_345__52_ <= r_n_345__52_;
      r_345__51_ <= r_n_345__51_;
      r_345__50_ <= r_n_345__50_;
      r_345__49_ <= r_n_345__49_;
      r_345__48_ <= r_n_345__48_;
      r_345__47_ <= r_n_345__47_;
      r_345__46_ <= r_n_345__46_;
      r_345__45_ <= r_n_345__45_;
      r_345__44_ <= r_n_345__44_;
      r_345__43_ <= r_n_345__43_;
      r_345__42_ <= r_n_345__42_;
      r_345__41_ <= r_n_345__41_;
      r_345__40_ <= r_n_345__40_;
      r_345__39_ <= r_n_345__39_;
      r_345__38_ <= r_n_345__38_;
      r_345__37_ <= r_n_345__37_;
      r_345__36_ <= r_n_345__36_;
      r_345__35_ <= r_n_345__35_;
      r_345__34_ <= r_n_345__34_;
      r_345__33_ <= r_n_345__33_;
      r_345__32_ <= r_n_345__32_;
      r_345__31_ <= r_n_345__31_;
      r_345__30_ <= r_n_345__30_;
      r_345__29_ <= r_n_345__29_;
      r_345__28_ <= r_n_345__28_;
      r_345__27_ <= r_n_345__27_;
      r_345__26_ <= r_n_345__26_;
      r_345__25_ <= r_n_345__25_;
      r_345__24_ <= r_n_345__24_;
      r_345__23_ <= r_n_345__23_;
      r_345__22_ <= r_n_345__22_;
      r_345__21_ <= r_n_345__21_;
      r_345__20_ <= r_n_345__20_;
      r_345__19_ <= r_n_345__19_;
      r_345__18_ <= r_n_345__18_;
      r_345__17_ <= r_n_345__17_;
      r_345__16_ <= r_n_345__16_;
      r_345__15_ <= r_n_345__15_;
      r_345__14_ <= r_n_345__14_;
      r_345__13_ <= r_n_345__13_;
      r_345__12_ <= r_n_345__12_;
      r_345__11_ <= r_n_345__11_;
      r_345__10_ <= r_n_345__10_;
      r_345__9_ <= r_n_345__9_;
      r_345__8_ <= r_n_345__8_;
      r_345__7_ <= r_n_345__7_;
      r_345__6_ <= r_n_345__6_;
      r_345__5_ <= r_n_345__5_;
      r_345__4_ <= r_n_345__4_;
      r_345__3_ <= r_n_345__3_;
      r_345__2_ <= r_n_345__2_;
      r_345__1_ <= r_n_345__1_;
      r_345__0_ <= r_n_345__0_;
    end 
    if(N3930) begin
      r_346__63_ <= r_n_346__63_;
      r_346__62_ <= r_n_346__62_;
      r_346__61_ <= r_n_346__61_;
      r_346__60_ <= r_n_346__60_;
      r_346__59_ <= r_n_346__59_;
      r_346__58_ <= r_n_346__58_;
      r_346__57_ <= r_n_346__57_;
      r_346__56_ <= r_n_346__56_;
      r_346__55_ <= r_n_346__55_;
      r_346__54_ <= r_n_346__54_;
      r_346__53_ <= r_n_346__53_;
      r_346__52_ <= r_n_346__52_;
      r_346__51_ <= r_n_346__51_;
      r_346__50_ <= r_n_346__50_;
      r_346__49_ <= r_n_346__49_;
      r_346__48_ <= r_n_346__48_;
      r_346__47_ <= r_n_346__47_;
      r_346__46_ <= r_n_346__46_;
      r_346__45_ <= r_n_346__45_;
      r_346__44_ <= r_n_346__44_;
      r_346__43_ <= r_n_346__43_;
      r_346__42_ <= r_n_346__42_;
      r_346__41_ <= r_n_346__41_;
      r_346__40_ <= r_n_346__40_;
      r_346__39_ <= r_n_346__39_;
      r_346__38_ <= r_n_346__38_;
      r_346__37_ <= r_n_346__37_;
      r_346__36_ <= r_n_346__36_;
      r_346__35_ <= r_n_346__35_;
      r_346__34_ <= r_n_346__34_;
      r_346__33_ <= r_n_346__33_;
      r_346__32_ <= r_n_346__32_;
      r_346__31_ <= r_n_346__31_;
      r_346__30_ <= r_n_346__30_;
      r_346__29_ <= r_n_346__29_;
      r_346__28_ <= r_n_346__28_;
      r_346__27_ <= r_n_346__27_;
      r_346__26_ <= r_n_346__26_;
      r_346__25_ <= r_n_346__25_;
      r_346__24_ <= r_n_346__24_;
      r_346__23_ <= r_n_346__23_;
      r_346__22_ <= r_n_346__22_;
      r_346__21_ <= r_n_346__21_;
      r_346__20_ <= r_n_346__20_;
      r_346__19_ <= r_n_346__19_;
      r_346__18_ <= r_n_346__18_;
      r_346__17_ <= r_n_346__17_;
      r_346__16_ <= r_n_346__16_;
      r_346__15_ <= r_n_346__15_;
      r_346__14_ <= r_n_346__14_;
      r_346__13_ <= r_n_346__13_;
      r_346__12_ <= r_n_346__12_;
      r_346__11_ <= r_n_346__11_;
      r_346__10_ <= r_n_346__10_;
      r_346__9_ <= r_n_346__9_;
      r_346__8_ <= r_n_346__8_;
      r_346__7_ <= r_n_346__7_;
      r_346__6_ <= r_n_346__6_;
      r_346__5_ <= r_n_346__5_;
      r_346__4_ <= r_n_346__4_;
      r_346__3_ <= r_n_346__3_;
      r_346__2_ <= r_n_346__2_;
      r_346__1_ <= r_n_346__1_;
      r_346__0_ <= r_n_346__0_;
    end 
    if(N3931) begin
      r_347__63_ <= r_n_347__63_;
      r_347__62_ <= r_n_347__62_;
      r_347__61_ <= r_n_347__61_;
      r_347__60_ <= r_n_347__60_;
      r_347__59_ <= r_n_347__59_;
      r_347__58_ <= r_n_347__58_;
      r_347__57_ <= r_n_347__57_;
      r_347__56_ <= r_n_347__56_;
      r_347__55_ <= r_n_347__55_;
      r_347__54_ <= r_n_347__54_;
      r_347__53_ <= r_n_347__53_;
      r_347__52_ <= r_n_347__52_;
      r_347__51_ <= r_n_347__51_;
      r_347__50_ <= r_n_347__50_;
      r_347__49_ <= r_n_347__49_;
      r_347__48_ <= r_n_347__48_;
      r_347__47_ <= r_n_347__47_;
      r_347__46_ <= r_n_347__46_;
      r_347__45_ <= r_n_347__45_;
      r_347__44_ <= r_n_347__44_;
      r_347__43_ <= r_n_347__43_;
      r_347__42_ <= r_n_347__42_;
      r_347__41_ <= r_n_347__41_;
      r_347__40_ <= r_n_347__40_;
      r_347__39_ <= r_n_347__39_;
      r_347__38_ <= r_n_347__38_;
      r_347__37_ <= r_n_347__37_;
      r_347__36_ <= r_n_347__36_;
      r_347__35_ <= r_n_347__35_;
      r_347__34_ <= r_n_347__34_;
      r_347__33_ <= r_n_347__33_;
      r_347__32_ <= r_n_347__32_;
      r_347__31_ <= r_n_347__31_;
      r_347__30_ <= r_n_347__30_;
      r_347__29_ <= r_n_347__29_;
      r_347__28_ <= r_n_347__28_;
      r_347__27_ <= r_n_347__27_;
      r_347__26_ <= r_n_347__26_;
      r_347__25_ <= r_n_347__25_;
      r_347__24_ <= r_n_347__24_;
      r_347__23_ <= r_n_347__23_;
      r_347__22_ <= r_n_347__22_;
      r_347__21_ <= r_n_347__21_;
      r_347__20_ <= r_n_347__20_;
      r_347__19_ <= r_n_347__19_;
      r_347__18_ <= r_n_347__18_;
      r_347__17_ <= r_n_347__17_;
      r_347__16_ <= r_n_347__16_;
      r_347__15_ <= r_n_347__15_;
      r_347__14_ <= r_n_347__14_;
      r_347__13_ <= r_n_347__13_;
      r_347__12_ <= r_n_347__12_;
      r_347__11_ <= r_n_347__11_;
      r_347__10_ <= r_n_347__10_;
      r_347__9_ <= r_n_347__9_;
      r_347__8_ <= r_n_347__8_;
      r_347__7_ <= r_n_347__7_;
      r_347__6_ <= r_n_347__6_;
      r_347__5_ <= r_n_347__5_;
      r_347__4_ <= r_n_347__4_;
      r_347__3_ <= r_n_347__3_;
      r_347__2_ <= r_n_347__2_;
      r_347__1_ <= r_n_347__1_;
      r_347__0_ <= r_n_347__0_;
    end 
    if(N3932) begin
      r_348__63_ <= r_n_348__63_;
      r_348__62_ <= r_n_348__62_;
      r_348__61_ <= r_n_348__61_;
      r_348__60_ <= r_n_348__60_;
      r_348__59_ <= r_n_348__59_;
      r_348__58_ <= r_n_348__58_;
      r_348__57_ <= r_n_348__57_;
      r_348__56_ <= r_n_348__56_;
      r_348__55_ <= r_n_348__55_;
      r_348__54_ <= r_n_348__54_;
      r_348__53_ <= r_n_348__53_;
      r_348__52_ <= r_n_348__52_;
      r_348__51_ <= r_n_348__51_;
      r_348__50_ <= r_n_348__50_;
      r_348__49_ <= r_n_348__49_;
      r_348__48_ <= r_n_348__48_;
      r_348__47_ <= r_n_348__47_;
      r_348__46_ <= r_n_348__46_;
      r_348__45_ <= r_n_348__45_;
      r_348__44_ <= r_n_348__44_;
      r_348__43_ <= r_n_348__43_;
      r_348__42_ <= r_n_348__42_;
      r_348__41_ <= r_n_348__41_;
      r_348__40_ <= r_n_348__40_;
      r_348__39_ <= r_n_348__39_;
      r_348__38_ <= r_n_348__38_;
      r_348__37_ <= r_n_348__37_;
      r_348__36_ <= r_n_348__36_;
      r_348__35_ <= r_n_348__35_;
      r_348__34_ <= r_n_348__34_;
      r_348__33_ <= r_n_348__33_;
      r_348__32_ <= r_n_348__32_;
      r_348__31_ <= r_n_348__31_;
      r_348__30_ <= r_n_348__30_;
      r_348__29_ <= r_n_348__29_;
      r_348__28_ <= r_n_348__28_;
      r_348__27_ <= r_n_348__27_;
      r_348__26_ <= r_n_348__26_;
      r_348__25_ <= r_n_348__25_;
      r_348__24_ <= r_n_348__24_;
      r_348__23_ <= r_n_348__23_;
      r_348__22_ <= r_n_348__22_;
      r_348__21_ <= r_n_348__21_;
      r_348__20_ <= r_n_348__20_;
      r_348__19_ <= r_n_348__19_;
      r_348__18_ <= r_n_348__18_;
      r_348__17_ <= r_n_348__17_;
      r_348__16_ <= r_n_348__16_;
      r_348__15_ <= r_n_348__15_;
      r_348__14_ <= r_n_348__14_;
      r_348__13_ <= r_n_348__13_;
      r_348__12_ <= r_n_348__12_;
      r_348__11_ <= r_n_348__11_;
      r_348__10_ <= r_n_348__10_;
      r_348__9_ <= r_n_348__9_;
      r_348__8_ <= r_n_348__8_;
      r_348__7_ <= r_n_348__7_;
      r_348__6_ <= r_n_348__6_;
      r_348__5_ <= r_n_348__5_;
      r_348__4_ <= r_n_348__4_;
      r_348__3_ <= r_n_348__3_;
      r_348__2_ <= r_n_348__2_;
      r_348__1_ <= r_n_348__1_;
      r_348__0_ <= r_n_348__0_;
    end 
    if(N3933) begin
      r_349__63_ <= r_n_349__63_;
      r_349__62_ <= r_n_349__62_;
      r_349__61_ <= r_n_349__61_;
      r_349__60_ <= r_n_349__60_;
      r_349__59_ <= r_n_349__59_;
      r_349__58_ <= r_n_349__58_;
      r_349__57_ <= r_n_349__57_;
      r_349__56_ <= r_n_349__56_;
      r_349__55_ <= r_n_349__55_;
      r_349__54_ <= r_n_349__54_;
      r_349__53_ <= r_n_349__53_;
      r_349__52_ <= r_n_349__52_;
      r_349__51_ <= r_n_349__51_;
      r_349__50_ <= r_n_349__50_;
      r_349__49_ <= r_n_349__49_;
      r_349__48_ <= r_n_349__48_;
      r_349__47_ <= r_n_349__47_;
      r_349__46_ <= r_n_349__46_;
      r_349__45_ <= r_n_349__45_;
      r_349__44_ <= r_n_349__44_;
      r_349__43_ <= r_n_349__43_;
      r_349__42_ <= r_n_349__42_;
      r_349__41_ <= r_n_349__41_;
      r_349__40_ <= r_n_349__40_;
      r_349__39_ <= r_n_349__39_;
      r_349__38_ <= r_n_349__38_;
      r_349__37_ <= r_n_349__37_;
      r_349__36_ <= r_n_349__36_;
      r_349__35_ <= r_n_349__35_;
      r_349__34_ <= r_n_349__34_;
      r_349__33_ <= r_n_349__33_;
      r_349__32_ <= r_n_349__32_;
      r_349__31_ <= r_n_349__31_;
      r_349__30_ <= r_n_349__30_;
      r_349__29_ <= r_n_349__29_;
      r_349__28_ <= r_n_349__28_;
      r_349__27_ <= r_n_349__27_;
      r_349__26_ <= r_n_349__26_;
      r_349__25_ <= r_n_349__25_;
      r_349__24_ <= r_n_349__24_;
      r_349__23_ <= r_n_349__23_;
      r_349__22_ <= r_n_349__22_;
      r_349__21_ <= r_n_349__21_;
      r_349__20_ <= r_n_349__20_;
      r_349__19_ <= r_n_349__19_;
      r_349__18_ <= r_n_349__18_;
      r_349__17_ <= r_n_349__17_;
      r_349__16_ <= r_n_349__16_;
      r_349__15_ <= r_n_349__15_;
      r_349__14_ <= r_n_349__14_;
      r_349__13_ <= r_n_349__13_;
      r_349__12_ <= r_n_349__12_;
      r_349__11_ <= r_n_349__11_;
      r_349__10_ <= r_n_349__10_;
      r_349__9_ <= r_n_349__9_;
      r_349__8_ <= r_n_349__8_;
      r_349__7_ <= r_n_349__7_;
      r_349__6_ <= r_n_349__6_;
      r_349__5_ <= r_n_349__5_;
      r_349__4_ <= r_n_349__4_;
      r_349__3_ <= r_n_349__3_;
      r_349__2_ <= r_n_349__2_;
      r_349__1_ <= r_n_349__1_;
      r_349__0_ <= r_n_349__0_;
    end 
    if(N3934) begin
      r_350__63_ <= r_n_350__63_;
      r_350__62_ <= r_n_350__62_;
      r_350__61_ <= r_n_350__61_;
      r_350__60_ <= r_n_350__60_;
      r_350__59_ <= r_n_350__59_;
      r_350__58_ <= r_n_350__58_;
      r_350__57_ <= r_n_350__57_;
      r_350__56_ <= r_n_350__56_;
      r_350__55_ <= r_n_350__55_;
      r_350__54_ <= r_n_350__54_;
      r_350__53_ <= r_n_350__53_;
      r_350__52_ <= r_n_350__52_;
      r_350__51_ <= r_n_350__51_;
      r_350__50_ <= r_n_350__50_;
      r_350__49_ <= r_n_350__49_;
      r_350__48_ <= r_n_350__48_;
      r_350__47_ <= r_n_350__47_;
      r_350__46_ <= r_n_350__46_;
      r_350__45_ <= r_n_350__45_;
      r_350__44_ <= r_n_350__44_;
      r_350__43_ <= r_n_350__43_;
      r_350__42_ <= r_n_350__42_;
      r_350__41_ <= r_n_350__41_;
      r_350__40_ <= r_n_350__40_;
      r_350__39_ <= r_n_350__39_;
      r_350__38_ <= r_n_350__38_;
      r_350__37_ <= r_n_350__37_;
      r_350__36_ <= r_n_350__36_;
      r_350__35_ <= r_n_350__35_;
      r_350__34_ <= r_n_350__34_;
      r_350__33_ <= r_n_350__33_;
      r_350__32_ <= r_n_350__32_;
      r_350__31_ <= r_n_350__31_;
      r_350__30_ <= r_n_350__30_;
      r_350__29_ <= r_n_350__29_;
      r_350__28_ <= r_n_350__28_;
      r_350__27_ <= r_n_350__27_;
      r_350__26_ <= r_n_350__26_;
      r_350__25_ <= r_n_350__25_;
      r_350__24_ <= r_n_350__24_;
      r_350__23_ <= r_n_350__23_;
      r_350__22_ <= r_n_350__22_;
      r_350__21_ <= r_n_350__21_;
      r_350__20_ <= r_n_350__20_;
      r_350__19_ <= r_n_350__19_;
      r_350__18_ <= r_n_350__18_;
      r_350__17_ <= r_n_350__17_;
      r_350__16_ <= r_n_350__16_;
      r_350__15_ <= r_n_350__15_;
      r_350__14_ <= r_n_350__14_;
      r_350__13_ <= r_n_350__13_;
      r_350__12_ <= r_n_350__12_;
      r_350__11_ <= r_n_350__11_;
      r_350__10_ <= r_n_350__10_;
      r_350__9_ <= r_n_350__9_;
      r_350__8_ <= r_n_350__8_;
      r_350__7_ <= r_n_350__7_;
      r_350__6_ <= r_n_350__6_;
      r_350__5_ <= r_n_350__5_;
      r_350__4_ <= r_n_350__4_;
      r_350__3_ <= r_n_350__3_;
      r_350__2_ <= r_n_350__2_;
      r_350__1_ <= r_n_350__1_;
      r_350__0_ <= r_n_350__0_;
    end 
    if(N3935) begin
      r_351__63_ <= r_n_351__63_;
      r_351__62_ <= r_n_351__62_;
      r_351__61_ <= r_n_351__61_;
      r_351__60_ <= r_n_351__60_;
      r_351__59_ <= r_n_351__59_;
      r_351__58_ <= r_n_351__58_;
      r_351__57_ <= r_n_351__57_;
      r_351__56_ <= r_n_351__56_;
      r_351__55_ <= r_n_351__55_;
      r_351__54_ <= r_n_351__54_;
      r_351__53_ <= r_n_351__53_;
      r_351__52_ <= r_n_351__52_;
      r_351__51_ <= r_n_351__51_;
      r_351__50_ <= r_n_351__50_;
      r_351__49_ <= r_n_351__49_;
      r_351__48_ <= r_n_351__48_;
      r_351__47_ <= r_n_351__47_;
      r_351__46_ <= r_n_351__46_;
      r_351__45_ <= r_n_351__45_;
      r_351__44_ <= r_n_351__44_;
      r_351__43_ <= r_n_351__43_;
      r_351__42_ <= r_n_351__42_;
      r_351__41_ <= r_n_351__41_;
      r_351__40_ <= r_n_351__40_;
      r_351__39_ <= r_n_351__39_;
      r_351__38_ <= r_n_351__38_;
      r_351__37_ <= r_n_351__37_;
      r_351__36_ <= r_n_351__36_;
      r_351__35_ <= r_n_351__35_;
      r_351__34_ <= r_n_351__34_;
      r_351__33_ <= r_n_351__33_;
      r_351__32_ <= r_n_351__32_;
      r_351__31_ <= r_n_351__31_;
      r_351__30_ <= r_n_351__30_;
      r_351__29_ <= r_n_351__29_;
      r_351__28_ <= r_n_351__28_;
      r_351__27_ <= r_n_351__27_;
      r_351__26_ <= r_n_351__26_;
      r_351__25_ <= r_n_351__25_;
      r_351__24_ <= r_n_351__24_;
      r_351__23_ <= r_n_351__23_;
      r_351__22_ <= r_n_351__22_;
      r_351__21_ <= r_n_351__21_;
      r_351__20_ <= r_n_351__20_;
      r_351__19_ <= r_n_351__19_;
      r_351__18_ <= r_n_351__18_;
      r_351__17_ <= r_n_351__17_;
      r_351__16_ <= r_n_351__16_;
      r_351__15_ <= r_n_351__15_;
      r_351__14_ <= r_n_351__14_;
      r_351__13_ <= r_n_351__13_;
      r_351__12_ <= r_n_351__12_;
      r_351__11_ <= r_n_351__11_;
      r_351__10_ <= r_n_351__10_;
      r_351__9_ <= r_n_351__9_;
      r_351__8_ <= r_n_351__8_;
      r_351__7_ <= r_n_351__7_;
      r_351__6_ <= r_n_351__6_;
      r_351__5_ <= r_n_351__5_;
      r_351__4_ <= r_n_351__4_;
      r_351__3_ <= r_n_351__3_;
      r_351__2_ <= r_n_351__2_;
      r_351__1_ <= r_n_351__1_;
      r_351__0_ <= r_n_351__0_;
    end 
    if(N3936) begin
      r_352__63_ <= r_n_352__63_;
      r_352__62_ <= r_n_352__62_;
      r_352__61_ <= r_n_352__61_;
      r_352__60_ <= r_n_352__60_;
      r_352__59_ <= r_n_352__59_;
      r_352__58_ <= r_n_352__58_;
      r_352__57_ <= r_n_352__57_;
      r_352__56_ <= r_n_352__56_;
      r_352__55_ <= r_n_352__55_;
      r_352__54_ <= r_n_352__54_;
      r_352__53_ <= r_n_352__53_;
      r_352__52_ <= r_n_352__52_;
      r_352__51_ <= r_n_352__51_;
      r_352__50_ <= r_n_352__50_;
      r_352__49_ <= r_n_352__49_;
      r_352__48_ <= r_n_352__48_;
      r_352__47_ <= r_n_352__47_;
      r_352__46_ <= r_n_352__46_;
      r_352__45_ <= r_n_352__45_;
      r_352__44_ <= r_n_352__44_;
      r_352__43_ <= r_n_352__43_;
      r_352__42_ <= r_n_352__42_;
      r_352__41_ <= r_n_352__41_;
      r_352__40_ <= r_n_352__40_;
      r_352__39_ <= r_n_352__39_;
      r_352__38_ <= r_n_352__38_;
      r_352__37_ <= r_n_352__37_;
      r_352__36_ <= r_n_352__36_;
      r_352__35_ <= r_n_352__35_;
      r_352__34_ <= r_n_352__34_;
      r_352__33_ <= r_n_352__33_;
      r_352__32_ <= r_n_352__32_;
      r_352__31_ <= r_n_352__31_;
      r_352__30_ <= r_n_352__30_;
      r_352__29_ <= r_n_352__29_;
      r_352__28_ <= r_n_352__28_;
      r_352__27_ <= r_n_352__27_;
      r_352__26_ <= r_n_352__26_;
      r_352__25_ <= r_n_352__25_;
      r_352__24_ <= r_n_352__24_;
      r_352__23_ <= r_n_352__23_;
      r_352__22_ <= r_n_352__22_;
      r_352__21_ <= r_n_352__21_;
      r_352__20_ <= r_n_352__20_;
      r_352__19_ <= r_n_352__19_;
      r_352__18_ <= r_n_352__18_;
      r_352__17_ <= r_n_352__17_;
      r_352__16_ <= r_n_352__16_;
      r_352__15_ <= r_n_352__15_;
      r_352__14_ <= r_n_352__14_;
      r_352__13_ <= r_n_352__13_;
      r_352__12_ <= r_n_352__12_;
      r_352__11_ <= r_n_352__11_;
      r_352__10_ <= r_n_352__10_;
      r_352__9_ <= r_n_352__9_;
      r_352__8_ <= r_n_352__8_;
      r_352__7_ <= r_n_352__7_;
      r_352__6_ <= r_n_352__6_;
      r_352__5_ <= r_n_352__5_;
      r_352__4_ <= r_n_352__4_;
      r_352__3_ <= r_n_352__3_;
      r_352__2_ <= r_n_352__2_;
      r_352__1_ <= r_n_352__1_;
      r_352__0_ <= r_n_352__0_;
    end 
    if(N3937) begin
      r_353__63_ <= r_n_353__63_;
      r_353__62_ <= r_n_353__62_;
      r_353__61_ <= r_n_353__61_;
      r_353__60_ <= r_n_353__60_;
      r_353__59_ <= r_n_353__59_;
      r_353__58_ <= r_n_353__58_;
      r_353__57_ <= r_n_353__57_;
      r_353__56_ <= r_n_353__56_;
      r_353__55_ <= r_n_353__55_;
      r_353__54_ <= r_n_353__54_;
      r_353__53_ <= r_n_353__53_;
      r_353__52_ <= r_n_353__52_;
      r_353__51_ <= r_n_353__51_;
      r_353__50_ <= r_n_353__50_;
      r_353__49_ <= r_n_353__49_;
      r_353__48_ <= r_n_353__48_;
      r_353__47_ <= r_n_353__47_;
      r_353__46_ <= r_n_353__46_;
      r_353__45_ <= r_n_353__45_;
      r_353__44_ <= r_n_353__44_;
      r_353__43_ <= r_n_353__43_;
      r_353__42_ <= r_n_353__42_;
      r_353__41_ <= r_n_353__41_;
      r_353__40_ <= r_n_353__40_;
      r_353__39_ <= r_n_353__39_;
      r_353__38_ <= r_n_353__38_;
      r_353__37_ <= r_n_353__37_;
      r_353__36_ <= r_n_353__36_;
      r_353__35_ <= r_n_353__35_;
      r_353__34_ <= r_n_353__34_;
      r_353__33_ <= r_n_353__33_;
      r_353__32_ <= r_n_353__32_;
      r_353__31_ <= r_n_353__31_;
      r_353__30_ <= r_n_353__30_;
      r_353__29_ <= r_n_353__29_;
      r_353__28_ <= r_n_353__28_;
      r_353__27_ <= r_n_353__27_;
      r_353__26_ <= r_n_353__26_;
      r_353__25_ <= r_n_353__25_;
      r_353__24_ <= r_n_353__24_;
      r_353__23_ <= r_n_353__23_;
      r_353__22_ <= r_n_353__22_;
      r_353__21_ <= r_n_353__21_;
      r_353__20_ <= r_n_353__20_;
      r_353__19_ <= r_n_353__19_;
      r_353__18_ <= r_n_353__18_;
      r_353__17_ <= r_n_353__17_;
      r_353__16_ <= r_n_353__16_;
      r_353__15_ <= r_n_353__15_;
      r_353__14_ <= r_n_353__14_;
      r_353__13_ <= r_n_353__13_;
      r_353__12_ <= r_n_353__12_;
      r_353__11_ <= r_n_353__11_;
      r_353__10_ <= r_n_353__10_;
      r_353__9_ <= r_n_353__9_;
      r_353__8_ <= r_n_353__8_;
      r_353__7_ <= r_n_353__7_;
      r_353__6_ <= r_n_353__6_;
      r_353__5_ <= r_n_353__5_;
      r_353__4_ <= r_n_353__4_;
      r_353__3_ <= r_n_353__3_;
      r_353__2_ <= r_n_353__2_;
      r_353__1_ <= r_n_353__1_;
      r_353__0_ <= r_n_353__0_;
    end 
    if(N3938) begin
      r_354__63_ <= r_n_354__63_;
      r_354__62_ <= r_n_354__62_;
      r_354__61_ <= r_n_354__61_;
      r_354__60_ <= r_n_354__60_;
      r_354__59_ <= r_n_354__59_;
      r_354__58_ <= r_n_354__58_;
      r_354__57_ <= r_n_354__57_;
      r_354__56_ <= r_n_354__56_;
      r_354__55_ <= r_n_354__55_;
      r_354__54_ <= r_n_354__54_;
      r_354__53_ <= r_n_354__53_;
      r_354__52_ <= r_n_354__52_;
      r_354__51_ <= r_n_354__51_;
      r_354__50_ <= r_n_354__50_;
      r_354__49_ <= r_n_354__49_;
      r_354__48_ <= r_n_354__48_;
      r_354__47_ <= r_n_354__47_;
      r_354__46_ <= r_n_354__46_;
      r_354__45_ <= r_n_354__45_;
      r_354__44_ <= r_n_354__44_;
      r_354__43_ <= r_n_354__43_;
      r_354__42_ <= r_n_354__42_;
      r_354__41_ <= r_n_354__41_;
      r_354__40_ <= r_n_354__40_;
      r_354__39_ <= r_n_354__39_;
      r_354__38_ <= r_n_354__38_;
      r_354__37_ <= r_n_354__37_;
      r_354__36_ <= r_n_354__36_;
      r_354__35_ <= r_n_354__35_;
      r_354__34_ <= r_n_354__34_;
      r_354__33_ <= r_n_354__33_;
      r_354__32_ <= r_n_354__32_;
      r_354__31_ <= r_n_354__31_;
      r_354__30_ <= r_n_354__30_;
      r_354__29_ <= r_n_354__29_;
      r_354__28_ <= r_n_354__28_;
      r_354__27_ <= r_n_354__27_;
      r_354__26_ <= r_n_354__26_;
      r_354__25_ <= r_n_354__25_;
      r_354__24_ <= r_n_354__24_;
      r_354__23_ <= r_n_354__23_;
      r_354__22_ <= r_n_354__22_;
      r_354__21_ <= r_n_354__21_;
      r_354__20_ <= r_n_354__20_;
      r_354__19_ <= r_n_354__19_;
      r_354__18_ <= r_n_354__18_;
      r_354__17_ <= r_n_354__17_;
      r_354__16_ <= r_n_354__16_;
      r_354__15_ <= r_n_354__15_;
      r_354__14_ <= r_n_354__14_;
      r_354__13_ <= r_n_354__13_;
      r_354__12_ <= r_n_354__12_;
      r_354__11_ <= r_n_354__11_;
      r_354__10_ <= r_n_354__10_;
      r_354__9_ <= r_n_354__9_;
      r_354__8_ <= r_n_354__8_;
      r_354__7_ <= r_n_354__7_;
      r_354__6_ <= r_n_354__6_;
      r_354__5_ <= r_n_354__5_;
      r_354__4_ <= r_n_354__4_;
      r_354__3_ <= r_n_354__3_;
      r_354__2_ <= r_n_354__2_;
      r_354__1_ <= r_n_354__1_;
      r_354__0_ <= r_n_354__0_;
    end 
    if(N3939) begin
      r_355__63_ <= r_n_355__63_;
      r_355__62_ <= r_n_355__62_;
      r_355__61_ <= r_n_355__61_;
      r_355__60_ <= r_n_355__60_;
      r_355__59_ <= r_n_355__59_;
      r_355__58_ <= r_n_355__58_;
      r_355__57_ <= r_n_355__57_;
      r_355__56_ <= r_n_355__56_;
      r_355__55_ <= r_n_355__55_;
      r_355__54_ <= r_n_355__54_;
      r_355__53_ <= r_n_355__53_;
      r_355__52_ <= r_n_355__52_;
      r_355__51_ <= r_n_355__51_;
      r_355__50_ <= r_n_355__50_;
      r_355__49_ <= r_n_355__49_;
      r_355__48_ <= r_n_355__48_;
      r_355__47_ <= r_n_355__47_;
      r_355__46_ <= r_n_355__46_;
      r_355__45_ <= r_n_355__45_;
      r_355__44_ <= r_n_355__44_;
      r_355__43_ <= r_n_355__43_;
      r_355__42_ <= r_n_355__42_;
      r_355__41_ <= r_n_355__41_;
      r_355__40_ <= r_n_355__40_;
      r_355__39_ <= r_n_355__39_;
      r_355__38_ <= r_n_355__38_;
      r_355__37_ <= r_n_355__37_;
      r_355__36_ <= r_n_355__36_;
      r_355__35_ <= r_n_355__35_;
      r_355__34_ <= r_n_355__34_;
      r_355__33_ <= r_n_355__33_;
      r_355__32_ <= r_n_355__32_;
      r_355__31_ <= r_n_355__31_;
      r_355__30_ <= r_n_355__30_;
      r_355__29_ <= r_n_355__29_;
      r_355__28_ <= r_n_355__28_;
      r_355__27_ <= r_n_355__27_;
      r_355__26_ <= r_n_355__26_;
      r_355__25_ <= r_n_355__25_;
      r_355__24_ <= r_n_355__24_;
      r_355__23_ <= r_n_355__23_;
      r_355__22_ <= r_n_355__22_;
      r_355__21_ <= r_n_355__21_;
      r_355__20_ <= r_n_355__20_;
      r_355__19_ <= r_n_355__19_;
      r_355__18_ <= r_n_355__18_;
      r_355__17_ <= r_n_355__17_;
      r_355__16_ <= r_n_355__16_;
      r_355__15_ <= r_n_355__15_;
      r_355__14_ <= r_n_355__14_;
      r_355__13_ <= r_n_355__13_;
      r_355__12_ <= r_n_355__12_;
      r_355__11_ <= r_n_355__11_;
      r_355__10_ <= r_n_355__10_;
      r_355__9_ <= r_n_355__9_;
      r_355__8_ <= r_n_355__8_;
      r_355__7_ <= r_n_355__7_;
      r_355__6_ <= r_n_355__6_;
      r_355__5_ <= r_n_355__5_;
      r_355__4_ <= r_n_355__4_;
      r_355__3_ <= r_n_355__3_;
      r_355__2_ <= r_n_355__2_;
      r_355__1_ <= r_n_355__1_;
      r_355__0_ <= r_n_355__0_;
    end 
    if(N3940) begin
      r_356__63_ <= r_n_356__63_;
      r_356__62_ <= r_n_356__62_;
      r_356__61_ <= r_n_356__61_;
      r_356__60_ <= r_n_356__60_;
      r_356__59_ <= r_n_356__59_;
      r_356__58_ <= r_n_356__58_;
      r_356__57_ <= r_n_356__57_;
      r_356__56_ <= r_n_356__56_;
      r_356__55_ <= r_n_356__55_;
      r_356__54_ <= r_n_356__54_;
      r_356__53_ <= r_n_356__53_;
      r_356__52_ <= r_n_356__52_;
      r_356__51_ <= r_n_356__51_;
      r_356__50_ <= r_n_356__50_;
      r_356__49_ <= r_n_356__49_;
      r_356__48_ <= r_n_356__48_;
      r_356__47_ <= r_n_356__47_;
      r_356__46_ <= r_n_356__46_;
      r_356__45_ <= r_n_356__45_;
      r_356__44_ <= r_n_356__44_;
      r_356__43_ <= r_n_356__43_;
      r_356__42_ <= r_n_356__42_;
      r_356__41_ <= r_n_356__41_;
      r_356__40_ <= r_n_356__40_;
      r_356__39_ <= r_n_356__39_;
      r_356__38_ <= r_n_356__38_;
      r_356__37_ <= r_n_356__37_;
      r_356__36_ <= r_n_356__36_;
      r_356__35_ <= r_n_356__35_;
      r_356__34_ <= r_n_356__34_;
      r_356__33_ <= r_n_356__33_;
      r_356__32_ <= r_n_356__32_;
      r_356__31_ <= r_n_356__31_;
      r_356__30_ <= r_n_356__30_;
      r_356__29_ <= r_n_356__29_;
      r_356__28_ <= r_n_356__28_;
      r_356__27_ <= r_n_356__27_;
      r_356__26_ <= r_n_356__26_;
      r_356__25_ <= r_n_356__25_;
      r_356__24_ <= r_n_356__24_;
      r_356__23_ <= r_n_356__23_;
      r_356__22_ <= r_n_356__22_;
      r_356__21_ <= r_n_356__21_;
      r_356__20_ <= r_n_356__20_;
      r_356__19_ <= r_n_356__19_;
      r_356__18_ <= r_n_356__18_;
      r_356__17_ <= r_n_356__17_;
      r_356__16_ <= r_n_356__16_;
      r_356__15_ <= r_n_356__15_;
      r_356__14_ <= r_n_356__14_;
      r_356__13_ <= r_n_356__13_;
      r_356__12_ <= r_n_356__12_;
      r_356__11_ <= r_n_356__11_;
      r_356__10_ <= r_n_356__10_;
      r_356__9_ <= r_n_356__9_;
      r_356__8_ <= r_n_356__8_;
      r_356__7_ <= r_n_356__7_;
      r_356__6_ <= r_n_356__6_;
      r_356__5_ <= r_n_356__5_;
      r_356__4_ <= r_n_356__4_;
      r_356__3_ <= r_n_356__3_;
      r_356__2_ <= r_n_356__2_;
      r_356__1_ <= r_n_356__1_;
      r_356__0_ <= r_n_356__0_;
    end 
    if(N3941) begin
      r_357__63_ <= r_n_357__63_;
      r_357__62_ <= r_n_357__62_;
      r_357__61_ <= r_n_357__61_;
      r_357__60_ <= r_n_357__60_;
      r_357__59_ <= r_n_357__59_;
      r_357__58_ <= r_n_357__58_;
      r_357__57_ <= r_n_357__57_;
      r_357__56_ <= r_n_357__56_;
      r_357__55_ <= r_n_357__55_;
      r_357__54_ <= r_n_357__54_;
      r_357__53_ <= r_n_357__53_;
      r_357__52_ <= r_n_357__52_;
      r_357__51_ <= r_n_357__51_;
      r_357__50_ <= r_n_357__50_;
      r_357__49_ <= r_n_357__49_;
      r_357__48_ <= r_n_357__48_;
      r_357__47_ <= r_n_357__47_;
      r_357__46_ <= r_n_357__46_;
      r_357__45_ <= r_n_357__45_;
      r_357__44_ <= r_n_357__44_;
      r_357__43_ <= r_n_357__43_;
      r_357__42_ <= r_n_357__42_;
      r_357__41_ <= r_n_357__41_;
      r_357__40_ <= r_n_357__40_;
      r_357__39_ <= r_n_357__39_;
      r_357__38_ <= r_n_357__38_;
      r_357__37_ <= r_n_357__37_;
      r_357__36_ <= r_n_357__36_;
      r_357__35_ <= r_n_357__35_;
      r_357__34_ <= r_n_357__34_;
      r_357__33_ <= r_n_357__33_;
      r_357__32_ <= r_n_357__32_;
      r_357__31_ <= r_n_357__31_;
      r_357__30_ <= r_n_357__30_;
      r_357__29_ <= r_n_357__29_;
      r_357__28_ <= r_n_357__28_;
      r_357__27_ <= r_n_357__27_;
      r_357__26_ <= r_n_357__26_;
      r_357__25_ <= r_n_357__25_;
      r_357__24_ <= r_n_357__24_;
      r_357__23_ <= r_n_357__23_;
      r_357__22_ <= r_n_357__22_;
      r_357__21_ <= r_n_357__21_;
      r_357__20_ <= r_n_357__20_;
      r_357__19_ <= r_n_357__19_;
      r_357__18_ <= r_n_357__18_;
      r_357__17_ <= r_n_357__17_;
      r_357__16_ <= r_n_357__16_;
      r_357__15_ <= r_n_357__15_;
      r_357__14_ <= r_n_357__14_;
      r_357__13_ <= r_n_357__13_;
      r_357__12_ <= r_n_357__12_;
      r_357__11_ <= r_n_357__11_;
      r_357__10_ <= r_n_357__10_;
      r_357__9_ <= r_n_357__9_;
      r_357__8_ <= r_n_357__8_;
      r_357__7_ <= r_n_357__7_;
      r_357__6_ <= r_n_357__6_;
      r_357__5_ <= r_n_357__5_;
      r_357__4_ <= r_n_357__4_;
      r_357__3_ <= r_n_357__3_;
      r_357__2_ <= r_n_357__2_;
      r_357__1_ <= r_n_357__1_;
      r_357__0_ <= r_n_357__0_;
    end 
    if(N3942) begin
      r_358__63_ <= r_n_358__63_;
      r_358__62_ <= r_n_358__62_;
      r_358__61_ <= r_n_358__61_;
      r_358__60_ <= r_n_358__60_;
      r_358__59_ <= r_n_358__59_;
      r_358__58_ <= r_n_358__58_;
      r_358__57_ <= r_n_358__57_;
      r_358__56_ <= r_n_358__56_;
      r_358__55_ <= r_n_358__55_;
      r_358__54_ <= r_n_358__54_;
      r_358__53_ <= r_n_358__53_;
      r_358__52_ <= r_n_358__52_;
      r_358__51_ <= r_n_358__51_;
      r_358__50_ <= r_n_358__50_;
      r_358__49_ <= r_n_358__49_;
      r_358__48_ <= r_n_358__48_;
      r_358__47_ <= r_n_358__47_;
      r_358__46_ <= r_n_358__46_;
      r_358__45_ <= r_n_358__45_;
      r_358__44_ <= r_n_358__44_;
      r_358__43_ <= r_n_358__43_;
      r_358__42_ <= r_n_358__42_;
      r_358__41_ <= r_n_358__41_;
      r_358__40_ <= r_n_358__40_;
      r_358__39_ <= r_n_358__39_;
      r_358__38_ <= r_n_358__38_;
      r_358__37_ <= r_n_358__37_;
      r_358__36_ <= r_n_358__36_;
      r_358__35_ <= r_n_358__35_;
      r_358__34_ <= r_n_358__34_;
      r_358__33_ <= r_n_358__33_;
      r_358__32_ <= r_n_358__32_;
      r_358__31_ <= r_n_358__31_;
      r_358__30_ <= r_n_358__30_;
      r_358__29_ <= r_n_358__29_;
      r_358__28_ <= r_n_358__28_;
      r_358__27_ <= r_n_358__27_;
      r_358__26_ <= r_n_358__26_;
      r_358__25_ <= r_n_358__25_;
      r_358__24_ <= r_n_358__24_;
      r_358__23_ <= r_n_358__23_;
      r_358__22_ <= r_n_358__22_;
      r_358__21_ <= r_n_358__21_;
      r_358__20_ <= r_n_358__20_;
      r_358__19_ <= r_n_358__19_;
      r_358__18_ <= r_n_358__18_;
      r_358__17_ <= r_n_358__17_;
      r_358__16_ <= r_n_358__16_;
      r_358__15_ <= r_n_358__15_;
      r_358__14_ <= r_n_358__14_;
      r_358__13_ <= r_n_358__13_;
      r_358__12_ <= r_n_358__12_;
      r_358__11_ <= r_n_358__11_;
      r_358__10_ <= r_n_358__10_;
      r_358__9_ <= r_n_358__9_;
      r_358__8_ <= r_n_358__8_;
      r_358__7_ <= r_n_358__7_;
      r_358__6_ <= r_n_358__6_;
      r_358__5_ <= r_n_358__5_;
      r_358__4_ <= r_n_358__4_;
      r_358__3_ <= r_n_358__3_;
      r_358__2_ <= r_n_358__2_;
      r_358__1_ <= r_n_358__1_;
      r_358__0_ <= r_n_358__0_;
    end 
    if(N3943) begin
      r_359__63_ <= r_n_359__63_;
      r_359__62_ <= r_n_359__62_;
      r_359__61_ <= r_n_359__61_;
      r_359__60_ <= r_n_359__60_;
      r_359__59_ <= r_n_359__59_;
      r_359__58_ <= r_n_359__58_;
      r_359__57_ <= r_n_359__57_;
      r_359__56_ <= r_n_359__56_;
      r_359__55_ <= r_n_359__55_;
      r_359__54_ <= r_n_359__54_;
      r_359__53_ <= r_n_359__53_;
      r_359__52_ <= r_n_359__52_;
      r_359__51_ <= r_n_359__51_;
      r_359__50_ <= r_n_359__50_;
      r_359__49_ <= r_n_359__49_;
      r_359__48_ <= r_n_359__48_;
      r_359__47_ <= r_n_359__47_;
      r_359__46_ <= r_n_359__46_;
      r_359__45_ <= r_n_359__45_;
      r_359__44_ <= r_n_359__44_;
      r_359__43_ <= r_n_359__43_;
      r_359__42_ <= r_n_359__42_;
      r_359__41_ <= r_n_359__41_;
      r_359__40_ <= r_n_359__40_;
      r_359__39_ <= r_n_359__39_;
      r_359__38_ <= r_n_359__38_;
      r_359__37_ <= r_n_359__37_;
      r_359__36_ <= r_n_359__36_;
      r_359__35_ <= r_n_359__35_;
      r_359__34_ <= r_n_359__34_;
      r_359__33_ <= r_n_359__33_;
      r_359__32_ <= r_n_359__32_;
      r_359__31_ <= r_n_359__31_;
      r_359__30_ <= r_n_359__30_;
      r_359__29_ <= r_n_359__29_;
      r_359__28_ <= r_n_359__28_;
      r_359__27_ <= r_n_359__27_;
      r_359__26_ <= r_n_359__26_;
      r_359__25_ <= r_n_359__25_;
      r_359__24_ <= r_n_359__24_;
      r_359__23_ <= r_n_359__23_;
      r_359__22_ <= r_n_359__22_;
      r_359__21_ <= r_n_359__21_;
      r_359__20_ <= r_n_359__20_;
      r_359__19_ <= r_n_359__19_;
      r_359__18_ <= r_n_359__18_;
      r_359__17_ <= r_n_359__17_;
      r_359__16_ <= r_n_359__16_;
      r_359__15_ <= r_n_359__15_;
      r_359__14_ <= r_n_359__14_;
      r_359__13_ <= r_n_359__13_;
      r_359__12_ <= r_n_359__12_;
      r_359__11_ <= r_n_359__11_;
      r_359__10_ <= r_n_359__10_;
      r_359__9_ <= r_n_359__9_;
      r_359__8_ <= r_n_359__8_;
      r_359__7_ <= r_n_359__7_;
      r_359__6_ <= r_n_359__6_;
      r_359__5_ <= r_n_359__5_;
      r_359__4_ <= r_n_359__4_;
      r_359__3_ <= r_n_359__3_;
      r_359__2_ <= r_n_359__2_;
      r_359__1_ <= r_n_359__1_;
      r_359__0_ <= r_n_359__0_;
    end 
    if(N3944) begin
      r_360__63_ <= r_n_360__63_;
      r_360__62_ <= r_n_360__62_;
      r_360__61_ <= r_n_360__61_;
      r_360__60_ <= r_n_360__60_;
      r_360__59_ <= r_n_360__59_;
      r_360__58_ <= r_n_360__58_;
      r_360__57_ <= r_n_360__57_;
      r_360__56_ <= r_n_360__56_;
      r_360__55_ <= r_n_360__55_;
      r_360__54_ <= r_n_360__54_;
      r_360__53_ <= r_n_360__53_;
      r_360__52_ <= r_n_360__52_;
      r_360__51_ <= r_n_360__51_;
      r_360__50_ <= r_n_360__50_;
      r_360__49_ <= r_n_360__49_;
      r_360__48_ <= r_n_360__48_;
      r_360__47_ <= r_n_360__47_;
      r_360__46_ <= r_n_360__46_;
      r_360__45_ <= r_n_360__45_;
      r_360__44_ <= r_n_360__44_;
      r_360__43_ <= r_n_360__43_;
      r_360__42_ <= r_n_360__42_;
      r_360__41_ <= r_n_360__41_;
      r_360__40_ <= r_n_360__40_;
      r_360__39_ <= r_n_360__39_;
      r_360__38_ <= r_n_360__38_;
      r_360__37_ <= r_n_360__37_;
      r_360__36_ <= r_n_360__36_;
      r_360__35_ <= r_n_360__35_;
      r_360__34_ <= r_n_360__34_;
      r_360__33_ <= r_n_360__33_;
      r_360__32_ <= r_n_360__32_;
      r_360__31_ <= r_n_360__31_;
      r_360__30_ <= r_n_360__30_;
      r_360__29_ <= r_n_360__29_;
      r_360__28_ <= r_n_360__28_;
      r_360__27_ <= r_n_360__27_;
      r_360__26_ <= r_n_360__26_;
      r_360__25_ <= r_n_360__25_;
      r_360__24_ <= r_n_360__24_;
      r_360__23_ <= r_n_360__23_;
      r_360__22_ <= r_n_360__22_;
      r_360__21_ <= r_n_360__21_;
      r_360__20_ <= r_n_360__20_;
      r_360__19_ <= r_n_360__19_;
      r_360__18_ <= r_n_360__18_;
      r_360__17_ <= r_n_360__17_;
      r_360__16_ <= r_n_360__16_;
      r_360__15_ <= r_n_360__15_;
      r_360__14_ <= r_n_360__14_;
      r_360__13_ <= r_n_360__13_;
      r_360__12_ <= r_n_360__12_;
      r_360__11_ <= r_n_360__11_;
      r_360__10_ <= r_n_360__10_;
      r_360__9_ <= r_n_360__9_;
      r_360__8_ <= r_n_360__8_;
      r_360__7_ <= r_n_360__7_;
      r_360__6_ <= r_n_360__6_;
      r_360__5_ <= r_n_360__5_;
      r_360__4_ <= r_n_360__4_;
      r_360__3_ <= r_n_360__3_;
      r_360__2_ <= r_n_360__2_;
      r_360__1_ <= r_n_360__1_;
      r_360__0_ <= r_n_360__0_;
    end 
    if(N3945) begin
      r_361__63_ <= r_n_361__63_;
      r_361__62_ <= r_n_361__62_;
      r_361__61_ <= r_n_361__61_;
      r_361__60_ <= r_n_361__60_;
      r_361__59_ <= r_n_361__59_;
      r_361__58_ <= r_n_361__58_;
      r_361__57_ <= r_n_361__57_;
      r_361__56_ <= r_n_361__56_;
      r_361__55_ <= r_n_361__55_;
      r_361__54_ <= r_n_361__54_;
      r_361__53_ <= r_n_361__53_;
      r_361__52_ <= r_n_361__52_;
      r_361__51_ <= r_n_361__51_;
      r_361__50_ <= r_n_361__50_;
      r_361__49_ <= r_n_361__49_;
      r_361__48_ <= r_n_361__48_;
      r_361__47_ <= r_n_361__47_;
      r_361__46_ <= r_n_361__46_;
      r_361__45_ <= r_n_361__45_;
      r_361__44_ <= r_n_361__44_;
      r_361__43_ <= r_n_361__43_;
      r_361__42_ <= r_n_361__42_;
      r_361__41_ <= r_n_361__41_;
      r_361__40_ <= r_n_361__40_;
      r_361__39_ <= r_n_361__39_;
      r_361__38_ <= r_n_361__38_;
      r_361__37_ <= r_n_361__37_;
      r_361__36_ <= r_n_361__36_;
      r_361__35_ <= r_n_361__35_;
      r_361__34_ <= r_n_361__34_;
      r_361__33_ <= r_n_361__33_;
      r_361__32_ <= r_n_361__32_;
      r_361__31_ <= r_n_361__31_;
      r_361__30_ <= r_n_361__30_;
      r_361__29_ <= r_n_361__29_;
      r_361__28_ <= r_n_361__28_;
      r_361__27_ <= r_n_361__27_;
      r_361__26_ <= r_n_361__26_;
      r_361__25_ <= r_n_361__25_;
      r_361__24_ <= r_n_361__24_;
      r_361__23_ <= r_n_361__23_;
      r_361__22_ <= r_n_361__22_;
      r_361__21_ <= r_n_361__21_;
      r_361__20_ <= r_n_361__20_;
      r_361__19_ <= r_n_361__19_;
      r_361__18_ <= r_n_361__18_;
      r_361__17_ <= r_n_361__17_;
      r_361__16_ <= r_n_361__16_;
      r_361__15_ <= r_n_361__15_;
      r_361__14_ <= r_n_361__14_;
      r_361__13_ <= r_n_361__13_;
      r_361__12_ <= r_n_361__12_;
      r_361__11_ <= r_n_361__11_;
      r_361__10_ <= r_n_361__10_;
      r_361__9_ <= r_n_361__9_;
      r_361__8_ <= r_n_361__8_;
      r_361__7_ <= r_n_361__7_;
      r_361__6_ <= r_n_361__6_;
      r_361__5_ <= r_n_361__5_;
      r_361__4_ <= r_n_361__4_;
      r_361__3_ <= r_n_361__3_;
      r_361__2_ <= r_n_361__2_;
      r_361__1_ <= r_n_361__1_;
      r_361__0_ <= r_n_361__0_;
    end 
    if(N3946) begin
      r_362__63_ <= r_n_362__63_;
      r_362__62_ <= r_n_362__62_;
      r_362__61_ <= r_n_362__61_;
      r_362__60_ <= r_n_362__60_;
      r_362__59_ <= r_n_362__59_;
      r_362__58_ <= r_n_362__58_;
      r_362__57_ <= r_n_362__57_;
      r_362__56_ <= r_n_362__56_;
      r_362__55_ <= r_n_362__55_;
      r_362__54_ <= r_n_362__54_;
      r_362__53_ <= r_n_362__53_;
      r_362__52_ <= r_n_362__52_;
      r_362__51_ <= r_n_362__51_;
      r_362__50_ <= r_n_362__50_;
      r_362__49_ <= r_n_362__49_;
      r_362__48_ <= r_n_362__48_;
      r_362__47_ <= r_n_362__47_;
      r_362__46_ <= r_n_362__46_;
      r_362__45_ <= r_n_362__45_;
      r_362__44_ <= r_n_362__44_;
      r_362__43_ <= r_n_362__43_;
      r_362__42_ <= r_n_362__42_;
      r_362__41_ <= r_n_362__41_;
      r_362__40_ <= r_n_362__40_;
      r_362__39_ <= r_n_362__39_;
      r_362__38_ <= r_n_362__38_;
      r_362__37_ <= r_n_362__37_;
      r_362__36_ <= r_n_362__36_;
      r_362__35_ <= r_n_362__35_;
      r_362__34_ <= r_n_362__34_;
      r_362__33_ <= r_n_362__33_;
      r_362__32_ <= r_n_362__32_;
      r_362__31_ <= r_n_362__31_;
      r_362__30_ <= r_n_362__30_;
      r_362__29_ <= r_n_362__29_;
      r_362__28_ <= r_n_362__28_;
      r_362__27_ <= r_n_362__27_;
      r_362__26_ <= r_n_362__26_;
      r_362__25_ <= r_n_362__25_;
      r_362__24_ <= r_n_362__24_;
      r_362__23_ <= r_n_362__23_;
      r_362__22_ <= r_n_362__22_;
      r_362__21_ <= r_n_362__21_;
      r_362__20_ <= r_n_362__20_;
      r_362__19_ <= r_n_362__19_;
      r_362__18_ <= r_n_362__18_;
      r_362__17_ <= r_n_362__17_;
      r_362__16_ <= r_n_362__16_;
      r_362__15_ <= r_n_362__15_;
      r_362__14_ <= r_n_362__14_;
      r_362__13_ <= r_n_362__13_;
      r_362__12_ <= r_n_362__12_;
      r_362__11_ <= r_n_362__11_;
      r_362__10_ <= r_n_362__10_;
      r_362__9_ <= r_n_362__9_;
      r_362__8_ <= r_n_362__8_;
      r_362__7_ <= r_n_362__7_;
      r_362__6_ <= r_n_362__6_;
      r_362__5_ <= r_n_362__5_;
      r_362__4_ <= r_n_362__4_;
      r_362__3_ <= r_n_362__3_;
      r_362__2_ <= r_n_362__2_;
      r_362__1_ <= r_n_362__1_;
      r_362__0_ <= r_n_362__0_;
    end 
    if(N3947) begin
      r_363__63_ <= r_n_363__63_;
      r_363__62_ <= r_n_363__62_;
      r_363__61_ <= r_n_363__61_;
      r_363__60_ <= r_n_363__60_;
      r_363__59_ <= r_n_363__59_;
      r_363__58_ <= r_n_363__58_;
      r_363__57_ <= r_n_363__57_;
      r_363__56_ <= r_n_363__56_;
      r_363__55_ <= r_n_363__55_;
      r_363__54_ <= r_n_363__54_;
      r_363__53_ <= r_n_363__53_;
      r_363__52_ <= r_n_363__52_;
      r_363__51_ <= r_n_363__51_;
      r_363__50_ <= r_n_363__50_;
      r_363__49_ <= r_n_363__49_;
      r_363__48_ <= r_n_363__48_;
      r_363__47_ <= r_n_363__47_;
      r_363__46_ <= r_n_363__46_;
      r_363__45_ <= r_n_363__45_;
      r_363__44_ <= r_n_363__44_;
      r_363__43_ <= r_n_363__43_;
      r_363__42_ <= r_n_363__42_;
      r_363__41_ <= r_n_363__41_;
      r_363__40_ <= r_n_363__40_;
      r_363__39_ <= r_n_363__39_;
      r_363__38_ <= r_n_363__38_;
      r_363__37_ <= r_n_363__37_;
      r_363__36_ <= r_n_363__36_;
      r_363__35_ <= r_n_363__35_;
      r_363__34_ <= r_n_363__34_;
      r_363__33_ <= r_n_363__33_;
      r_363__32_ <= r_n_363__32_;
      r_363__31_ <= r_n_363__31_;
      r_363__30_ <= r_n_363__30_;
      r_363__29_ <= r_n_363__29_;
      r_363__28_ <= r_n_363__28_;
      r_363__27_ <= r_n_363__27_;
      r_363__26_ <= r_n_363__26_;
      r_363__25_ <= r_n_363__25_;
      r_363__24_ <= r_n_363__24_;
      r_363__23_ <= r_n_363__23_;
      r_363__22_ <= r_n_363__22_;
      r_363__21_ <= r_n_363__21_;
      r_363__20_ <= r_n_363__20_;
      r_363__19_ <= r_n_363__19_;
      r_363__18_ <= r_n_363__18_;
      r_363__17_ <= r_n_363__17_;
      r_363__16_ <= r_n_363__16_;
      r_363__15_ <= r_n_363__15_;
      r_363__14_ <= r_n_363__14_;
      r_363__13_ <= r_n_363__13_;
      r_363__12_ <= r_n_363__12_;
      r_363__11_ <= r_n_363__11_;
      r_363__10_ <= r_n_363__10_;
      r_363__9_ <= r_n_363__9_;
      r_363__8_ <= r_n_363__8_;
      r_363__7_ <= r_n_363__7_;
      r_363__6_ <= r_n_363__6_;
      r_363__5_ <= r_n_363__5_;
      r_363__4_ <= r_n_363__4_;
      r_363__3_ <= r_n_363__3_;
      r_363__2_ <= r_n_363__2_;
      r_363__1_ <= r_n_363__1_;
      r_363__0_ <= r_n_363__0_;
    end 
    if(N3948) begin
      r_364__63_ <= r_n_364__63_;
      r_364__62_ <= r_n_364__62_;
      r_364__61_ <= r_n_364__61_;
      r_364__60_ <= r_n_364__60_;
      r_364__59_ <= r_n_364__59_;
      r_364__58_ <= r_n_364__58_;
      r_364__57_ <= r_n_364__57_;
      r_364__56_ <= r_n_364__56_;
      r_364__55_ <= r_n_364__55_;
      r_364__54_ <= r_n_364__54_;
      r_364__53_ <= r_n_364__53_;
      r_364__52_ <= r_n_364__52_;
      r_364__51_ <= r_n_364__51_;
      r_364__50_ <= r_n_364__50_;
      r_364__49_ <= r_n_364__49_;
      r_364__48_ <= r_n_364__48_;
      r_364__47_ <= r_n_364__47_;
      r_364__46_ <= r_n_364__46_;
      r_364__45_ <= r_n_364__45_;
      r_364__44_ <= r_n_364__44_;
      r_364__43_ <= r_n_364__43_;
      r_364__42_ <= r_n_364__42_;
      r_364__41_ <= r_n_364__41_;
      r_364__40_ <= r_n_364__40_;
      r_364__39_ <= r_n_364__39_;
      r_364__38_ <= r_n_364__38_;
      r_364__37_ <= r_n_364__37_;
      r_364__36_ <= r_n_364__36_;
      r_364__35_ <= r_n_364__35_;
      r_364__34_ <= r_n_364__34_;
      r_364__33_ <= r_n_364__33_;
      r_364__32_ <= r_n_364__32_;
      r_364__31_ <= r_n_364__31_;
      r_364__30_ <= r_n_364__30_;
      r_364__29_ <= r_n_364__29_;
      r_364__28_ <= r_n_364__28_;
      r_364__27_ <= r_n_364__27_;
      r_364__26_ <= r_n_364__26_;
      r_364__25_ <= r_n_364__25_;
      r_364__24_ <= r_n_364__24_;
      r_364__23_ <= r_n_364__23_;
      r_364__22_ <= r_n_364__22_;
      r_364__21_ <= r_n_364__21_;
      r_364__20_ <= r_n_364__20_;
      r_364__19_ <= r_n_364__19_;
      r_364__18_ <= r_n_364__18_;
      r_364__17_ <= r_n_364__17_;
      r_364__16_ <= r_n_364__16_;
      r_364__15_ <= r_n_364__15_;
      r_364__14_ <= r_n_364__14_;
      r_364__13_ <= r_n_364__13_;
      r_364__12_ <= r_n_364__12_;
      r_364__11_ <= r_n_364__11_;
      r_364__10_ <= r_n_364__10_;
      r_364__9_ <= r_n_364__9_;
      r_364__8_ <= r_n_364__8_;
      r_364__7_ <= r_n_364__7_;
      r_364__6_ <= r_n_364__6_;
      r_364__5_ <= r_n_364__5_;
      r_364__4_ <= r_n_364__4_;
      r_364__3_ <= r_n_364__3_;
      r_364__2_ <= r_n_364__2_;
      r_364__1_ <= r_n_364__1_;
      r_364__0_ <= r_n_364__0_;
    end 
    if(N3949) begin
      r_365__63_ <= r_n_365__63_;
      r_365__62_ <= r_n_365__62_;
      r_365__61_ <= r_n_365__61_;
      r_365__60_ <= r_n_365__60_;
      r_365__59_ <= r_n_365__59_;
      r_365__58_ <= r_n_365__58_;
      r_365__57_ <= r_n_365__57_;
      r_365__56_ <= r_n_365__56_;
      r_365__55_ <= r_n_365__55_;
      r_365__54_ <= r_n_365__54_;
      r_365__53_ <= r_n_365__53_;
      r_365__52_ <= r_n_365__52_;
      r_365__51_ <= r_n_365__51_;
      r_365__50_ <= r_n_365__50_;
      r_365__49_ <= r_n_365__49_;
      r_365__48_ <= r_n_365__48_;
      r_365__47_ <= r_n_365__47_;
      r_365__46_ <= r_n_365__46_;
      r_365__45_ <= r_n_365__45_;
      r_365__44_ <= r_n_365__44_;
      r_365__43_ <= r_n_365__43_;
      r_365__42_ <= r_n_365__42_;
      r_365__41_ <= r_n_365__41_;
      r_365__40_ <= r_n_365__40_;
      r_365__39_ <= r_n_365__39_;
      r_365__38_ <= r_n_365__38_;
      r_365__37_ <= r_n_365__37_;
      r_365__36_ <= r_n_365__36_;
      r_365__35_ <= r_n_365__35_;
      r_365__34_ <= r_n_365__34_;
      r_365__33_ <= r_n_365__33_;
      r_365__32_ <= r_n_365__32_;
      r_365__31_ <= r_n_365__31_;
      r_365__30_ <= r_n_365__30_;
      r_365__29_ <= r_n_365__29_;
      r_365__28_ <= r_n_365__28_;
      r_365__27_ <= r_n_365__27_;
      r_365__26_ <= r_n_365__26_;
      r_365__25_ <= r_n_365__25_;
      r_365__24_ <= r_n_365__24_;
      r_365__23_ <= r_n_365__23_;
      r_365__22_ <= r_n_365__22_;
      r_365__21_ <= r_n_365__21_;
      r_365__20_ <= r_n_365__20_;
      r_365__19_ <= r_n_365__19_;
      r_365__18_ <= r_n_365__18_;
      r_365__17_ <= r_n_365__17_;
      r_365__16_ <= r_n_365__16_;
      r_365__15_ <= r_n_365__15_;
      r_365__14_ <= r_n_365__14_;
      r_365__13_ <= r_n_365__13_;
      r_365__12_ <= r_n_365__12_;
      r_365__11_ <= r_n_365__11_;
      r_365__10_ <= r_n_365__10_;
      r_365__9_ <= r_n_365__9_;
      r_365__8_ <= r_n_365__8_;
      r_365__7_ <= r_n_365__7_;
      r_365__6_ <= r_n_365__6_;
      r_365__5_ <= r_n_365__5_;
      r_365__4_ <= r_n_365__4_;
      r_365__3_ <= r_n_365__3_;
      r_365__2_ <= r_n_365__2_;
      r_365__1_ <= r_n_365__1_;
      r_365__0_ <= r_n_365__0_;
    end 
    if(N3950) begin
      r_366__63_ <= r_n_366__63_;
      r_366__62_ <= r_n_366__62_;
      r_366__61_ <= r_n_366__61_;
      r_366__60_ <= r_n_366__60_;
      r_366__59_ <= r_n_366__59_;
      r_366__58_ <= r_n_366__58_;
      r_366__57_ <= r_n_366__57_;
      r_366__56_ <= r_n_366__56_;
      r_366__55_ <= r_n_366__55_;
      r_366__54_ <= r_n_366__54_;
      r_366__53_ <= r_n_366__53_;
      r_366__52_ <= r_n_366__52_;
      r_366__51_ <= r_n_366__51_;
      r_366__50_ <= r_n_366__50_;
      r_366__49_ <= r_n_366__49_;
      r_366__48_ <= r_n_366__48_;
      r_366__47_ <= r_n_366__47_;
      r_366__46_ <= r_n_366__46_;
      r_366__45_ <= r_n_366__45_;
      r_366__44_ <= r_n_366__44_;
      r_366__43_ <= r_n_366__43_;
      r_366__42_ <= r_n_366__42_;
      r_366__41_ <= r_n_366__41_;
      r_366__40_ <= r_n_366__40_;
      r_366__39_ <= r_n_366__39_;
      r_366__38_ <= r_n_366__38_;
      r_366__37_ <= r_n_366__37_;
      r_366__36_ <= r_n_366__36_;
      r_366__35_ <= r_n_366__35_;
      r_366__34_ <= r_n_366__34_;
      r_366__33_ <= r_n_366__33_;
      r_366__32_ <= r_n_366__32_;
      r_366__31_ <= r_n_366__31_;
      r_366__30_ <= r_n_366__30_;
      r_366__29_ <= r_n_366__29_;
      r_366__28_ <= r_n_366__28_;
      r_366__27_ <= r_n_366__27_;
      r_366__26_ <= r_n_366__26_;
      r_366__25_ <= r_n_366__25_;
      r_366__24_ <= r_n_366__24_;
      r_366__23_ <= r_n_366__23_;
      r_366__22_ <= r_n_366__22_;
      r_366__21_ <= r_n_366__21_;
      r_366__20_ <= r_n_366__20_;
      r_366__19_ <= r_n_366__19_;
      r_366__18_ <= r_n_366__18_;
      r_366__17_ <= r_n_366__17_;
      r_366__16_ <= r_n_366__16_;
      r_366__15_ <= r_n_366__15_;
      r_366__14_ <= r_n_366__14_;
      r_366__13_ <= r_n_366__13_;
      r_366__12_ <= r_n_366__12_;
      r_366__11_ <= r_n_366__11_;
      r_366__10_ <= r_n_366__10_;
      r_366__9_ <= r_n_366__9_;
      r_366__8_ <= r_n_366__8_;
      r_366__7_ <= r_n_366__7_;
      r_366__6_ <= r_n_366__6_;
      r_366__5_ <= r_n_366__5_;
      r_366__4_ <= r_n_366__4_;
      r_366__3_ <= r_n_366__3_;
      r_366__2_ <= r_n_366__2_;
      r_366__1_ <= r_n_366__1_;
      r_366__0_ <= r_n_366__0_;
    end 
    if(N3951) begin
      r_367__63_ <= r_n_367__63_;
      r_367__62_ <= r_n_367__62_;
      r_367__61_ <= r_n_367__61_;
      r_367__60_ <= r_n_367__60_;
      r_367__59_ <= r_n_367__59_;
      r_367__58_ <= r_n_367__58_;
      r_367__57_ <= r_n_367__57_;
      r_367__56_ <= r_n_367__56_;
      r_367__55_ <= r_n_367__55_;
      r_367__54_ <= r_n_367__54_;
      r_367__53_ <= r_n_367__53_;
      r_367__52_ <= r_n_367__52_;
      r_367__51_ <= r_n_367__51_;
      r_367__50_ <= r_n_367__50_;
      r_367__49_ <= r_n_367__49_;
      r_367__48_ <= r_n_367__48_;
      r_367__47_ <= r_n_367__47_;
      r_367__46_ <= r_n_367__46_;
      r_367__45_ <= r_n_367__45_;
      r_367__44_ <= r_n_367__44_;
      r_367__43_ <= r_n_367__43_;
      r_367__42_ <= r_n_367__42_;
      r_367__41_ <= r_n_367__41_;
      r_367__40_ <= r_n_367__40_;
      r_367__39_ <= r_n_367__39_;
      r_367__38_ <= r_n_367__38_;
      r_367__37_ <= r_n_367__37_;
      r_367__36_ <= r_n_367__36_;
      r_367__35_ <= r_n_367__35_;
      r_367__34_ <= r_n_367__34_;
      r_367__33_ <= r_n_367__33_;
      r_367__32_ <= r_n_367__32_;
      r_367__31_ <= r_n_367__31_;
      r_367__30_ <= r_n_367__30_;
      r_367__29_ <= r_n_367__29_;
      r_367__28_ <= r_n_367__28_;
      r_367__27_ <= r_n_367__27_;
      r_367__26_ <= r_n_367__26_;
      r_367__25_ <= r_n_367__25_;
      r_367__24_ <= r_n_367__24_;
      r_367__23_ <= r_n_367__23_;
      r_367__22_ <= r_n_367__22_;
      r_367__21_ <= r_n_367__21_;
      r_367__20_ <= r_n_367__20_;
      r_367__19_ <= r_n_367__19_;
      r_367__18_ <= r_n_367__18_;
      r_367__17_ <= r_n_367__17_;
      r_367__16_ <= r_n_367__16_;
      r_367__15_ <= r_n_367__15_;
      r_367__14_ <= r_n_367__14_;
      r_367__13_ <= r_n_367__13_;
      r_367__12_ <= r_n_367__12_;
      r_367__11_ <= r_n_367__11_;
      r_367__10_ <= r_n_367__10_;
      r_367__9_ <= r_n_367__9_;
      r_367__8_ <= r_n_367__8_;
      r_367__7_ <= r_n_367__7_;
      r_367__6_ <= r_n_367__6_;
      r_367__5_ <= r_n_367__5_;
      r_367__4_ <= r_n_367__4_;
      r_367__3_ <= r_n_367__3_;
      r_367__2_ <= r_n_367__2_;
      r_367__1_ <= r_n_367__1_;
      r_367__0_ <= r_n_367__0_;
    end 
    if(N3952) begin
      r_368__63_ <= r_n_368__63_;
      r_368__62_ <= r_n_368__62_;
      r_368__61_ <= r_n_368__61_;
      r_368__60_ <= r_n_368__60_;
      r_368__59_ <= r_n_368__59_;
      r_368__58_ <= r_n_368__58_;
      r_368__57_ <= r_n_368__57_;
      r_368__56_ <= r_n_368__56_;
      r_368__55_ <= r_n_368__55_;
      r_368__54_ <= r_n_368__54_;
      r_368__53_ <= r_n_368__53_;
      r_368__52_ <= r_n_368__52_;
      r_368__51_ <= r_n_368__51_;
      r_368__50_ <= r_n_368__50_;
      r_368__49_ <= r_n_368__49_;
      r_368__48_ <= r_n_368__48_;
      r_368__47_ <= r_n_368__47_;
      r_368__46_ <= r_n_368__46_;
      r_368__45_ <= r_n_368__45_;
      r_368__44_ <= r_n_368__44_;
      r_368__43_ <= r_n_368__43_;
      r_368__42_ <= r_n_368__42_;
      r_368__41_ <= r_n_368__41_;
      r_368__40_ <= r_n_368__40_;
      r_368__39_ <= r_n_368__39_;
      r_368__38_ <= r_n_368__38_;
      r_368__37_ <= r_n_368__37_;
      r_368__36_ <= r_n_368__36_;
      r_368__35_ <= r_n_368__35_;
      r_368__34_ <= r_n_368__34_;
      r_368__33_ <= r_n_368__33_;
      r_368__32_ <= r_n_368__32_;
      r_368__31_ <= r_n_368__31_;
      r_368__30_ <= r_n_368__30_;
      r_368__29_ <= r_n_368__29_;
      r_368__28_ <= r_n_368__28_;
      r_368__27_ <= r_n_368__27_;
      r_368__26_ <= r_n_368__26_;
      r_368__25_ <= r_n_368__25_;
      r_368__24_ <= r_n_368__24_;
      r_368__23_ <= r_n_368__23_;
      r_368__22_ <= r_n_368__22_;
      r_368__21_ <= r_n_368__21_;
      r_368__20_ <= r_n_368__20_;
      r_368__19_ <= r_n_368__19_;
      r_368__18_ <= r_n_368__18_;
      r_368__17_ <= r_n_368__17_;
      r_368__16_ <= r_n_368__16_;
      r_368__15_ <= r_n_368__15_;
      r_368__14_ <= r_n_368__14_;
      r_368__13_ <= r_n_368__13_;
      r_368__12_ <= r_n_368__12_;
      r_368__11_ <= r_n_368__11_;
      r_368__10_ <= r_n_368__10_;
      r_368__9_ <= r_n_368__9_;
      r_368__8_ <= r_n_368__8_;
      r_368__7_ <= r_n_368__7_;
      r_368__6_ <= r_n_368__6_;
      r_368__5_ <= r_n_368__5_;
      r_368__4_ <= r_n_368__4_;
      r_368__3_ <= r_n_368__3_;
      r_368__2_ <= r_n_368__2_;
      r_368__1_ <= r_n_368__1_;
      r_368__0_ <= r_n_368__0_;
    end 
    if(N3953) begin
      r_369__63_ <= r_n_369__63_;
      r_369__62_ <= r_n_369__62_;
      r_369__61_ <= r_n_369__61_;
      r_369__60_ <= r_n_369__60_;
      r_369__59_ <= r_n_369__59_;
      r_369__58_ <= r_n_369__58_;
      r_369__57_ <= r_n_369__57_;
      r_369__56_ <= r_n_369__56_;
      r_369__55_ <= r_n_369__55_;
      r_369__54_ <= r_n_369__54_;
      r_369__53_ <= r_n_369__53_;
      r_369__52_ <= r_n_369__52_;
      r_369__51_ <= r_n_369__51_;
      r_369__50_ <= r_n_369__50_;
      r_369__49_ <= r_n_369__49_;
      r_369__48_ <= r_n_369__48_;
      r_369__47_ <= r_n_369__47_;
      r_369__46_ <= r_n_369__46_;
      r_369__45_ <= r_n_369__45_;
      r_369__44_ <= r_n_369__44_;
      r_369__43_ <= r_n_369__43_;
      r_369__42_ <= r_n_369__42_;
      r_369__41_ <= r_n_369__41_;
      r_369__40_ <= r_n_369__40_;
      r_369__39_ <= r_n_369__39_;
      r_369__38_ <= r_n_369__38_;
      r_369__37_ <= r_n_369__37_;
      r_369__36_ <= r_n_369__36_;
      r_369__35_ <= r_n_369__35_;
      r_369__34_ <= r_n_369__34_;
      r_369__33_ <= r_n_369__33_;
      r_369__32_ <= r_n_369__32_;
      r_369__31_ <= r_n_369__31_;
      r_369__30_ <= r_n_369__30_;
      r_369__29_ <= r_n_369__29_;
      r_369__28_ <= r_n_369__28_;
      r_369__27_ <= r_n_369__27_;
      r_369__26_ <= r_n_369__26_;
      r_369__25_ <= r_n_369__25_;
      r_369__24_ <= r_n_369__24_;
      r_369__23_ <= r_n_369__23_;
      r_369__22_ <= r_n_369__22_;
      r_369__21_ <= r_n_369__21_;
      r_369__20_ <= r_n_369__20_;
      r_369__19_ <= r_n_369__19_;
      r_369__18_ <= r_n_369__18_;
      r_369__17_ <= r_n_369__17_;
      r_369__16_ <= r_n_369__16_;
      r_369__15_ <= r_n_369__15_;
      r_369__14_ <= r_n_369__14_;
      r_369__13_ <= r_n_369__13_;
      r_369__12_ <= r_n_369__12_;
      r_369__11_ <= r_n_369__11_;
      r_369__10_ <= r_n_369__10_;
      r_369__9_ <= r_n_369__9_;
      r_369__8_ <= r_n_369__8_;
      r_369__7_ <= r_n_369__7_;
      r_369__6_ <= r_n_369__6_;
      r_369__5_ <= r_n_369__5_;
      r_369__4_ <= r_n_369__4_;
      r_369__3_ <= r_n_369__3_;
      r_369__2_ <= r_n_369__2_;
      r_369__1_ <= r_n_369__1_;
      r_369__0_ <= r_n_369__0_;
    end 
    if(N3954) begin
      r_370__63_ <= r_n_370__63_;
      r_370__62_ <= r_n_370__62_;
      r_370__61_ <= r_n_370__61_;
      r_370__60_ <= r_n_370__60_;
      r_370__59_ <= r_n_370__59_;
      r_370__58_ <= r_n_370__58_;
      r_370__57_ <= r_n_370__57_;
      r_370__56_ <= r_n_370__56_;
      r_370__55_ <= r_n_370__55_;
      r_370__54_ <= r_n_370__54_;
      r_370__53_ <= r_n_370__53_;
      r_370__52_ <= r_n_370__52_;
      r_370__51_ <= r_n_370__51_;
      r_370__50_ <= r_n_370__50_;
      r_370__49_ <= r_n_370__49_;
      r_370__48_ <= r_n_370__48_;
      r_370__47_ <= r_n_370__47_;
      r_370__46_ <= r_n_370__46_;
      r_370__45_ <= r_n_370__45_;
      r_370__44_ <= r_n_370__44_;
      r_370__43_ <= r_n_370__43_;
      r_370__42_ <= r_n_370__42_;
      r_370__41_ <= r_n_370__41_;
      r_370__40_ <= r_n_370__40_;
      r_370__39_ <= r_n_370__39_;
      r_370__38_ <= r_n_370__38_;
      r_370__37_ <= r_n_370__37_;
      r_370__36_ <= r_n_370__36_;
      r_370__35_ <= r_n_370__35_;
      r_370__34_ <= r_n_370__34_;
      r_370__33_ <= r_n_370__33_;
      r_370__32_ <= r_n_370__32_;
      r_370__31_ <= r_n_370__31_;
      r_370__30_ <= r_n_370__30_;
      r_370__29_ <= r_n_370__29_;
      r_370__28_ <= r_n_370__28_;
      r_370__27_ <= r_n_370__27_;
      r_370__26_ <= r_n_370__26_;
      r_370__25_ <= r_n_370__25_;
      r_370__24_ <= r_n_370__24_;
      r_370__23_ <= r_n_370__23_;
      r_370__22_ <= r_n_370__22_;
      r_370__21_ <= r_n_370__21_;
      r_370__20_ <= r_n_370__20_;
      r_370__19_ <= r_n_370__19_;
      r_370__18_ <= r_n_370__18_;
      r_370__17_ <= r_n_370__17_;
      r_370__16_ <= r_n_370__16_;
      r_370__15_ <= r_n_370__15_;
      r_370__14_ <= r_n_370__14_;
      r_370__13_ <= r_n_370__13_;
      r_370__12_ <= r_n_370__12_;
      r_370__11_ <= r_n_370__11_;
      r_370__10_ <= r_n_370__10_;
      r_370__9_ <= r_n_370__9_;
      r_370__8_ <= r_n_370__8_;
      r_370__7_ <= r_n_370__7_;
      r_370__6_ <= r_n_370__6_;
      r_370__5_ <= r_n_370__5_;
      r_370__4_ <= r_n_370__4_;
      r_370__3_ <= r_n_370__3_;
      r_370__2_ <= r_n_370__2_;
      r_370__1_ <= r_n_370__1_;
      r_370__0_ <= r_n_370__0_;
    end 
    if(N3955) begin
      r_371__63_ <= r_n_371__63_;
      r_371__62_ <= r_n_371__62_;
      r_371__61_ <= r_n_371__61_;
      r_371__60_ <= r_n_371__60_;
      r_371__59_ <= r_n_371__59_;
      r_371__58_ <= r_n_371__58_;
      r_371__57_ <= r_n_371__57_;
      r_371__56_ <= r_n_371__56_;
      r_371__55_ <= r_n_371__55_;
      r_371__54_ <= r_n_371__54_;
      r_371__53_ <= r_n_371__53_;
      r_371__52_ <= r_n_371__52_;
      r_371__51_ <= r_n_371__51_;
      r_371__50_ <= r_n_371__50_;
      r_371__49_ <= r_n_371__49_;
      r_371__48_ <= r_n_371__48_;
      r_371__47_ <= r_n_371__47_;
      r_371__46_ <= r_n_371__46_;
      r_371__45_ <= r_n_371__45_;
      r_371__44_ <= r_n_371__44_;
      r_371__43_ <= r_n_371__43_;
      r_371__42_ <= r_n_371__42_;
      r_371__41_ <= r_n_371__41_;
      r_371__40_ <= r_n_371__40_;
      r_371__39_ <= r_n_371__39_;
      r_371__38_ <= r_n_371__38_;
      r_371__37_ <= r_n_371__37_;
      r_371__36_ <= r_n_371__36_;
      r_371__35_ <= r_n_371__35_;
      r_371__34_ <= r_n_371__34_;
      r_371__33_ <= r_n_371__33_;
      r_371__32_ <= r_n_371__32_;
      r_371__31_ <= r_n_371__31_;
      r_371__30_ <= r_n_371__30_;
      r_371__29_ <= r_n_371__29_;
      r_371__28_ <= r_n_371__28_;
      r_371__27_ <= r_n_371__27_;
      r_371__26_ <= r_n_371__26_;
      r_371__25_ <= r_n_371__25_;
      r_371__24_ <= r_n_371__24_;
      r_371__23_ <= r_n_371__23_;
      r_371__22_ <= r_n_371__22_;
      r_371__21_ <= r_n_371__21_;
      r_371__20_ <= r_n_371__20_;
      r_371__19_ <= r_n_371__19_;
      r_371__18_ <= r_n_371__18_;
      r_371__17_ <= r_n_371__17_;
      r_371__16_ <= r_n_371__16_;
      r_371__15_ <= r_n_371__15_;
      r_371__14_ <= r_n_371__14_;
      r_371__13_ <= r_n_371__13_;
      r_371__12_ <= r_n_371__12_;
      r_371__11_ <= r_n_371__11_;
      r_371__10_ <= r_n_371__10_;
      r_371__9_ <= r_n_371__9_;
      r_371__8_ <= r_n_371__8_;
      r_371__7_ <= r_n_371__7_;
      r_371__6_ <= r_n_371__6_;
      r_371__5_ <= r_n_371__5_;
      r_371__4_ <= r_n_371__4_;
      r_371__3_ <= r_n_371__3_;
      r_371__2_ <= r_n_371__2_;
      r_371__1_ <= r_n_371__1_;
      r_371__0_ <= r_n_371__0_;
    end 
    if(N3956) begin
      r_372__63_ <= r_n_372__63_;
      r_372__62_ <= r_n_372__62_;
      r_372__61_ <= r_n_372__61_;
      r_372__60_ <= r_n_372__60_;
      r_372__59_ <= r_n_372__59_;
      r_372__58_ <= r_n_372__58_;
      r_372__57_ <= r_n_372__57_;
      r_372__56_ <= r_n_372__56_;
      r_372__55_ <= r_n_372__55_;
      r_372__54_ <= r_n_372__54_;
      r_372__53_ <= r_n_372__53_;
      r_372__52_ <= r_n_372__52_;
      r_372__51_ <= r_n_372__51_;
      r_372__50_ <= r_n_372__50_;
      r_372__49_ <= r_n_372__49_;
      r_372__48_ <= r_n_372__48_;
      r_372__47_ <= r_n_372__47_;
      r_372__46_ <= r_n_372__46_;
      r_372__45_ <= r_n_372__45_;
      r_372__44_ <= r_n_372__44_;
      r_372__43_ <= r_n_372__43_;
      r_372__42_ <= r_n_372__42_;
      r_372__41_ <= r_n_372__41_;
      r_372__40_ <= r_n_372__40_;
      r_372__39_ <= r_n_372__39_;
      r_372__38_ <= r_n_372__38_;
      r_372__37_ <= r_n_372__37_;
      r_372__36_ <= r_n_372__36_;
      r_372__35_ <= r_n_372__35_;
      r_372__34_ <= r_n_372__34_;
      r_372__33_ <= r_n_372__33_;
      r_372__32_ <= r_n_372__32_;
      r_372__31_ <= r_n_372__31_;
      r_372__30_ <= r_n_372__30_;
      r_372__29_ <= r_n_372__29_;
      r_372__28_ <= r_n_372__28_;
      r_372__27_ <= r_n_372__27_;
      r_372__26_ <= r_n_372__26_;
      r_372__25_ <= r_n_372__25_;
      r_372__24_ <= r_n_372__24_;
      r_372__23_ <= r_n_372__23_;
      r_372__22_ <= r_n_372__22_;
      r_372__21_ <= r_n_372__21_;
      r_372__20_ <= r_n_372__20_;
      r_372__19_ <= r_n_372__19_;
      r_372__18_ <= r_n_372__18_;
      r_372__17_ <= r_n_372__17_;
      r_372__16_ <= r_n_372__16_;
      r_372__15_ <= r_n_372__15_;
      r_372__14_ <= r_n_372__14_;
      r_372__13_ <= r_n_372__13_;
      r_372__12_ <= r_n_372__12_;
      r_372__11_ <= r_n_372__11_;
      r_372__10_ <= r_n_372__10_;
      r_372__9_ <= r_n_372__9_;
      r_372__8_ <= r_n_372__8_;
      r_372__7_ <= r_n_372__7_;
      r_372__6_ <= r_n_372__6_;
      r_372__5_ <= r_n_372__5_;
      r_372__4_ <= r_n_372__4_;
      r_372__3_ <= r_n_372__3_;
      r_372__2_ <= r_n_372__2_;
      r_372__1_ <= r_n_372__1_;
      r_372__0_ <= r_n_372__0_;
    end 
    if(N3957) begin
      r_373__63_ <= r_n_373__63_;
      r_373__62_ <= r_n_373__62_;
      r_373__61_ <= r_n_373__61_;
      r_373__60_ <= r_n_373__60_;
      r_373__59_ <= r_n_373__59_;
      r_373__58_ <= r_n_373__58_;
      r_373__57_ <= r_n_373__57_;
      r_373__56_ <= r_n_373__56_;
      r_373__55_ <= r_n_373__55_;
      r_373__54_ <= r_n_373__54_;
      r_373__53_ <= r_n_373__53_;
      r_373__52_ <= r_n_373__52_;
      r_373__51_ <= r_n_373__51_;
      r_373__50_ <= r_n_373__50_;
      r_373__49_ <= r_n_373__49_;
      r_373__48_ <= r_n_373__48_;
      r_373__47_ <= r_n_373__47_;
      r_373__46_ <= r_n_373__46_;
      r_373__45_ <= r_n_373__45_;
      r_373__44_ <= r_n_373__44_;
      r_373__43_ <= r_n_373__43_;
      r_373__42_ <= r_n_373__42_;
      r_373__41_ <= r_n_373__41_;
      r_373__40_ <= r_n_373__40_;
      r_373__39_ <= r_n_373__39_;
      r_373__38_ <= r_n_373__38_;
      r_373__37_ <= r_n_373__37_;
      r_373__36_ <= r_n_373__36_;
      r_373__35_ <= r_n_373__35_;
      r_373__34_ <= r_n_373__34_;
      r_373__33_ <= r_n_373__33_;
      r_373__32_ <= r_n_373__32_;
      r_373__31_ <= r_n_373__31_;
      r_373__30_ <= r_n_373__30_;
      r_373__29_ <= r_n_373__29_;
      r_373__28_ <= r_n_373__28_;
      r_373__27_ <= r_n_373__27_;
      r_373__26_ <= r_n_373__26_;
      r_373__25_ <= r_n_373__25_;
      r_373__24_ <= r_n_373__24_;
      r_373__23_ <= r_n_373__23_;
      r_373__22_ <= r_n_373__22_;
      r_373__21_ <= r_n_373__21_;
      r_373__20_ <= r_n_373__20_;
      r_373__19_ <= r_n_373__19_;
      r_373__18_ <= r_n_373__18_;
      r_373__17_ <= r_n_373__17_;
      r_373__16_ <= r_n_373__16_;
      r_373__15_ <= r_n_373__15_;
      r_373__14_ <= r_n_373__14_;
      r_373__13_ <= r_n_373__13_;
      r_373__12_ <= r_n_373__12_;
      r_373__11_ <= r_n_373__11_;
      r_373__10_ <= r_n_373__10_;
      r_373__9_ <= r_n_373__9_;
      r_373__8_ <= r_n_373__8_;
      r_373__7_ <= r_n_373__7_;
      r_373__6_ <= r_n_373__6_;
      r_373__5_ <= r_n_373__5_;
      r_373__4_ <= r_n_373__4_;
      r_373__3_ <= r_n_373__3_;
      r_373__2_ <= r_n_373__2_;
      r_373__1_ <= r_n_373__1_;
      r_373__0_ <= r_n_373__0_;
    end 
    if(N3958) begin
      r_374__63_ <= r_n_374__63_;
      r_374__62_ <= r_n_374__62_;
      r_374__61_ <= r_n_374__61_;
      r_374__60_ <= r_n_374__60_;
      r_374__59_ <= r_n_374__59_;
      r_374__58_ <= r_n_374__58_;
      r_374__57_ <= r_n_374__57_;
      r_374__56_ <= r_n_374__56_;
      r_374__55_ <= r_n_374__55_;
      r_374__54_ <= r_n_374__54_;
      r_374__53_ <= r_n_374__53_;
      r_374__52_ <= r_n_374__52_;
      r_374__51_ <= r_n_374__51_;
      r_374__50_ <= r_n_374__50_;
      r_374__49_ <= r_n_374__49_;
      r_374__48_ <= r_n_374__48_;
      r_374__47_ <= r_n_374__47_;
      r_374__46_ <= r_n_374__46_;
      r_374__45_ <= r_n_374__45_;
      r_374__44_ <= r_n_374__44_;
      r_374__43_ <= r_n_374__43_;
      r_374__42_ <= r_n_374__42_;
      r_374__41_ <= r_n_374__41_;
      r_374__40_ <= r_n_374__40_;
      r_374__39_ <= r_n_374__39_;
      r_374__38_ <= r_n_374__38_;
      r_374__37_ <= r_n_374__37_;
      r_374__36_ <= r_n_374__36_;
      r_374__35_ <= r_n_374__35_;
      r_374__34_ <= r_n_374__34_;
      r_374__33_ <= r_n_374__33_;
      r_374__32_ <= r_n_374__32_;
      r_374__31_ <= r_n_374__31_;
      r_374__30_ <= r_n_374__30_;
      r_374__29_ <= r_n_374__29_;
      r_374__28_ <= r_n_374__28_;
      r_374__27_ <= r_n_374__27_;
      r_374__26_ <= r_n_374__26_;
      r_374__25_ <= r_n_374__25_;
      r_374__24_ <= r_n_374__24_;
      r_374__23_ <= r_n_374__23_;
      r_374__22_ <= r_n_374__22_;
      r_374__21_ <= r_n_374__21_;
      r_374__20_ <= r_n_374__20_;
      r_374__19_ <= r_n_374__19_;
      r_374__18_ <= r_n_374__18_;
      r_374__17_ <= r_n_374__17_;
      r_374__16_ <= r_n_374__16_;
      r_374__15_ <= r_n_374__15_;
      r_374__14_ <= r_n_374__14_;
      r_374__13_ <= r_n_374__13_;
      r_374__12_ <= r_n_374__12_;
      r_374__11_ <= r_n_374__11_;
      r_374__10_ <= r_n_374__10_;
      r_374__9_ <= r_n_374__9_;
      r_374__8_ <= r_n_374__8_;
      r_374__7_ <= r_n_374__7_;
      r_374__6_ <= r_n_374__6_;
      r_374__5_ <= r_n_374__5_;
      r_374__4_ <= r_n_374__4_;
      r_374__3_ <= r_n_374__3_;
      r_374__2_ <= r_n_374__2_;
      r_374__1_ <= r_n_374__1_;
      r_374__0_ <= r_n_374__0_;
    end 
    if(N3959) begin
      r_375__63_ <= r_n_375__63_;
      r_375__62_ <= r_n_375__62_;
      r_375__61_ <= r_n_375__61_;
      r_375__60_ <= r_n_375__60_;
      r_375__59_ <= r_n_375__59_;
      r_375__58_ <= r_n_375__58_;
      r_375__57_ <= r_n_375__57_;
      r_375__56_ <= r_n_375__56_;
      r_375__55_ <= r_n_375__55_;
      r_375__54_ <= r_n_375__54_;
      r_375__53_ <= r_n_375__53_;
      r_375__52_ <= r_n_375__52_;
      r_375__51_ <= r_n_375__51_;
      r_375__50_ <= r_n_375__50_;
      r_375__49_ <= r_n_375__49_;
      r_375__48_ <= r_n_375__48_;
      r_375__47_ <= r_n_375__47_;
      r_375__46_ <= r_n_375__46_;
      r_375__45_ <= r_n_375__45_;
      r_375__44_ <= r_n_375__44_;
      r_375__43_ <= r_n_375__43_;
      r_375__42_ <= r_n_375__42_;
      r_375__41_ <= r_n_375__41_;
      r_375__40_ <= r_n_375__40_;
      r_375__39_ <= r_n_375__39_;
      r_375__38_ <= r_n_375__38_;
      r_375__37_ <= r_n_375__37_;
      r_375__36_ <= r_n_375__36_;
      r_375__35_ <= r_n_375__35_;
      r_375__34_ <= r_n_375__34_;
      r_375__33_ <= r_n_375__33_;
      r_375__32_ <= r_n_375__32_;
      r_375__31_ <= r_n_375__31_;
      r_375__30_ <= r_n_375__30_;
      r_375__29_ <= r_n_375__29_;
      r_375__28_ <= r_n_375__28_;
      r_375__27_ <= r_n_375__27_;
      r_375__26_ <= r_n_375__26_;
      r_375__25_ <= r_n_375__25_;
      r_375__24_ <= r_n_375__24_;
      r_375__23_ <= r_n_375__23_;
      r_375__22_ <= r_n_375__22_;
      r_375__21_ <= r_n_375__21_;
      r_375__20_ <= r_n_375__20_;
      r_375__19_ <= r_n_375__19_;
      r_375__18_ <= r_n_375__18_;
      r_375__17_ <= r_n_375__17_;
      r_375__16_ <= r_n_375__16_;
      r_375__15_ <= r_n_375__15_;
      r_375__14_ <= r_n_375__14_;
      r_375__13_ <= r_n_375__13_;
      r_375__12_ <= r_n_375__12_;
      r_375__11_ <= r_n_375__11_;
      r_375__10_ <= r_n_375__10_;
      r_375__9_ <= r_n_375__9_;
      r_375__8_ <= r_n_375__8_;
      r_375__7_ <= r_n_375__7_;
      r_375__6_ <= r_n_375__6_;
      r_375__5_ <= r_n_375__5_;
      r_375__4_ <= r_n_375__4_;
      r_375__3_ <= r_n_375__3_;
      r_375__2_ <= r_n_375__2_;
      r_375__1_ <= r_n_375__1_;
      r_375__0_ <= r_n_375__0_;
    end 
    if(N3960) begin
      r_376__63_ <= r_n_376__63_;
      r_376__62_ <= r_n_376__62_;
      r_376__61_ <= r_n_376__61_;
      r_376__60_ <= r_n_376__60_;
      r_376__59_ <= r_n_376__59_;
      r_376__58_ <= r_n_376__58_;
      r_376__57_ <= r_n_376__57_;
      r_376__56_ <= r_n_376__56_;
      r_376__55_ <= r_n_376__55_;
      r_376__54_ <= r_n_376__54_;
      r_376__53_ <= r_n_376__53_;
      r_376__52_ <= r_n_376__52_;
      r_376__51_ <= r_n_376__51_;
      r_376__50_ <= r_n_376__50_;
      r_376__49_ <= r_n_376__49_;
      r_376__48_ <= r_n_376__48_;
      r_376__47_ <= r_n_376__47_;
      r_376__46_ <= r_n_376__46_;
      r_376__45_ <= r_n_376__45_;
      r_376__44_ <= r_n_376__44_;
      r_376__43_ <= r_n_376__43_;
      r_376__42_ <= r_n_376__42_;
      r_376__41_ <= r_n_376__41_;
      r_376__40_ <= r_n_376__40_;
      r_376__39_ <= r_n_376__39_;
      r_376__38_ <= r_n_376__38_;
      r_376__37_ <= r_n_376__37_;
      r_376__36_ <= r_n_376__36_;
      r_376__35_ <= r_n_376__35_;
      r_376__34_ <= r_n_376__34_;
      r_376__33_ <= r_n_376__33_;
      r_376__32_ <= r_n_376__32_;
      r_376__31_ <= r_n_376__31_;
      r_376__30_ <= r_n_376__30_;
      r_376__29_ <= r_n_376__29_;
      r_376__28_ <= r_n_376__28_;
      r_376__27_ <= r_n_376__27_;
      r_376__26_ <= r_n_376__26_;
      r_376__25_ <= r_n_376__25_;
      r_376__24_ <= r_n_376__24_;
      r_376__23_ <= r_n_376__23_;
      r_376__22_ <= r_n_376__22_;
      r_376__21_ <= r_n_376__21_;
      r_376__20_ <= r_n_376__20_;
      r_376__19_ <= r_n_376__19_;
      r_376__18_ <= r_n_376__18_;
      r_376__17_ <= r_n_376__17_;
      r_376__16_ <= r_n_376__16_;
      r_376__15_ <= r_n_376__15_;
      r_376__14_ <= r_n_376__14_;
      r_376__13_ <= r_n_376__13_;
      r_376__12_ <= r_n_376__12_;
      r_376__11_ <= r_n_376__11_;
      r_376__10_ <= r_n_376__10_;
      r_376__9_ <= r_n_376__9_;
      r_376__8_ <= r_n_376__8_;
      r_376__7_ <= r_n_376__7_;
      r_376__6_ <= r_n_376__6_;
      r_376__5_ <= r_n_376__5_;
      r_376__4_ <= r_n_376__4_;
      r_376__3_ <= r_n_376__3_;
      r_376__2_ <= r_n_376__2_;
      r_376__1_ <= r_n_376__1_;
      r_376__0_ <= r_n_376__0_;
    end 
    if(N3961) begin
      r_377__63_ <= r_n_377__63_;
      r_377__62_ <= r_n_377__62_;
      r_377__61_ <= r_n_377__61_;
      r_377__60_ <= r_n_377__60_;
      r_377__59_ <= r_n_377__59_;
      r_377__58_ <= r_n_377__58_;
      r_377__57_ <= r_n_377__57_;
      r_377__56_ <= r_n_377__56_;
      r_377__55_ <= r_n_377__55_;
      r_377__54_ <= r_n_377__54_;
      r_377__53_ <= r_n_377__53_;
      r_377__52_ <= r_n_377__52_;
      r_377__51_ <= r_n_377__51_;
      r_377__50_ <= r_n_377__50_;
      r_377__49_ <= r_n_377__49_;
      r_377__48_ <= r_n_377__48_;
      r_377__47_ <= r_n_377__47_;
      r_377__46_ <= r_n_377__46_;
      r_377__45_ <= r_n_377__45_;
      r_377__44_ <= r_n_377__44_;
      r_377__43_ <= r_n_377__43_;
      r_377__42_ <= r_n_377__42_;
      r_377__41_ <= r_n_377__41_;
      r_377__40_ <= r_n_377__40_;
      r_377__39_ <= r_n_377__39_;
      r_377__38_ <= r_n_377__38_;
      r_377__37_ <= r_n_377__37_;
      r_377__36_ <= r_n_377__36_;
      r_377__35_ <= r_n_377__35_;
      r_377__34_ <= r_n_377__34_;
      r_377__33_ <= r_n_377__33_;
      r_377__32_ <= r_n_377__32_;
      r_377__31_ <= r_n_377__31_;
      r_377__30_ <= r_n_377__30_;
      r_377__29_ <= r_n_377__29_;
      r_377__28_ <= r_n_377__28_;
      r_377__27_ <= r_n_377__27_;
      r_377__26_ <= r_n_377__26_;
      r_377__25_ <= r_n_377__25_;
      r_377__24_ <= r_n_377__24_;
      r_377__23_ <= r_n_377__23_;
      r_377__22_ <= r_n_377__22_;
      r_377__21_ <= r_n_377__21_;
      r_377__20_ <= r_n_377__20_;
      r_377__19_ <= r_n_377__19_;
      r_377__18_ <= r_n_377__18_;
      r_377__17_ <= r_n_377__17_;
      r_377__16_ <= r_n_377__16_;
      r_377__15_ <= r_n_377__15_;
      r_377__14_ <= r_n_377__14_;
      r_377__13_ <= r_n_377__13_;
      r_377__12_ <= r_n_377__12_;
      r_377__11_ <= r_n_377__11_;
      r_377__10_ <= r_n_377__10_;
      r_377__9_ <= r_n_377__9_;
      r_377__8_ <= r_n_377__8_;
      r_377__7_ <= r_n_377__7_;
      r_377__6_ <= r_n_377__6_;
      r_377__5_ <= r_n_377__5_;
      r_377__4_ <= r_n_377__4_;
      r_377__3_ <= r_n_377__3_;
      r_377__2_ <= r_n_377__2_;
      r_377__1_ <= r_n_377__1_;
      r_377__0_ <= r_n_377__0_;
    end 
    if(N3962) begin
      r_378__63_ <= r_n_378__63_;
      r_378__62_ <= r_n_378__62_;
      r_378__61_ <= r_n_378__61_;
      r_378__60_ <= r_n_378__60_;
      r_378__59_ <= r_n_378__59_;
      r_378__58_ <= r_n_378__58_;
      r_378__57_ <= r_n_378__57_;
      r_378__56_ <= r_n_378__56_;
      r_378__55_ <= r_n_378__55_;
      r_378__54_ <= r_n_378__54_;
      r_378__53_ <= r_n_378__53_;
      r_378__52_ <= r_n_378__52_;
      r_378__51_ <= r_n_378__51_;
      r_378__50_ <= r_n_378__50_;
      r_378__49_ <= r_n_378__49_;
      r_378__48_ <= r_n_378__48_;
      r_378__47_ <= r_n_378__47_;
      r_378__46_ <= r_n_378__46_;
      r_378__45_ <= r_n_378__45_;
      r_378__44_ <= r_n_378__44_;
      r_378__43_ <= r_n_378__43_;
      r_378__42_ <= r_n_378__42_;
      r_378__41_ <= r_n_378__41_;
      r_378__40_ <= r_n_378__40_;
      r_378__39_ <= r_n_378__39_;
      r_378__38_ <= r_n_378__38_;
      r_378__37_ <= r_n_378__37_;
      r_378__36_ <= r_n_378__36_;
      r_378__35_ <= r_n_378__35_;
      r_378__34_ <= r_n_378__34_;
      r_378__33_ <= r_n_378__33_;
      r_378__32_ <= r_n_378__32_;
      r_378__31_ <= r_n_378__31_;
      r_378__30_ <= r_n_378__30_;
      r_378__29_ <= r_n_378__29_;
      r_378__28_ <= r_n_378__28_;
      r_378__27_ <= r_n_378__27_;
      r_378__26_ <= r_n_378__26_;
      r_378__25_ <= r_n_378__25_;
      r_378__24_ <= r_n_378__24_;
      r_378__23_ <= r_n_378__23_;
      r_378__22_ <= r_n_378__22_;
      r_378__21_ <= r_n_378__21_;
      r_378__20_ <= r_n_378__20_;
      r_378__19_ <= r_n_378__19_;
      r_378__18_ <= r_n_378__18_;
      r_378__17_ <= r_n_378__17_;
      r_378__16_ <= r_n_378__16_;
      r_378__15_ <= r_n_378__15_;
      r_378__14_ <= r_n_378__14_;
      r_378__13_ <= r_n_378__13_;
      r_378__12_ <= r_n_378__12_;
      r_378__11_ <= r_n_378__11_;
      r_378__10_ <= r_n_378__10_;
      r_378__9_ <= r_n_378__9_;
      r_378__8_ <= r_n_378__8_;
      r_378__7_ <= r_n_378__7_;
      r_378__6_ <= r_n_378__6_;
      r_378__5_ <= r_n_378__5_;
      r_378__4_ <= r_n_378__4_;
      r_378__3_ <= r_n_378__3_;
      r_378__2_ <= r_n_378__2_;
      r_378__1_ <= r_n_378__1_;
      r_378__0_ <= r_n_378__0_;
    end 
    if(N3963) begin
      r_379__63_ <= r_n_379__63_;
      r_379__62_ <= r_n_379__62_;
      r_379__61_ <= r_n_379__61_;
      r_379__60_ <= r_n_379__60_;
      r_379__59_ <= r_n_379__59_;
      r_379__58_ <= r_n_379__58_;
      r_379__57_ <= r_n_379__57_;
      r_379__56_ <= r_n_379__56_;
      r_379__55_ <= r_n_379__55_;
      r_379__54_ <= r_n_379__54_;
      r_379__53_ <= r_n_379__53_;
      r_379__52_ <= r_n_379__52_;
      r_379__51_ <= r_n_379__51_;
      r_379__50_ <= r_n_379__50_;
      r_379__49_ <= r_n_379__49_;
      r_379__48_ <= r_n_379__48_;
      r_379__47_ <= r_n_379__47_;
      r_379__46_ <= r_n_379__46_;
      r_379__45_ <= r_n_379__45_;
      r_379__44_ <= r_n_379__44_;
      r_379__43_ <= r_n_379__43_;
      r_379__42_ <= r_n_379__42_;
      r_379__41_ <= r_n_379__41_;
      r_379__40_ <= r_n_379__40_;
      r_379__39_ <= r_n_379__39_;
      r_379__38_ <= r_n_379__38_;
      r_379__37_ <= r_n_379__37_;
      r_379__36_ <= r_n_379__36_;
      r_379__35_ <= r_n_379__35_;
      r_379__34_ <= r_n_379__34_;
      r_379__33_ <= r_n_379__33_;
      r_379__32_ <= r_n_379__32_;
      r_379__31_ <= r_n_379__31_;
      r_379__30_ <= r_n_379__30_;
      r_379__29_ <= r_n_379__29_;
      r_379__28_ <= r_n_379__28_;
      r_379__27_ <= r_n_379__27_;
      r_379__26_ <= r_n_379__26_;
      r_379__25_ <= r_n_379__25_;
      r_379__24_ <= r_n_379__24_;
      r_379__23_ <= r_n_379__23_;
      r_379__22_ <= r_n_379__22_;
      r_379__21_ <= r_n_379__21_;
      r_379__20_ <= r_n_379__20_;
      r_379__19_ <= r_n_379__19_;
      r_379__18_ <= r_n_379__18_;
      r_379__17_ <= r_n_379__17_;
      r_379__16_ <= r_n_379__16_;
      r_379__15_ <= r_n_379__15_;
      r_379__14_ <= r_n_379__14_;
      r_379__13_ <= r_n_379__13_;
      r_379__12_ <= r_n_379__12_;
      r_379__11_ <= r_n_379__11_;
      r_379__10_ <= r_n_379__10_;
      r_379__9_ <= r_n_379__9_;
      r_379__8_ <= r_n_379__8_;
      r_379__7_ <= r_n_379__7_;
      r_379__6_ <= r_n_379__6_;
      r_379__5_ <= r_n_379__5_;
      r_379__4_ <= r_n_379__4_;
      r_379__3_ <= r_n_379__3_;
      r_379__2_ <= r_n_379__2_;
      r_379__1_ <= r_n_379__1_;
      r_379__0_ <= r_n_379__0_;
    end 
    if(N3964) begin
      r_380__63_ <= r_n_380__63_;
      r_380__62_ <= r_n_380__62_;
      r_380__61_ <= r_n_380__61_;
      r_380__60_ <= r_n_380__60_;
      r_380__59_ <= r_n_380__59_;
      r_380__58_ <= r_n_380__58_;
      r_380__57_ <= r_n_380__57_;
      r_380__56_ <= r_n_380__56_;
      r_380__55_ <= r_n_380__55_;
      r_380__54_ <= r_n_380__54_;
      r_380__53_ <= r_n_380__53_;
      r_380__52_ <= r_n_380__52_;
      r_380__51_ <= r_n_380__51_;
      r_380__50_ <= r_n_380__50_;
      r_380__49_ <= r_n_380__49_;
      r_380__48_ <= r_n_380__48_;
      r_380__47_ <= r_n_380__47_;
      r_380__46_ <= r_n_380__46_;
      r_380__45_ <= r_n_380__45_;
      r_380__44_ <= r_n_380__44_;
      r_380__43_ <= r_n_380__43_;
      r_380__42_ <= r_n_380__42_;
      r_380__41_ <= r_n_380__41_;
      r_380__40_ <= r_n_380__40_;
      r_380__39_ <= r_n_380__39_;
      r_380__38_ <= r_n_380__38_;
      r_380__37_ <= r_n_380__37_;
      r_380__36_ <= r_n_380__36_;
      r_380__35_ <= r_n_380__35_;
      r_380__34_ <= r_n_380__34_;
      r_380__33_ <= r_n_380__33_;
      r_380__32_ <= r_n_380__32_;
      r_380__31_ <= r_n_380__31_;
      r_380__30_ <= r_n_380__30_;
      r_380__29_ <= r_n_380__29_;
      r_380__28_ <= r_n_380__28_;
      r_380__27_ <= r_n_380__27_;
      r_380__26_ <= r_n_380__26_;
      r_380__25_ <= r_n_380__25_;
      r_380__24_ <= r_n_380__24_;
      r_380__23_ <= r_n_380__23_;
      r_380__22_ <= r_n_380__22_;
      r_380__21_ <= r_n_380__21_;
      r_380__20_ <= r_n_380__20_;
      r_380__19_ <= r_n_380__19_;
      r_380__18_ <= r_n_380__18_;
      r_380__17_ <= r_n_380__17_;
      r_380__16_ <= r_n_380__16_;
      r_380__15_ <= r_n_380__15_;
      r_380__14_ <= r_n_380__14_;
      r_380__13_ <= r_n_380__13_;
      r_380__12_ <= r_n_380__12_;
      r_380__11_ <= r_n_380__11_;
      r_380__10_ <= r_n_380__10_;
      r_380__9_ <= r_n_380__9_;
      r_380__8_ <= r_n_380__8_;
      r_380__7_ <= r_n_380__7_;
      r_380__6_ <= r_n_380__6_;
      r_380__5_ <= r_n_380__5_;
      r_380__4_ <= r_n_380__4_;
      r_380__3_ <= r_n_380__3_;
      r_380__2_ <= r_n_380__2_;
      r_380__1_ <= r_n_380__1_;
      r_380__0_ <= r_n_380__0_;
    end 
    if(N3965) begin
      r_381__63_ <= r_n_381__63_;
      r_381__62_ <= r_n_381__62_;
      r_381__61_ <= r_n_381__61_;
      r_381__60_ <= r_n_381__60_;
      r_381__59_ <= r_n_381__59_;
      r_381__58_ <= r_n_381__58_;
      r_381__57_ <= r_n_381__57_;
      r_381__56_ <= r_n_381__56_;
      r_381__55_ <= r_n_381__55_;
      r_381__54_ <= r_n_381__54_;
      r_381__53_ <= r_n_381__53_;
      r_381__52_ <= r_n_381__52_;
      r_381__51_ <= r_n_381__51_;
      r_381__50_ <= r_n_381__50_;
      r_381__49_ <= r_n_381__49_;
      r_381__48_ <= r_n_381__48_;
      r_381__47_ <= r_n_381__47_;
      r_381__46_ <= r_n_381__46_;
      r_381__45_ <= r_n_381__45_;
      r_381__44_ <= r_n_381__44_;
      r_381__43_ <= r_n_381__43_;
      r_381__42_ <= r_n_381__42_;
      r_381__41_ <= r_n_381__41_;
      r_381__40_ <= r_n_381__40_;
      r_381__39_ <= r_n_381__39_;
      r_381__38_ <= r_n_381__38_;
      r_381__37_ <= r_n_381__37_;
      r_381__36_ <= r_n_381__36_;
      r_381__35_ <= r_n_381__35_;
      r_381__34_ <= r_n_381__34_;
      r_381__33_ <= r_n_381__33_;
      r_381__32_ <= r_n_381__32_;
      r_381__31_ <= r_n_381__31_;
      r_381__30_ <= r_n_381__30_;
      r_381__29_ <= r_n_381__29_;
      r_381__28_ <= r_n_381__28_;
      r_381__27_ <= r_n_381__27_;
      r_381__26_ <= r_n_381__26_;
      r_381__25_ <= r_n_381__25_;
      r_381__24_ <= r_n_381__24_;
      r_381__23_ <= r_n_381__23_;
      r_381__22_ <= r_n_381__22_;
      r_381__21_ <= r_n_381__21_;
      r_381__20_ <= r_n_381__20_;
      r_381__19_ <= r_n_381__19_;
      r_381__18_ <= r_n_381__18_;
      r_381__17_ <= r_n_381__17_;
      r_381__16_ <= r_n_381__16_;
      r_381__15_ <= r_n_381__15_;
      r_381__14_ <= r_n_381__14_;
      r_381__13_ <= r_n_381__13_;
      r_381__12_ <= r_n_381__12_;
      r_381__11_ <= r_n_381__11_;
      r_381__10_ <= r_n_381__10_;
      r_381__9_ <= r_n_381__9_;
      r_381__8_ <= r_n_381__8_;
      r_381__7_ <= r_n_381__7_;
      r_381__6_ <= r_n_381__6_;
      r_381__5_ <= r_n_381__5_;
      r_381__4_ <= r_n_381__4_;
      r_381__3_ <= r_n_381__3_;
      r_381__2_ <= r_n_381__2_;
      r_381__1_ <= r_n_381__1_;
      r_381__0_ <= r_n_381__0_;
    end 
    if(N3966) begin
      r_382__63_ <= r_n_382__63_;
      r_382__62_ <= r_n_382__62_;
      r_382__61_ <= r_n_382__61_;
      r_382__60_ <= r_n_382__60_;
      r_382__59_ <= r_n_382__59_;
      r_382__58_ <= r_n_382__58_;
      r_382__57_ <= r_n_382__57_;
      r_382__56_ <= r_n_382__56_;
      r_382__55_ <= r_n_382__55_;
      r_382__54_ <= r_n_382__54_;
      r_382__53_ <= r_n_382__53_;
      r_382__52_ <= r_n_382__52_;
      r_382__51_ <= r_n_382__51_;
      r_382__50_ <= r_n_382__50_;
      r_382__49_ <= r_n_382__49_;
      r_382__48_ <= r_n_382__48_;
      r_382__47_ <= r_n_382__47_;
      r_382__46_ <= r_n_382__46_;
      r_382__45_ <= r_n_382__45_;
      r_382__44_ <= r_n_382__44_;
      r_382__43_ <= r_n_382__43_;
      r_382__42_ <= r_n_382__42_;
      r_382__41_ <= r_n_382__41_;
      r_382__40_ <= r_n_382__40_;
      r_382__39_ <= r_n_382__39_;
      r_382__38_ <= r_n_382__38_;
      r_382__37_ <= r_n_382__37_;
      r_382__36_ <= r_n_382__36_;
      r_382__35_ <= r_n_382__35_;
      r_382__34_ <= r_n_382__34_;
      r_382__33_ <= r_n_382__33_;
      r_382__32_ <= r_n_382__32_;
      r_382__31_ <= r_n_382__31_;
      r_382__30_ <= r_n_382__30_;
      r_382__29_ <= r_n_382__29_;
      r_382__28_ <= r_n_382__28_;
      r_382__27_ <= r_n_382__27_;
      r_382__26_ <= r_n_382__26_;
      r_382__25_ <= r_n_382__25_;
      r_382__24_ <= r_n_382__24_;
      r_382__23_ <= r_n_382__23_;
      r_382__22_ <= r_n_382__22_;
      r_382__21_ <= r_n_382__21_;
      r_382__20_ <= r_n_382__20_;
      r_382__19_ <= r_n_382__19_;
      r_382__18_ <= r_n_382__18_;
      r_382__17_ <= r_n_382__17_;
      r_382__16_ <= r_n_382__16_;
      r_382__15_ <= r_n_382__15_;
      r_382__14_ <= r_n_382__14_;
      r_382__13_ <= r_n_382__13_;
      r_382__12_ <= r_n_382__12_;
      r_382__11_ <= r_n_382__11_;
      r_382__10_ <= r_n_382__10_;
      r_382__9_ <= r_n_382__9_;
      r_382__8_ <= r_n_382__8_;
      r_382__7_ <= r_n_382__7_;
      r_382__6_ <= r_n_382__6_;
      r_382__5_ <= r_n_382__5_;
      r_382__4_ <= r_n_382__4_;
      r_382__3_ <= r_n_382__3_;
      r_382__2_ <= r_n_382__2_;
      r_382__1_ <= r_n_382__1_;
      r_382__0_ <= r_n_382__0_;
    end 
    if(N3967) begin
      r_383__63_ <= r_n_383__63_;
      r_383__62_ <= r_n_383__62_;
      r_383__61_ <= r_n_383__61_;
      r_383__60_ <= r_n_383__60_;
      r_383__59_ <= r_n_383__59_;
      r_383__58_ <= r_n_383__58_;
      r_383__57_ <= r_n_383__57_;
      r_383__56_ <= r_n_383__56_;
      r_383__55_ <= r_n_383__55_;
      r_383__54_ <= r_n_383__54_;
      r_383__53_ <= r_n_383__53_;
      r_383__52_ <= r_n_383__52_;
      r_383__51_ <= r_n_383__51_;
      r_383__50_ <= r_n_383__50_;
      r_383__49_ <= r_n_383__49_;
      r_383__48_ <= r_n_383__48_;
      r_383__47_ <= r_n_383__47_;
      r_383__46_ <= r_n_383__46_;
      r_383__45_ <= r_n_383__45_;
      r_383__44_ <= r_n_383__44_;
      r_383__43_ <= r_n_383__43_;
      r_383__42_ <= r_n_383__42_;
      r_383__41_ <= r_n_383__41_;
      r_383__40_ <= r_n_383__40_;
      r_383__39_ <= r_n_383__39_;
      r_383__38_ <= r_n_383__38_;
      r_383__37_ <= r_n_383__37_;
      r_383__36_ <= r_n_383__36_;
      r_383__35_ <= r_n_383__35_;
      r_383__34_ <= r_n_383__34_;
      r_383__33_ <= r_n_383__33_;
      r_383__32_ <= r_n_383__32_;
      r_383__31_ <= r_n_383__31_;
      r_383__30_ <= r_n_383__30_;
      r_383__29_ <= r_n_383__29_;
      r_383__28_ <= r_n_383__28_;
      r_383__27_ <= r_n_383__27_;
      r_383__26_ <= r_n_383__26_;
      r_383__25_ <= r_n_383__25_;
      r_383__24_ <= r_n_383__24_;
      r_383__23_ <= r_n_383__23_;
      r_383__22_ <= r_n_383__22_;
      r_383__21_ <= r_n_383__21_;
      r_383__20_ <= r_n_383__20_;
      r_383__19_ <= r_n_383__19_;
      r_383__18_ <= r_n_383__18_;
      r_383__17_ <= r_n_383__17_;
      r_383__16_ <= r_n_383__16_;
      r_383__15_ <= r_n_383__15_;
      r_383__14_ <= r_n_383__14_;
      r_383__13_ <= r_n_383__13_;
      r_383__12_ <= r_n_383__12_;
      r_383__11_ <= r_n_383__11_;
      r_383__10_ <= r_n_383__10_;
      r_383__9_ <= r_n_383__9_;
      r_383__8_ <= r_n_383__8_;
      r_383__7_ <= r_n_383__7_;
      r_383__6_ <= r_n_383__6_;
      r_383__5_ <= r_n_383__5_;
      r_383__4_ <= r_n_383__4_;
      r_383__3_ <= r_n_383__3_;
      r_383__2_ <= r_n_383__2_;
      r_383__1_ <= r_n_383__1_;
      r_383__0_ <= r_n_383__0_;
    end 
    if(N3968) begin
      r_384__63_ <= r_n_384__63_;
      r_384__62_ <= r_n_384__62_;
      r_384__61_ <= r_n_384__61_;
      r_384__60_ <= r_n_384__60_;
      r_384__59_ <= r_n_384__59_;
      r_384__58_ <= r_n_384__58_;
      r_384__57_ <= r_n_384__57_;
      r_384__56_ <= r_n_384__56_;
      r_384__55_ <= r_n_384__55_;
      r_384__54_ <= r_n_384__54_;
      r_384__53_ <= r_n_384__53_;
      r_384__52_ <= r_n_384__52_;
      r_384__51_ <= r_n_384__51_;
      r_384__50_ <= r_n_384__50_;
      r_384__49_ <= r_n_384__49_;
      r_384__48_ <= r_n_384__48_;
      r_384__47_ <= r_n_384__47_;
      r_384__46_ <= r_n_384__46_;
      r_384__45_ <= r_n_384__45_;
      r_384__44_ <= r_n_384__44_;
      r_384__43_ <= r_n_384__43_;
      r_384__42_ <= r_n_384__42_;
      r_384__41_ <= r_n_384__41_;
      r_384__40_ <= r_n_384__40_;
      r_384__39_ <= r_n_384__39_;
      r_384__38_ <= r_n_384__38_;
      r_384__37_ <= r_n_384__37_;
      r_384__36_ <= r_n_384__36_;
      r_384__35_ <= r_n_384__35_;
      r_384__34_ <= r_n_384__34_;
      r_384__33_ <= r_n_384__33_;
      r_384__32_ <= r_n_384__32_;
      r_384__31_ <= r_n_384__31_;
      r_384__30_ <= r_n_384__30_;
      r_384__29_ <= r_n_384__29_;
      r_384__28_ <= r_n_384__28_;
      r_384__27_ <= r_n_384__27_;
      r_384__26_ <= r_n_384__26_;
      r_384__25_ <= r_n_384__25_;
      r_384__24_ <= r_n_384__24_;
      r_384__23_ <= r_n_384__23_;
      r_384__22_ <= r_n_384__22_;
      r_384__21_ <= r_n_384__21_;
      r_384__20_ <= r_n_384__20_;
      r_384__19_ <= r_n_384__19_;
      r_384__18_ <= r_n_384__18_;
      r_384__17_ <= r_n_384__17_;
      r_384__16_ <= r_n_384__16_;
      r_384__15_ <= r_n_384__15_;
      r_384__14_ <= r_n_384__14_;
      r_384__13_ <= r_n_384__13_;
      r_384__12_ <= r_n_384__12_;
      r_384__11_ <= r_n_384__11_;
      r_384__10_ <= r_n_384__10_;
      r_384__9_ <= r_n_384__9_;
      r_384__8_ <= r_n_384__8_;
      r_384__7_ <= r_n_384__7_;
      r_384__6_ <= r_n_384__6_;
      r_384__5_ <= r_n_384__5_;
      r_384__4_ <= r_n_384__4_;
      r_384__3_ <= r_n_384__3_;
      r_384__2_ <= r_n_384__2_;
      r_384__1_ <= r_n_384__1_;
      r_384__0_ <= r_n_384__0_;
    end 
    if(N3969) begin
      r_385__63_ <= r_n_385__63_;
      r_385__62_ <= r_n_385__62_;
      r_385__61_ <= r_n_385__61_;
      r_385__60_ <= r_n_385__60_;
      r_385__59_ <= r_n_385__59_;
      r_385__58_ <= r_n_385__58_;
      r_385__57_ <= r_n_385__57_;
      r_385__56_ <= r_n_385__56_;
      r_385__55_ <= r_n_385__55_;
      r_385__54_ <= r_n_385__54_;
      r_385__53_ <= r_n_385__53_;
      r_385__52_ <= r_n_385__52_;
      r_385__51_ <= r_n_385__51_;
      r_385__50_ <= r_n_385__50_;
      r_385__49_ <= r_n_385__49_;
      r_385__48_ <= r_n_385__48_;
      r_385__47_ <= r_n_385__47_;
      r_385__46_ <= r_n_385__46_;
      r_385__45_ <= r_n_385__45_;
      r_385__44_ <= r_n_385__44_;
      r_385__43_ <= r_n_385__43_;
      r_385__42_ <= r_n_385__42_;
      r_385__41_ <= r_n_385__41_;
      r_385__40_ <= r_n_385__40_;
      r_385__39_ <= r_n_385__39_;
      r_385__38_ <= r_n_385__38_;
      r_385__37_ <= r_n_385__37_;
      r_385__36_ <= r_n_385__36_;
      r_385__35_ <= r_n_385__35_;
      r_385__34_ <= r_n_385__34_;
      r_385__33_ <= r_n_385__33_;
      r_385__32_ <= r_n_385__32_;
      r_385__31_ <= r_n_385__31_;
      r_385__30_ <= r_n_385__30_;
      r_385__29_ <= r_n_385__29_;
      r_385__28_ <= r_n_385__28_;
      r_385__27_ <= r_n_385__27_;
      r_385__26_ <= r_n_385__26_;
      r_385__25_ <= r_n_385__25_;
      r_385__24_ <= r_n_385__24_;
      r_385__23_ <= r_n_385__23_;
      r_385__22_ <= r_n_385__22_;
      r_385__21_ <= r_n_385__21_;
      r_385__20_ <= r_n_385__20_;
      r_385__19_ <= r_n_385__19_;
      r_385__18_ <= r_n_385__18_;
      r_385__17_ <= r_n_385__17_;
      r_385__16_ <= r_n_385__16_;
      r_385__15_ <= r_n_385__15_;
      r_385__14_ <= r_n_385__14_;
      r_385__13_ <= r_n_385__13_;
      r_385__12_ <= r_n_385__12_;
      r_385__11_ <= r_n_385__11_;
      r_385__10_ <= r_n_385__10_;
      r_385__9_ <= r_n_385__9_;
      r_385__8_ <= r_n_385__8_;
      r_385__7_ <= r_n_385__7_;
      r_385__6_ <= r_n_385__6_;
      r_385__5_ <= r_n_385__5_;
      r_385__4_ <= r_n_385__4_;
      r_385__3_ <= r_n_385__3_;
      r_385__2_ <= r_n_385__2_;
      r_385__1_ <= r_n_385__1_;
      r_385__0_ <= r_n_385__0_;
    end 
    if(N3970) begin
      r_386__63_ <= r_n_386__63_;
      r_386__62_ <= r_n_386__62_;
      r_386__61_ <= r_n_386__61_;
      r_386__60_ <= r_n_386__60_;
      r_386__59_ <= r_n_386__59_;
      r_386__58_ <= r_n_386__58_;
      r_386__57_ <= r_n_386__57_;
      r_386__56_ <= r_n_386__56_;
      r_386__55_ <= r_n_386__55_;
      r_386__54_ <= r_n_386__54_;
      r_386__53_ <= r_n_386__53_;
      r_386__52_ <= r_n_386__52_;
      r_386__51_ <= r_n_386__51_;
      r_386__50_ <= r_n_386__50_;
      r_386__49_ <= r_n_386__49_;
      r_386__48_ <= r_n_386__48_;
      r_386__47_ <= r_n_386__47_;
      r_386__46_ <= r_n_386__46_;
      r_386__45_ <= r_n_386__45_;
      r_386__44_ <= r_n_386__44_;
      r_386__43_ <= r_n_386__43_;
      r_386__42_ <= r_n_386__42_;
      r_386__41_ <= r_n_386__41_;
      r_386__40_ <= r_n_386__40_;
      r_386__39_ <= r_n_386__39_;
      r_386__38_ <= r_n_386__38_;
      r_386__37_ <= r_n_386__37_;
      r_386__36_ <= r_n_386__36_;
      r_386__35_ <= r_n_386__35_;
      r_386__34_ <= r_n_386__34_;
      r_386__33_ <= r_n_386__33_;
      r_386__32_ <= r_n_386__32_;
      r_386__31_ <= r_n_386__31_;
      r_386__30_ <= r_n_386__30_;
      r_386__29_ <= r_n_386__29_;
      r_386__28_ <= r_n_386__28_;
      r_386__27_ <= r_n_386__27_;
      r_386__26_ <= r_n_386__26_;
      r_386__25_ <= r_n_386__25_;
      r_386__24_ <= r_n_386__24_;
      r_386__23_ <= r_n_386__23_;
      r_386__22_ <= r_n_386__22_;
      r_386__21_ <= r_n_386__21_;
      r_386__20_ <= r_n_386__20_;
      r_386__19_ <= r_n_386__19_;
      r_386__18_ <= r_n_386__18_;
      r_386__17_ <= r_n_386__17_;
      r_386__16_ <= r_n_386__16_;
      r_386__15_ <= r_n_386__15_;
      r_386__14_ <= r_n_386__14_;
      r_386__13_ <= r_n_386__13_;
      r_386__12_ <= r_n_386__12_;
      r_386__11_ <= r_n_386__11_;
      r_386__10_ <= r_n_386__10_;
      r_386__9_ <= r_n_386__9_;
      r_386__8_ <= r_n_386__8_;
      r_386__7_ <= r_n_386__7_;
      r_386__6_ <= r_n_386__6_;
      r_386__5_ <= r_n_386__5_;
      r_386__4_ <= r_n_386__4_;
      r_386__3_ <= r_n_386__3_;
      r_386__2_ <= r_n_386__2_;
      r_386__1_ <= r_n_386__1_;
      r_386__0_ <= r_n_386__0_;
    end 
    if(N3971) begin
      r_387__63_ <= r_n_387__63_;
      r_387__62_ <= r_n_387__62_;
      r_387__61_ <= r_n_387__61_;
      r_387__60_ <= r_n_387__60_;
      r_387__59_ <= r_n_387__59_;
      r_387__58_ <= r_n_387__58_;
      r_387__57_ <= r_n_387__57_;
      r_387__56_ <= r_n_387__56_;
      r_387__55_ <= r_n_387__55_;
      r_387__54_ <= r_n_387__54_;
      r_387__53_ <= r_n_387__53_;
      r_387__52_ <= r_n_387__52_;
      r_387__51_ <= r_n_387__51_;
      r_387__50_ <= r_n_387__50_;
      r_387__49_ <= r_n_387__49_;
      r_387__48_ <= r_n_387__48_;
      r_387__47_ <= r_n_387__47_;
      r_387__46_ <= r_n_387__46_;
      r_387__45_ <= r_n_387__45_;
      r_387__44_ <= r_n_387__44_;
      r_387__43_ <= r_n_387__43_;
      r_387__42_ <= r_n_387__42_;
      r_387__41_ <= r_n_387__41_;
      r_387__40_ <= r_n_387__40_;
      r_387__39_ <= r_n_387__39_;
      r_387__38_ <= r_n_387__38_;
      r_387__37_ <= r_n_387__37_;
      r_387__36_ <= r_n_387__36_;
      r_387__35_ <= r_n_387__35_;
      r_387__34_ <= r_n_387__34_;
      r_387__33_ <= r_n_387__33_;
      r_387__32_ <= r_n_387__32_;
      r_387__31_ <= r_n_387__31_;
      r_387__30_ <= r_n_387__30_;
      r_387__29_ <= r_n_387__29_;
      r_387__28_ <= r_n_387__28_;
      r_387__27_ <= r_n_387__27_;
      r_387__26_ <= r_n_387__26_;
      r_387__25_ <= r_n_387__25_;
      r_387__24_ <= r_n_387__24_;
      r_387__23_ <= r_n_387__23_;
      r_387__22_ <= r_n_387__22_;
      r_387__21_ <= r_n_387__21_;
      r_387__20_ <= r_n_387__20_;
      r_387__19_ <= r_n_387__19_;
      r_387__18_ <= r_n_387__18_;
      r_387__17_ <= r_n_387__17_;
      r_387__16_ <= r_n_387__16_;
      r_387__15_ <= r_n_387__15_;
      r_387__14_ <= r_n_387__14_;
      r_387__13_ <= r_n_387__13_;
      r_387__12_ <= r_n_387__12_;
      r_387__11_ <= r_n_387__11_;
      r_387__10_ <= r_n_387__10_;
      r_387__9_ <= r_n_387__9_;
      r_387__8_ <= r_n_387__8_;
      r_387__7_ <= r_n_387__7_;
      r_387__6_ <= r_n_387__6_;
      r_387__5_ <= r_n_387__5_;
      r_387__4_ <= r_n_387__4_;
      r_387__3_ <= r_n_387__3_;
      r_387__2_ <= r_n_387__2_;
      r_387__1_ <= r_n_387__1_;
      r_387__0_ <= r_n_387__0_;
    end 
    if(N3972) begin
      r_388__63_ <= r_n_388__63_;
      r_388__62_ <= r_n_388__62_;
      r_388__61_ <= r_n_388__61_;
      r_388__60_ <= r_n_388__60_;
      r_388__59_ <= r_n_388__59_;
      r_388__58_ <= r_n_388__58_;
      r_388__57_ <= r_n_388__57_;
      r_388__56_ <= r_n_388__56_;
      r_388__55_ <= r_n_388__55_;
      r_388__54_ <= r_n_388__54_;
      r_388__53_ <= r_n_388__53_;
      r_388__52_ <= r_n_388__52_;
      r_388__51_ <= r_n_388__51_;
      r_388__50_ <= r_n_388__50_;
      r_388__49_ <= r_n_388__49_;
      r_388__48_ <= r_n_388__48_;
      r_388__47_ <= r_n_388__47_;
      r_388__46_ <= r_n_388__46_;
      r_388__45_ <= r_n_388__45_;
      r_388__44_ <= r_n_388__44_;
      r_388__43_ <= r_n_388__43_;
      r_388__42_ <= r_n_388__42_;
      r_388__41_ <= r_n_388__41_;
      r_388__40_ <= r_n_388__40_;
      r_388__39_ <= r_n_388__39_;
      r_388__38_ <= r_n_388__38_;
      r_388__37_ <= r_n_388__37_;
      r_388__36_ <= r_n_388__36_;
      r_388__35_ <= r_n_388__35_;
      r_388__34_ <= r_n_388__34_;
      r_388__33_ <= r_n_388__33_;
      r_388__32_ <= r_n_388__32_;
      r_388__31_ <= r_n_388__31_;
      r_388__30_ <= r_n_388__30_;
      r_388__29_ <= r_n_388__29_;
      r_388__28_ <= r_n_388__28_;
      r_388__27_ <= r_n_388__27_;
      r_388__26_ <= r_n_388__26_;
      r_388__25_ <= r_n_388__25_;
      r_388__24_ <= r_n_388__24_;
      r_388__23_ <= r_n_388__23_;
      r_388__22_ <= r_n_388__22_;
      r_388__21_ <= r_n_388__21_;
      r_388__20_ <= r_n_388__20_;
      r_388__19_ <= r_n_388__19_;
      r_388__18_ <= r_n_388__18_;
      r_388__17_ <= r_n_388__17_;
      r_388__16_ <= r_n_388__16_;
      r_388__15_ <= r_n_388__15_;
      r_388__14_ <= r_n_388__14_;
      r_388__13_ <= r_n_388__13_;
      r_388__12_ <= r_n_388__12_;
      r_388__11_ <= r_n_388__11_;
      r_388__10_ <= r_n_388__10_;
      r_388__9_ <= r_n_388__9_;
      r_388__8_ <= r_n_388__8_;
      r_388__7_ <= r_n_388__7_;
      r_388__6_ <= r_n_388__6_;
      r_388__5_ <= r_n_388__5_;
      r_388__4_ <= r_n_388__4_;
      r_388__3_ <= r_n_388__3_;
      r_388__2_ <= r_n_388__2_;
      r_388__1_ <= r_n_388__1_;
      r_388__0_ <= r_n_388__0_;
    end 
    if(N3973) begin
      r_389__63_ <= r_n_389__63_;
      r_389__62_ <= r_n_389__62_;
      r_389__61_ <= r_n_389__61_;
      r_389__60_ <= r_n_389__60_;
      r_389__59_ <= r_n_389__59_;
      r_389__58_ <= r_n_389__58_;
      r_389__57_ <= r_n_389__57_;
      r_389__56_ <= r_n_389__56_;
      r_389__55_ <= r_n_389__55_;
      r_389__54_ <= r_n_389__54_;
      r_389__53_ <= r_n_389__53_;
      r_389__52_ <= r_n_389__52_;
      r_389__51_ <= r_n_389__51_;
      r_389__50_ <= r_n_389__50_;
      r_389__49_ <= r_n_389__49_;
      r_389__48_ <= r_n_389__48_;
      r_389__47_ <= r_n_389__47_;
      r_389__46_ <= r_n_389__46_;
      r_389__45_ <= r_n_389__45_;
      r_389__44_ <= r_n_389__44_;
      r_389__43_ <= r_n_389__43_;
      r_389__42_ <= r_n_389__42_;
      r_389__41_ <= r_n_389__41_;
      r_389__40_ <= r_n_389__40_;
      r_389__39_ <= r_n_389__39_;
      r_389__38_ <= r_n_389__38_;
      r_389__37_ <= r_n_389__37_;
      r_389__36_ <= r_n_389__36_;
      r_389__35_ <= r_n_389__35_;
      r_389__34_ <= r_n_389__34_;
      r_389__33_ <= r_n_389__33_;
      r_389__32_ <= r_n_389__32_;
      r_389__31_ <= r_n_389__31_;
      r_389__30_ <= r_n_389__30_;
      r_389__29_ <= r_n_389__29_;
      r_389__28_ <= r_n_389__28_;
      r_389__27_ <= r_n_389__27_;
      r_389__26_ <= r_n_389__26_;
      r_389__25_ <= r_n_389__25_;
      r_389__24_ <= r_n_389__24_;
      r_389__23_ <= r_n_389__23_;
      r_389__22_ <= r_n_389__22_;
      r_389__21_ <= r_n_389__21_;
      r_389__20_ <= r_n_389__20_;
      r_389__19_ <= r_n_389__19_;
      r_389__18_ <= r_n_389__18_;
      r_389__17_ <= r_n_389__17_;
      r_389__16_ <= r_n_389__16_;
      r_389__15_ <= r_n_389__15_;
      r_389__14_ <= r_n_389__14_;
      r_389__13_ <= r_n_389__13_;
      r_389__12_ <= r_n_389__12_;
      r_389__11_ <= r_n_389__11_;
      r_389__10_ <= r_n_389__10_;
      r_389__9_ <= r_n_389__9_;
      r_389__8_ <= r_n_389__8_;
      r_389__7_ <= r_n_389__7_;
      r_389__6_ <= r_n_389__6_;
      r_389__5_ <= r_n_389__5_;
      r_389__4_ <= r_n_389__4_;
      r_389__3_ <= r_n_389__3_;
      r_389__2_ <= r_n_389__2_;
      r_389__1_ <= r_n_389__1_;
      r_389__0_ <= r_n_389__0_;
    end 
    if(N3974) begin
      r_390__63_ <= r_n_390__63_;
      r_390__62_ <= r_n_390__62_;
      r_390__61_ <= r_n_390__61_;
      r_390__60_ <= r_n_390__60_;
      r_390__59_ <= r_n_390__59_;
      r_390__58_ <= r_n_390__58_;
      r_390__57_ <= r_n_390__57_;
      r_390__56_ <= r_n_390__56_;
      r_390__55_ <= r_n_390__55_;
      r_390__54_ <= r_n_390__54_;
      r_390__53_ <= r_n_390__53_;
      r_390__52_ <= r_n_390__52_;
      r_390__51_ <= r_n_390__51_;
      r_390__50_ <= r_n_390__50_;
      r_390__49_ <= r_n_390__49_;
      r_390__48_ <= r_n_390__48_;
      r_390__47_ <= r_n_390__47_;
      r_390__46_ <= r_n_390__46_;
      r_390__45_ <= r_n_390__45_;
      r_390__44_ <= r_n_390__44_;
      r_390__43_ <= r_n_390__43_;
      r_390__42_ <= r_n_390__42_;
      r_390__41_ <= r_n_390__41_;
      r_390__40_ <= r_n_390__40_;
      r_390__39_ <= r_n_390__39_;
      r_390__38_ <= r_n_390__38_;
      r_390__37_ <= r_n_390__37_;
      r_390__36_ <= r_n_390__36_;
      r_390__35_ <= r_n_390__35_;
      r_390__34_ <= r_n_390__34_;
      r_390__33_ <= r_n_390__33_;
      r_390__32_ <= r_n_390__32_;
      r_390__31_ <= r_n_390__31_;
      r_390__30_ <= r_n_390__30_;
      r_390__29_ <= r_n_390__29_;
      r_390__28_ <= r_n_390__28_;
      r_390__27_ <= r_n_390__27_;
      r_390__26_ <= r_n_390__26_;
      r_390__25_ <= r_n_390__25_;
      r_390__24_ <= r_n_390__24_;
      r_390__23_ <= r_n_390__23_;
      r_390__22_ <= r_n_390__22_;
      r_390__21_ <= r_n_390__21_;
      r_390__20_ <= r_n_390__20_;
      r_390__19_ <= r_n_390__19_;
      r_390__18_ <= r_n_390__18_;
      r_390__17_ <= r_n_390__17_;
      r_390__16_ <= r_n_390__16_;
      r_390__15_ <= r_n_390__15_;
      r_390__14_ <= r_n_390__14_;
      r_390__13_ <= r_n_390__13_;
      r_390__12_ <= r_n_390__12_;
      r_390__11_ <= r_n_390__11_;
      r_390__10_ <= r_n_390__10_;
      r_390__9_ <= r_n_390__9_;
      r_390__8_ <= r_n_390__8_;
      r_390__7_ <= r_n_390__7_;
      r_390__6_ <= r_n_390__6_;
      r_390__5_ <= r_n_390__5_;
      r_390__4_ <= r_n_390__4_;
      r_390__3_ <= r_n_390__3_;
      r_390__2_ <= r_n_390__2_;
      r_390__1_ <= r_n_390__1_;
      r_390__0_ <= r_n_390__0_;
    end 
    if(N3975) begin
      r_391__63_ <= r_n_391__63_;
      r_391__62_ <= r_n_391__62_;
      r_391__61_ <= r_n_391__61_;
      r_391__60_ <= r_n_391__60_;
      r_391__59_ <= r_n_391__59_;
      r_391__58_ <= r_n_391__58_;
      r_391__57_ <= r_n_391__57_;
      r_391__56_ <= r_n_391__56_;
      r_391__55_ <= r_n_391__55_;
      r_391__54_ <= r_n_391__54_;
      r_391__53_ <= r_n_391__53_;
      r_391__52_ <= r_n_391__52_;
      r_391__51_ <= r_n_391__51_;
      r_391__50_ <= r_n_391__50_;
      r_391__49_ <= r_n_391__49_;
      r_391__48_ <= r_n_391__48_;
      r_391__47_ <= r_n_391__47_;
      r_391__46_ <= r_n_391__46_;
      r_391__45_ <= r_n_391__45_;
      r_391__44_ <= r_n_391__44_;
      r_391__43_ <= r_n_391__43_;
      r_391__42_ <= r_n_391__42_;
      r_391__41_ <= r_n_391__41_;
      r_391__40_ <= r_n_391__40_;
      r_391__39_ <= r_n_391__39_;
      r_391__38_ <= r_n_391__38_;
      r_391__37_ <= r_n_391__37_;
      r_391__36_ <= r_n_391__36_;
      r_391__35_ <= r_n_391__35_;
      r_391__34_ <= r_n_391__34_;
      r_391__33_ <= r_n_391__33_;
      r_391__32_ <= r_n_391__32_;
      r_391__31_ <= r_n_391__31_;
      r_391__30_ <= r_n_391__30_;
      r_391__29_ <= r_n_391__29_;
      r_391__28_ <= r_n_391__28_;
      r_391__27_ <= r_n_391__27_;
      r_391__26_ <= r_n_391__26_;
      r_391__25_ <= r_n_391__25_;
      r_391__24_ <= r_n_391__24_;
      r_391__23_ <= r_n_391__23_;
      r_391__22_ <= r_n_391__22_;
      r_391__21_ <= r_n_391__21_;
      r_391__20_ <= r_n_391__20_;
      r_391__19_ <= r_n_391__19_;
      r_391__18_ <= r_n_391__18_;
      r_391__17_ <= r_n_391__17_;
      r_391__16_ <= r_n_391__16_;
      r_391__15_ <= r_n_391__15_;
      r_391__14_ <= r_n_391__14_;
      r_391__13_ <= r_n_391__13_;
      r_391__12_ <= r_n_391__12_;
      r_391__11_ <= r_n_391__11_;
      r_391__10_ <= r_n_391__10_;
      r_391__9_ <= r_n_391__9_;
      r_391__8_ <= r_n_391__8_;
      r_391__7_ <= r_n_391__7_;
      r_391__6_ <= r_n_391__6_;
      r_391__5_ <= r_n_391__5_;
      r_391__4_ <= r_n_391__4_;
      r_391__3_ <= r_n_391__3_;
      r_391__2_ <= r_n_391__2_;
      r_391__1_ <= r_n_391__1_;
      r_391__0_ <= r_n_391__0_;
    end 
    if(N3976) begin
      r_392__63_ <= r_n_392__63_;
      r_392__62_ <= r_n_392__62_;
      r_392__61_ <= r_n_392__61_;
      r_392__60_ <= r_n_392__60_;
      r_392__59_ <= r_n_392__59_;
      r_392__58_ <= r_n_392__58_;
      r_392__57_ <= r_n_392__57_;
      r_392__56_ <= r_n_392__56_;
      r_392__55_ <= r_n_392__55_;
      r_392__54_ <= r_n_392__54_;
      r_392__53_ <= r_n_392__53_;
      r_392__52_ <= r_n_392__52_;
      r_392__51_ <= r_n_392__51_;
      r_392__50_ <= r_n_392__50_;
      r_392__49_ <= r_n_392__49_;
      r_392__48_ <= r_n_392__48_;
      r_392__47_ <= r_n_392__47_;
      r_392__46_ <= r_n_392__46_;
      r_392__45_ <= r_n_392__45_;
      r_392__44_ <= r_n_392__44_;
      r_392__43_ <= r_n_392__43_;
      r_392__42_ <= r_n_392__42_;
      r_392__41_ <= r_n_392__41_;
      r_392__40_ <= r_n_392__40_;
      r_392__39_ <= r_n_392__39_;
      r_392__38_ <= r_n_392__38_;
      r_392__37_ <= r_n_392__37_;
      r_392__36_ <= r_n_392__36_;
      r_392__35_ <= r_n_392__35_;
      r_392__34_ <= r_n_392__34_;
      r_392__33_ <= r_n_392__33_;
      r_392__32_ <= r_n_392__32_;
      r_392__31_ <= r_n_392__31_;
      r_392__30_ <= r_n_392__30_;
      r_392__29_ <= r_n_392__29_;
      r_392__28_ <= r_n_392__28_;
      r_392__27_ <= r_n_392__27_;
      r_392__26_ <= r_n_392__26_;
      r_392__25_ <= r_n_392__25_;
      r_392__24_ <= r_n_392__24_;
      r_392__23_ <= r_n_392__23_;
      r_392__22_ <= r_n_392__22_;
      r_392__21_ <= r_n_392__21_;
      r_392__20_ <= r_n_392__20_;
      r_392__19_ <= r_n_392__19_;
      r_392__18_ <= r_n_392__18_;
      r_392__17_ <= r_n_392__17_;
      r_392__16_ <= r_n_392__16_;
      r_392__15_ <= r_n_392__15_;
      r_392__14_ <= r_n_392__14_;
      r_392__13_ <= r_n_392__13_;
      r_392__12_ <= r_n_392__12_;
      r_392__11_ <= r_n_392__11_;
      r_392__10_ <= r_n_392__10_;
      r_392__9_ <= r_n_392__9_;
      r_392__8_ <= r_n_392__8_;
      r_392__7_ <= r_n_392__7_;
      r_392__6_ <= r_n_392__6_;
      r_392__5_ <= r_n_392__5_;
      r_392__4_ <= r_n_392__4_;
      r_392__3_ <= r_n_392__3_;
      r_392__2_ <= r_n_392__2_;
      r_392__1_ <= r_n_392__1_;
      r_392__0_ <= r_n_392__0_;
    end 
    if(N3977) begin
      r_393__63_ <= r_n_393__63_;
      r_393__62_ <= r_n_393__62_;
      r_393__61_ <= r_n_393__61_;
      r_393__60_ <= r_n_393__60_;
      r_393__59_ <= r_n_393__59_;
      r_393__58_ <= r_n_393__58_;
      r_393__57_ <= r_n_393__57_;
      r_393__56_ <= r_n_393__56_;
      r_393__55_ <= r_n_393__55_;
      r_393__54_ <= r_n_393__54_;
      r_393__53_ <= r_n_393__53_;
      r_393__52_ <= r_n_393__52_;
      r_393__51_ <= r_n_393__51_;
      r_393__50_ <= r_n_393__50_;
      r_393__49_ <= r_n_393__49_;
      r_393__48_ <= r_n_393__48_;
      r_393__47_ <= r_n_393__47_;
      r_393__46_ <= r_n_393__46_;
      r_393__45_ <= r_n_393__45_;
      r_393__44_ <= r_n_393__44_;
      r_393__43_ <= r_n_393__43_;
      r_393__42_ <= r_n_393__42_;
      r_393__41_ <= r_n_393__41_;
      r_393__40_ <= r_n_393__40_;
      r_393__39_ <= r_n_393__39_;
      r_393__38_ <= r_n_393__38_;
      r_393__37_ <= r_n_393__37_;
      r_393__36_ <= r_n_393__36_;
      r_393__35_ <= r_n_393__35_;
      r_393__34_ <= r_n_393__34_;
      r_393__33_ <= r_n_393__33_;
      r_393__32_ <= r_n_393__32_;
      r_393__31_ <= r_n_393__31_;
      r_393__30_ <= r_n_393__30_;
      r_393__29_ <= r_n_393__29_;
      r_393__28_ <= r_n_393__28_;
      r_393__27_ <= r_n_393__27_;
      r_393__26_ <= r_n_393__26_;
      r_393__25_ <= r_n_393__25_;
      r_393__24_ <= r_n_393__24_;
      r_393__23_ <= r_n_393__23_;
      r_393__22_ <= r_n_393__22_;
      r_393__21_ <= r_n_393__21_;
      r_393__20_ <= r_n_393__20_;
      r_393__19_ <= r_n_393__19_;
      r_393__18_ <= r_n_393__18_;
      r_393__17_ <= r_n_393__17_;
      r_393__16_ <= r_n_393__16_;
      r_393__15_ <= r_n_393__15_;
      r_393__14_ <= r_n_393__14_;
      r_393__13_ <= r_n_393__13_;
      r_393__12_ <= r_n_393__12_;
      r_393__11_ <= r_n_393__11_;
      r_393__10_ <= r_n_393__10_;
      r_393__9_ <= r_n_393__9_;
      r_393__8_ <= r_n_393__8_;
      r_393__7_ <= r_n_393__7_;
      r_393__6_ <= r_n_393__6_;
      r_393__5_ <= r_n_393__5_;
      r_393__4_ <= r_n_393__4_;
      r_393__3_ <= r_n_393__3_;
      r_393__2_ <= r_n_393__2_;
      r_393__1_ <= r_n_393__1_;
      r_393__0_ <= r_n_393__0_;
    end 
    if(N3978) begin
      r_394__63_ <= r_n_394__63_;
      r_394__62_ <= r_n_394__62_;
      r_394__61_ <= r_n_394__61_;
      r_394__60_ <= r_n_394__60_;
      r_394__59_ <= r_n_394__59_;
      r_394__58_ <= r_n_394__58_;
      r_394__57_ <= r_n_394__57_;
      r_394__56_ <= r_n_394__56_;
      r_394__55_ <= r_n_394__55_;
      r_394__54_ <= r_n_394__54_;
      r_394__53_ <= r_n_394__53_;
      r_394__52_ <= r_n_394__52_;
      r_394__51_ <= r_n_394__51_;
      r_394__50_ <= r_n_394__50_;
      r_394__49_ <= r_n_394__49_;
      r_394__48_ <= r_n_394__48_;
      r_394__47_ <= r_n_394__47_;
      r_394__46_ <= r_n_394__46_;
      r_394__45_ <= r_n_394__45_;
      r_394__44_ <= r_n_394__44_;
      r_394__43_ <= r_n_394__43_;
      r_394__42_ <= r_n_394__42_;
      r_394__41_ <= r_n_394__41_;
      r_394__40_ <= r_n_394__40_;
      r_394__39_ <= r_n_394__39_;
      r_394__38_ <= r_n_394__38_;
      r_394__37_ <= r_n_394__37_;
      r_394__36_ <= r_n_394__36_;
      r_394__35_ <= r_n_394__35_;
      r_394__34_ <= r_n_394__34_;
      r_394__33_ <= r_n_394__33_;
      r_394__32_ <= r_n_394__32_;
      r_394__31_ <= r_n_394__31_;
      r_394__30_ <= r_n_394__30_;
      r_394__29_ <= r_n_394__29_;
      r_394__28_ <= r_n_394__28_;
      r_394__27_ <= r_n_394__27_;
      r_394__26_ <= r_n_394__26_;
      r_394__25_ <= r_n_394__25_;
      r_394__24_ <= r_n_394__24_;
      r_394__23_ <= r_n_394__23_;
      r_394__22_ <= r_n_394__22_;
      r_394__21_ <= r_n_394__21_;
      r_394__20_ <= r_n_394__20_;
      r_394__19_ <= r_n_394__19_;
      r_394__18_ <= r_n_394__18_;
      r_394__17_ <= r_n_394__17_;
      r_394__16_ <= r_n_394__16_;
      r_394__15_ <= r_n_394__15_;
      r_394__14_ <= r_n_394__14_;
      r_394__13_ <= r_n_394__13_;
      r_394__12_ <= r_n_394__12_;
      r_394__11_ <= r_n_394__11_;
      r_394__10_ <= r_n_394__10_;
      r_394__9_ <= r_n_394__9_;
      r_394__8_ <= r_n_394__8_;
      r_394__7_ <= r_n_394__7_;
      r_394__6_ <= r_n_394__6_;
      r_394__5_ <= r_n_394__5_;
      r_394__4_ <= r_n_394__4_;
      r_394__3_ <= r_n_394__3_;
      r_394__2_ <= r_n_394__2_;
      r_394__1_ <= r_n_394__1_;
      r_394__0_ <= r_n_394__0_;
    end 
    if(N3979) begin
      r_395__63_ <= r_n_395__63_;
      r_395__62_ <= r_n_395__62_;
      r_395__61_ <= r_n_395__61_;
      r_395__60_ <= r_n_395__60_;
      r_395__59_ <= r_n_395__59_;
      r_395__58_ <= r_n_395__58_;
      r_395__57_ <= r_n_395__57_;
      r_395__56_ <= r_n_395__56_;
      r_395__55_ <= r_n_395__55_;
      r_395__54_ <= r_n_395__54_;
      r_395__53_ <= r_n_395__53_;
      r_395__52_ <= r_n_395__52_;
      r_395__51_ <= r_n_395__51_;
      r_395__50_ <= r_n_395__50_;
      r_395__49_ <= r_n_395__49_;
      r_395__48_ <= r_n_395__48_;
      r_395__47_ <= r_n_395__47_;
      r_395__46_ <= r_n_395__46_;
      r_395__45_ <= r_n_395__45_;
      r_395__44_ <= r_n_395__44_;
      r_395__43_ <= r_n_395__43_;
      r_395__42_ <= r_n_395__42_;
      r_395__41_ <= r_n_395__41_;
      r_395__40_ <= r_n_395__40_;
      r_395__39_ <= r_n_395__39_;
      r_395__38_ <= r_n_395__38_;
      r_395__37_ <= r_n_395__37_;
      r_395__36_ <= r_n_395__36_;
      r_395__35_ <= r_n_395__35_;
      r_395__34_ <= r_n_395__34_;
      r_395__33_ <= r_n_395__33_;
      r_395__32_ <= r_n_395__32_;
      r_395__31_ <= r_n_395__31_;
      r_395__30_ <= r_n_395__30_;
      r_395__29_ <= r_n_395__29_;
      r_395__28_ <= r_n_395__28_;
      r_395__27_ <= r_n_395__27_;
      r_395__26_ <= r_n_395__26_;
      r_395__25_ <= r_n_395__25_;
      r_395__24_ <= r_n_395__24_;
      r_395__23_ <= r_n_395__23_;
      r_395__22_ <= r_n_395__22_;
      r_395__21_ <= r_n_395__21_;
      r_395__20_ <= r_n_395__20_;
      r_395__19_ <= r_n_395__19_;
      r_395__18_ <= r_n_395__18_;
      r_395__17_ <= r_n_395__17_;
      r_395__16_ <= r_n_395__16_;
      r_395__15_ <= r_n_395__15_;
      r_395__14_ <= r_n_395__14_;
      r_395__13_ <= r_n_395__13_;
      r_395__12_ <= r_n_395__12_;
      r_395__11_ <= r_n_395__11_;
      r_395__10_ <= r_n_395__10_;
      r_395__9_ <= r_n_395__9_;
      r_395__8_ <= r_n_395__8_;
      r_395__7_ <= r_n_395__7_;
      r_395__6_ <= r_n_395__6_;
      r_395__5_ <= r_n_395__5_;
      r_395__4_ <= r_n_395__4_;
      r_395__3_ <= r_n_395__3_;
      r_395__2_ <= r_n_395__2_;
      r_395__1_ <= r_n_395__1_;
      r_395__0_ <= r_n_395__0_;
    end 
    if(N3980) begin
      r_396__63_ <= r_n_396__63_;
      r_396__62_ <= r_n_396__62_;
      r_396__61_ <= r_n_396__61_;
      r_396__60_ <= r_n_396__60_;
      r_396__59_ <= r_n_396__59_;
      r_396__58_ <= r_n_396__58_;
      r_396__57_ <= r_n_396__57_;
      r_396__56_ <= r_n_396__56_;
      r_396__55_ <= r_n_396__55_;
      r_396__54_ <= r_n_396__54_;
      r_396__53_ <= r_n_396__53_;
      r_396__52_ <= r_n_396__52_;
      r_396__51_ <= r_n_396__51_;
      r_396__50_ <= r_n_396__50_;
      r_396__49_ <= r_n_396__49_;
      r_396__48_ <= r_n_396__48_;
      r_396__47_ <= r_n_396__47_;
      r_396__46_ <= r_n_396__46_;
      r_396__45_ <= r_n_396__45_;
      r_396__44_ <= r_n_396__44_;
      r_396__43_ <= r_n_396__43_;
      r_396__42_ <= r_n_396__42_;
      r_396__41_ <= r_n_396__41_;
      r_396__40_ <= r_n_396__40_;
      r_396__39_ <= r_n_396__39_;
      r_396__38_ <= r_n_396__38_;
      r_396__37_ <= r_n_396__37_;
      r_396__36_ <= r_n_396__36_;
      r_396__35_ <= r_n_396__35_;
      r_396__34_ <= r_n_396__34_;
      r_396__33_ <= r_n_396__33_;
      r_396__32_ <= r_n_396__32_;
      r_396__31_ <= r_n_396__31_;
      r_396__30_ <= r_n_396__30_;
      r_396__29_ <= r_n_396__29_;
      r_396__28_ <= r_n_396__28_;
      r_396__27_ <= r_n_396__27_;
      r_396__26_ <= r_n_396__26_;
      r_396__25_ <= r_n_396__25_;
      r_396__24_ <= r_n_396__24_;
      r_396__23_ <= r_n_396__23_;
      r_396__22_ <= r_n_396__22_;
      r_396__21_ <= r_n_396__21_;
      r_396__20_ <= r_n_396__20_;
      r_396__19_ <= r_n_396__19_;
      r_396__18_ <= r_n_396__18_;
      r_396__17_ <= r_n_396__17_;
      r_396__16_ <= r_n_396__16_;
      r_396__15_ <= r_n_396__15_;
      r_396__14_ <= r_n_396__14_;
      r_396__13_ <= r_n_396__13_;
      r_396__12_ <= r_n_396__12_;
      r_396__11_ <= r_n_396__11_;
      r_396__10_ <= r_n_396__10_;
      r_396__9_ <= r_n_396__9_;
      r_396__8_ <= r_n_396__8_;
      r_396__7_ <= r_n_396__7_;
      r_396__6_ <= r_n_396__6_;
      r_396__5_ <= r_n_396__5_;
      r_396__4_ <= r_n_396__4_;
      r_396__3_ <= r_n_396__3_;
      r_396__2_ <= r_n_396__2_;
      r_396__1_ <= r_n_396__1_;
      r_396__0_ <= r_n_396__0_;
    end 
    if(N3981) begin
      r_397__63_ <= r_n_397__63_;
      r_397__62_ <= r_n_397__62_;
      r_397__61_ <= r_n_397__61_;
      r_397__60_ <= r_n_397__60_;
      r_397__59_ <= r_n_397__59_;
      r_397__58_ <= r_n_397__58_;
      r_397__57_ <= r_n_397__57_;
      r_397__56_ <= r_n_397__56_;
      r_397__55_ <= r_n_397__55_;
      r_397__54_ <= r_n_397__54_;
      r_397__53_ <= r_n_397__53_;
      r_397__52_ <= r_n_397__52_;
      r_397__51_ <= r_n_397__51_;
      r_397__50_ <= r_n_397__50_;
      r_397__49_ <= r_n_397__49_;
      r_397__48_ <= r_n_397__48_;
      r_397__47_ <= r_n_397__47_;
      r_397__46_ <= r_n_397__46_;
      r_397__45_ <= r_n_397__45_;
      r_397__44_ <= r_n_397__44_;
      r_397__43_ <= r_n_397__43_;
      r_397__42_ <= r_n_397__42_;
      r_397__41_ <= r_n_397__41_;
      r_397__40_ <= r_n_397__40_;
      r_397__39_ <= r_n_397__39_;
      r_397__38_ <= r_n_397__38_;
      r_397__37_ <= r_n_397__37_;
      r_397__36_ <= r_n_397__36_;
      r_397__35_ <= r_n_397__35_;
      r_397__34_ <= r_n_397__34_;
      r_397__33_ <= r_n_397__33_;
      r_397__32_ <= r_n_397__32_;
      r_397__31_ <= r_n_397__31_;
      r_397__30_ <= r_n_397__30_;
      r_397__29_ <= r_n_397__29_;
      r_397__28_ <= r_n_397__28_;
      r_397__27_ <= r_n_397__27_;
      r_397__26_ <= r_n_397__26_;
      r_397__25_ <= r_n_397__25_;
      r_397__24_ <= r_n_397__24_;
      r_397__23_ <= r_n_397__23_;
      r_397__22_ <= r_n_397__22_;
      r_397__21_ <= r_n_397__21_;
      r_397__20_ <= r_n_397__20_;
      r_397__19_ <= r_n_397__19_;
      r_397__18_ <= r_n_397__18_;
      r_397__17_ <= r_n_397__17_;
      r_397__16_ <= r_n_397__16_;
      r_397__15_ <= r_n_397__15_;
      r_397__14_ <= r_n_397__14_;
      r_397__13_ <= r_n_397__13_;
      r_397__12_ <= r_n_397__12_;
      r_397__11_ <= r_n_397__11_;
      r_397__10_ <= r_n_397__10_;
      r_397__9_ <= r_n_397__9_;
      r_397__8_ <= r_n_397__8_;
      r_397__7_ <= r_n_397__7_;
      r_397__6_ <= r_n_397__6_;
      r_397__5_ <= r_n_397__5_;
      r_397__4_ <= r_n_397__4_;
      r_397__3_ <= r_n_397__3_;
      r_397__2_ <= r_n_397__2_;
      r_397__1_ <= r_n_397__1_;
      r_397__0_ <= r_n_397__0_;
    end 
    if(N3982) begin
      r_398__63_ <= r_n_398__63_;
      r_398__62_ <= r_n_398__62_;
      r_398__61_ <= r_n_398__61_;
      r_398__60_ <= r_n_398__60_;
      r_398__59_ <= r_n_398__59_;
      r_398__58_ <= r_n_398__58_;
      r_398__57_ <= r_n_398__57_;
      r_398__56_ <= r_n_398__56_;
      r_398__55_ <= r_n_398__55_;
      r_398__54_ <= r_n_398__54_;
      r_398__53_ <= r_n_398__53_;
      r_398__52_ <= r_n_398__52_;
      r_398__51_ <= r_n_398__51_;
      r_398__50_ <= r_n_398__50_;
      r_398__49_ <= r_n_398__49_;
      r_398__48_ <= r_n_398__48_;
      r_398__47_ <= r_n_398__47_;
      r_398__46_ <= r_n_398__46_;
      r_398__45_ <= r_n_398__45_;
      r_398__44_ <= r_n_398__44_;
      r_398__43_ <= r_n_398__43_;
      r_398__42_ <= r_n_398__42_;
      r_398__41_ <= r_n_398__41_;
      r_398__40_ <= r_n_398__40_;
      r_398__39_ <= r_n_398__39_;
      r_398__38_ <= r_n_398__38_;
      r_398__37_ <= r_n_398__37_;
      r_398__36_ <= r_n_398__36_;
      r_398__35_ <= r_n_398__35_;
      r_398__34_ <= r_n_398__34_;
      r_398__33_ <= r_n_398__33_;
      r_398__32_ <= r_n_398__32_;
      r_398__31_ <= r_n_398__31_;
      r_398__30_ <= r_n_398__30_;
      r_398__29_ <= r_n_398__29_;
      r_398__28_ <= r_n_398__28_;
      r_398__27_ <= r_n_398__27_;
      r_398__26_ <= r_n_398__26_;
      r_398__25_ <= r_n_398__25_;
      r_398__24_ <= r_n_398__24_;
      r_398__23_ <= r_n_398__23_;
      r_398__22_ <= r_n_398__22_;
      r_398__21_ <= r_n_398__21_;
      r_398__20_ <= r_n_398__20_;
      r_398__19_ <= r_n_398__19_;
      r_398__18_ <= r_n_398__18_;
      r_398__17_ <= r_n_398__17_;
      r_398__16_ <= r_n_398__16_;
      r_398__15_ <= r_n_398__15_;
      r_398__14_ <= r_n_398__14_;
      r_398__13_ <= r_n_398__13_;
      r_398__12_ <= r_n_398__12_;
      r_398__11_ <= r_n_398__11_;
      r_398__10_ <= r_n_398__10_;
      r_398__9_ <= r_n_398__9_;
      r_398__8_ <= r_n_398__8_;
      r_398__7_ <= r_n_398__7_;
      r_398__6_ <= r_n_398__6_;
      r_398__5_ <= r_n_398__5_;
      r_398__4_ <= r_n_398__4_;
      r_398__3_ <= r_n_398__3_;
      r_398__2_ <= r_n_398__2_;
      r_398__1_ <= r_n_398__1_;
      r_398__0_ <= r_n_398__0_;
    end 
    if(N3983) begin
      r_399__63_ <= r_n_399__63_;
      r_399__62_ <= r_n_399__62_;
      r_399__61_ <= r_n_399__61_;
      r_399__60_ <= r_n_399__60_;
      r_399__59_ <= r_n_399__59_;
      r_399__58_ <= r_n_399__58_;
      r_399__57_ <= r_n_399__57_;
      r_399__56_ <= r_n_399__56_;
      r_399__55_ <= r_n_399__55_;
      r_399__54_ <= r_n_399__54_;
      r_399__53_ <= r_n_399__53_;
      r_399__52_ <= r_n_399__52_;
      r_399__51_ <= r_n_399__51_;
      r_399__50_ <= r_n_399__50_;
      r_399__49_ <= r_n_399__49_;
      r_399__48_ <= r_n_399__48_;
      r_399__47_ <= r_n_399__47_;
      r_399__46_ <= r_n_399__46_;
      r_399__45_ <= r_n_399__45_;
      r_399__44_ <= r_n_399__44_;
      r_399__43_ <= r_n_399__43_;
      r_399__42_ <= r_n_399__42_;
      r_399__41_ <= r_n_399__41_;
      r_399__40_ <= r_n_399__40_;
      r_399__39_ <= r_n_399__39_;
      r_399__38_ <= r_n_399__38_;
      r_399__37_ <= r_n_399__37_;
      r_399__36_ <= r_n_399__36_;
      r_399__35_ <= r_n_399__35_;
      r_399__34_ <= r_n_399__34_;
      r_399__33_ <= r_n_399__33_;
      r_399__32_ <= r_n_399__32_;
      r_399__31_ <= r_n_399__31_;
      r_399__30_ <= r_n_399__30_;
      r_399__29_ <= r_n_399__29_;
      r_399__28_ <= r_n_399__28_;
      r_399__27_ <= r_n_399__27_;
      r_399__26_ <= r_n_399__26_;
      r_399__25_ <= r_n_399__25_;
      r_399__24_ <= r_n_399__24_;
      r_399__23_ <= r_n_399__23_;
      r_399__22_ <= r_n_399__22_;
      r_399__21_ <= r_n_399__21_;
      r_399__20_ <= r_n_399__20_;
      r_399__19_ <= r_n_399__19_;
      r_399__18_ <= r_n_399__18_;
      r_399__17_ <= r_n_399__17_;
      r_399__16_ <= r_n_399__16_;
      r_399__15_ <= r_n_399__15_;
      r_399__14_ <= r_n_399__14_;
      r_399__13_ <= r_n_399__13_;
      r_399__12_ <= r_n_399__12_;
      r_399__11_ <= r_n_399__11_;
      r_399__10_ <= r_n_399__10_;
      r_399__9_ <= r_n_399__9_;
      r_399__8_ <= r_n_399__8_;
      r_399__7_ <= r_n_399__7_;
      r_399__6_ <= r_n_399__6_;
      r_399__5_ <= r_n_399__5_;
      r_399__4_ <= r_n_399__4_;
      r_399__3_ <= r_n_399__3_;
      r_399__2_ <= r_n_399__2_;
      r_399__1_ <= r_n_399__1_;
      r_399__0_ <= r_n_399__0_;
    end 
    if(N3984) begin
      r_400__63_ <= r_n_400__63_;
      r_400__62_ <= r_n_400__62_;
      r_400__61_ <= r_n_400__61_;
      r_400__60_ <= r_n_400__60_;
      r_400__59_ <= r_n_400__59_;
      r_400__58_ <= r_n_400__58_;
      r_400__57_ <= r_n_400__57_;
      r_400__56_ <= r_n_400__56_;
      r_400__55_ <= r_n_400__55_;
      r_400__54_ <= r_n_400__54_;
      r_400__53_ <= r_n_400__53_;
      r_400__52_ <= r_n_400__52_;
      r_400__51_ <= r_n_400__51_;
      r_400__50_ <= r_n_400__50_;
      r_400__49_ <= r_n_400__49_;
      r_400__48_ <= r_n_400__48_;
      r_400__47_ <= r_n_400__47_;
      r_400__46_ <= r_n_400__46_;
      r_400__45_ <= r_n_400__45_;
      r_400__44_ <= r_n_400__44_;
      r_400__43_ <= r_n_400__43_;
      r_400__42_ <= r_n_400__42_;
      r_400__41_ <= r_n_400__41_;
      r_400__40_ <= r_n_400__40_;
      r_400__39_ <= r_n_400__39_;
      r_400__38_ <= r_n_400__38_;
      r_400__37_ <= r_n_400__37_;
      r_400__36_ <= r_n_400__36_;
      r_400__35_ <= r_n_400__35_;
      r_400__34_ <= r_n_400__34_;
      r_400__33_ <= r_n_400__33_;
      r_400__32_ <= r_n_400__32_;
      r_400__31_ <= r_n_400__31_;
      r_400__30_ <= r_n_400__30_;
      r_400__29_ <= r_n_400__29_;
      r_400__28_ <= r_n_400__28_;
      r_400__27_ <= r_n_400__27_;
      r_400__26_ <= r_n_400__26_;
      r_400__25_ <= r_n_400__25_;
      r_400__24_ <= r_n_400__24_;
      r_400__23_ <= r_n_400__23_;
      r_400__22_ <= r_n_400__22_;
      r_400__21_ <= r_n_400__21_;
      r_400__20_ <= r_n_400__20_;
      r_400__19_ <= r_n_400__19_;
      r_400__18_ <= r_n_400__18_;
      r_400__17_ <= r_n_400__17_;
      r_400__16_ <= r_n_400__16_;
      r_400__15_ <= r_n_400__15_;
      r_400__14_ <= r_n_400__14_;
      r_400__13_ <= r_n_400__13_;
      r_400__12_ <= r_n_400__12_;
      r_400__11_ <= r_n_400__11_;
      r_400__10_ <= r_n_400__10_;
      r_400__9_ <= r_n_400__9_;
      r_400__8_ <= r_n_400__8_;
      r_400__7_ <= r_n_400__7_;
      r_400__6_ <= r_n_400__6_;
      r_400__5_ <= r_n_400__5_;
      r_400__4_ <= r_n_400__4_;
      r_400__3_ <= r_n_400__3_;
      r_400__2_ <= r_n_400__2_;
      r_400__1_ <= r_n_400__1_;
      r_400__0_ <= r_n_400__0_;
    end 
    if(N3985) begin
      r_401__63_ <= r_n_401__63_;
      r_401__62_ <= r_n_401__62_;
      r_401__61_ <= r_n_401__61_;
      r_401__60_ <= r_n_401__60_;
      r_401__59_ <= r_n_401__59_;
      r_401__58_ <= r_n_401__58_;
      r_401__57_ <= r_n_401__57_;
      r_401__56_ <= r_n_401__56_;
      r_401__55_ <= r_n_401__55_;
      r_401__54_ <= r_n_401__54_;
      r_401__53_ <= r_n_401__53_;
      r_401__52_ <= r_n_401__52_;
      r_401__51_ <= r_n_401__51_;
      r_401__50_ <= r_n_401__50_;
      r_401__49_ <= r_n_401__49_;
      r_401__48_ <= r_n_401__48_;
      r_401__47_ <= r_n_401__47_;
      r_401__46_ <= r_n_401__46_;
      r_401__45_ <= r_n_401__45_;
      r_401__44_ <= r_n_401__44_;
      r_401__43_ <= r_n_401__43_;
      r_401__42_ <= r_n_401__42_;
      r_401__41_ <= r_n_401__41_;
      r_401__40_ <= r_n_401__40_;
      r_401__39_ <= r_n_401__39_;
      r_401__38_ <= r_n_401__38_;
      r_401__37_ <= r_n_401__37_;
      r_401__36_ <= r_n_401__36_;
      r_401__35_ <= r_n_401__35_;
      r_401__34_ <= r_n_401__34_;
      r_401__33_ <= r_n_401__33_;
      r_401__32_ <= r_n_401__32_;
      r_401__31_ <= r_n_401__31_;
      r_401__30_ <= r_n_401__30_;
      r_401__29_ <= r_n_401__29_;
      r_401__28_ <= r_n_401__28_;
      r_401__27_ <= r_n_401__27_;
      r_401__26_ <= r_n_401__26_;
      r_401__25_ <= r_n_401__25_;
      r_401__24_ <= r_n_401__24_;
      r_401__23_ <= r_n_401__23_;
      r_401__22_ <= r_n_401__22_;
      r_401__21_ <= r_n_401__21_;
      r_401__20_ <= r_n_401__20_;
      r_401__19_ <= r_n_401__19_;
      r_401__18_ <= r_n_401__18_;
      r_401__17_ <= r_n_401__17_;
      r_401__16_ <= r_n_401__16_;
      r_401__15_ <= r_n_401__15_;
      r_401__14_ <= r_n_401__14_;
      r_401__13_ <= r_n_401__13_;
      r_401__12_ <= r_n_401__12_;
      r_401__11_ <= r_n_401__11_;
      r_401__10_ <= r_n_401__10_;
      r_401__9_ <= r_n_401__9_;
      r_401__8_ <= r_n_401__8_;
      r_401__7_ <= r_n_401__7_;
      r_401__6_ <= r_n_401__6_;
      r_401__5_ <= r_n_401__5_;
      r_401__4_ <= r_n_401__4_;
      r_401__3_ <= r_n_401__3_;
      r_401__2_ <= r_n_401__2_;
      r_401__1_ <= r_n_401__1_;
      r_401__0_ <= r_n_401__0_;
    end 
    if(N3986) begin
      r_402__63_ <= r_n_402__63_;
      r_402__62_ <= r_n_402__62_;
      r_402__61_ <= r_n_402__61_;
      r_402__60_ <= r_n_402__60_;
      r_402__59_ <= r_n_402__59_;
      r_402__58_ <= r_n_402__58_;
      r_402__57_ <= r_n_402__57_;
      r_402__56_ <= r_n_402__56_;
      r_402__55_ <= r_n_402__55_;
      r_402__54_ <= r_n_402__54_;
      r_402__53_ <= r_n_402__53_;
      r_402__52_ <= r_n_402__52_;
      r_402__51_ <= r_n_402__51_;
      r_402__50_ <= r_n_402__50_;
      r_402__49_ <= r_n_402__49_;
      r_402__48_ <= r_n_402__48_;
      r_402__47_ <= r_n_402__47_;
      r_402__46_ <= r_n_402__46_;
      r_402__45_ <= r_n_402__45_;
      r_402__44_ <= r_n_402__44_;
      r_402__43_ <= r_n_402__43_;
      r_402__42_ <= r_n_402__42_;
      r_402__41_ <= r_n_402__41_;
      r_402__40_ <= r_n_402__40_;
      r_402__39_ <= r_n_402__39_;
      r_402__38_ <= r_n_402__38_;
      r_402__37_ <= r_n_402__37_;
      r_402__36_ <= r_n_402__36_;
      r_402__35_ <= r_n_402__35_;
      r_402__34_ <= r_n_402__34_;
      r_402__33_ <= r_n_402__33_;
      r_402__32_ <= r_n_402__32_;
      r_402__31_ <= r_n_402__31_;
      r_402__30_ <= r_n_402__30_;
      r_402__29_ <= r_n_402__29_;
      r_402__28_ <= r_n_402__28_;
      r_402__27_ <= r_n_402__27_;
      r_402__26_ <= r_n_402__26_;
      r_402__25_ <= r_n_402__25_;
      r_402__24_ <= r_n_402__24_;
      r_402__23_ <= r_n_402__23_;
      r_402__22_ <= r_n_402__22_;
      r_402__21_ <= r_n_402__21_;
      r_402__20_ <= r_n_402__20_;
      r_402__19_ <= r_n_402__19_;
      r_402__18_ <= r_n_402__18_;
      r_402__17_ <= r_n_402__17_;
      r_402__16_ <= r_n_402__16_;
      r_402__15_ <= r_n_402__15_;
      r_402__14_ <= r_n_402__14_;
      r_402__13_ <= r_n_402__13_;
      r_402__12_ <= r_n_402__12_;
      r_402__11_ <= r_n_402__11_;
      r_402__10_ <= r_n_402__10_;
      r_402__9_ <= r_n_402__9_;
      r_402__8_ <= r_n_402__8_;
      r_402__7_ <= r_n_402__7_;
      r_402__6_ <= r_n_402__6_;
      r_402__5_ <= r_n_402__5_;
      r_402__4_ <= r_n_402__4_;
      r_402__3_ <= r_n_402__3_;
      r_402__2_ <= r_n_402__2_;
      r_402__1_ <= r_n_402__1_;
      r_402__0_ <= r_n_402__0_;
    end 
    if(N3987) begin
      r_403__63_ <= r_n_403__63_;
      r_403__62_ <= r_n_403__62_;
      r_403__61_ <= r_n_403__61_;
      r_403__60_ <= r_n_403__60_;
      r_403__59_ <= r_n_403__59_;
      r_403__58_ <= r_n_403__58_;
      r_403__57_ <= r_n_403__57_;
      r_403__56_ <= r_n_403__56_;
      r_403__55_ <= r_n_403__55_;
      r_403__54_ <= r_n_403__54_;
      r_403__53_ <= r_n_403__53_;
      r_403__52_ <= r_n_403__52_;
      r_403__51_ <= r_n_403__51_;
      r_403__50_ <= r_n_403__50_;
      r_403__49_ <= r_n_403__49_;
      r_403__48_ <= r_n_403__48_;
      r_403__47_ <= r_n_403__47_;
      r_403__46_ <= r_n_403__46_;
      r_403__45_ <= r_n_403__45_;
      r_403__44_ <= r_n_403__44_;
      r_403__43_ <= r_n_403__43_;
      r_403__42_ <= r_n_403__42_;
      r_403__41_ <= r_n_403__41_;
      r_403__40_ <= r_n_403__40_;
      r_403__39_ <= r_n_403__39_;
      r_403__38_ <= r_n_403__38_;
      r_403__37_ <= r_n_403__37_;
      r_403__36_ <= r_n_403__36_;
      r_403__35_ <= r_n_403__35_;
      r_403__34_ <= r_n_403__34_;
      r_403__33_ <= r_n_403__33_;
      r_403__32_ <= r_n_403__32_;
      r_403__31_ <= r_n_403__31_;
      r_403__30_ <= r_n_403__30_;
      r_403__29_ <= r_n_403__29_;
      r_403__28_ <= r_n_403__28_;
      r_403__27_ <= r_n_403__27_;
      r_403__26_ <= r_n_403__26_;
      r_403__25_ <= r_n_403__25_;
      r_403__24_ <= r_n_403__24_;
      r_403__23_ <= r_n_403__23_;
      r_403__22_ <= r_n_403__22_;
      r_403__21_ <= r_n_403__21_;
      r_403__20_ <= r_n_403__20_;
      r_403__19_ <= r_n_403__19_;
      r_403__18_ <= r_n_403__18_;
      r_403__17_ <= r_n_403__17_;
      r_403__16_ <= r_n_403__16_;
      r_403__15_ <= r_n_403__15_;
      r_403__14_ <= r_n_403__14_;
      r_403__13_ <= r_n_403__13_;
      r_403__12_ <= r_n_403__12_;
      r_403__11_ <= r_n_403__11_;
      r_403__10_ <= r_n_403__10_;
      r_403__9_ <= r_n_403__9_;
      r_403__8_ <= r_n_403__8_;
      r_403__7_ <= r_n_403__7_;
      r_403__6_ <= r_n_403__6_;
      r_403__5_ <= r_n_403__5_;
      r_403__4_ <= r_n_403__4_;
      r_403__3_ <= r_n_403__3_;
      r_403__2_ <= r_n_403__2_;
      r_403__1_ <= r_n_403__1_;
      r_403__0_ <= r_n_403__0_;
    end 
    if(N3988) begin
      r_404__63_ <= r_n_404__63_;
      r_404__62_ <= r_n_404__62_;
      r_404__61_ <= r_n_404__61_;
      r_404__60_ <= r_n_404__60_;
      r_404__59_ <= r_n_404__59_;
      r_404__58_ <= r_n_404__58_;
      r_404__57_ <= r_n_404__57_;
      r_404__56_ <= r_n_404__56_;
      r_404__55_ <= r_n_404__55_;
      r_404__54_ <= r_n_404__54_;
      r_404__53_ <= r_n_404__53_;
      r_404__52_ <= r_n_404__52_;
      r_404__51_ <= r_n_404__51_;
      r_404__50_ <= r_n_404__50_;
      r_404__49_ <= r_n_404__49_;
      r_404__48_ <= r_n_404__48_;
      r_404__47_ <= r_n_404__47_;
      r_404__46_ <= r_n_404__46_;
      r_404__45_ <= r_n_404__45_;
      r_404__44_ <= r_n_404__44_;
      r_404__43_ <= r_n_404__43_;
      r_404__42_ <= r_n_404__42_;
      r_404__41_ <= r_n_404__41_;
      r_404__40_ <= r_n_404__40_;
      r_404__39_ <= r_n_404__39_;
      r_404__38_ <= r_n_404__38_;
      r_404__37_ <= r_n_404__37_;
      r_404__36_ <= r_n_404__36_;
      r_404__35_ <= r_n_404__35_;
      r_404__34_ <= r_n_404__34_;
      r_404__33_ <= r_n_404__33_;
      r_404__32_ <= r_n_404__32_;
      r_404__31_ <= r_n_404__31_;
      r_404__30_ <= r_n_404__30_;
      r_404__29_ <= r_n_404__29_;
      r_404__28_ <= r_n_404__28_;
      r_404__27_ <= r_n_404__27_;
      r_404__26_ <= r_n_404__26_;
      r_404__25_ <= r_n_404__25_;
      r_404__24_ <= r_n_404__24_;
      r_404__23_ <= r_n_404__23_;
      r_404__22_ <= r_n_404__22_;
      r_404__21_ <= r_n_404__21_;
      r_404__20_ <= r_n_404__20_;
      r_404__19_ <= r_n_404__19_;
      r_404__18_ <= r_n_404__18_;
      r_404__17_ <= r_n_404__17_;
      r_404__16_ <= r_n_404__16_;
      r_404__15_ <= r_n_404__15_;
      r_404__14_ <= r_n_404__14_;
      r_404__13_ <= r_n_404__13_;
      r_404__12_ <= r_n_404__12_;
      r_404__11_ <= r_n_404__11_;
      r_404__10_ <= r_n_404__10_;
      r_404__9_ <= r_n_404__9_;
      r_404__8_ <= r_n_404__8_;
      r_404__7_ <= r_n_404__7_;
      r_404__6_ <= r_n_404__6_;
      r_404__5_ <= r_n_404__5_;
      r_404__4_ <= r_n_404__4_;
      r_404__3_ <= r_n_404__3_;
      r_404__2_ <= r_n_404__2_;
      r_404__1_ <= r_n_404__1_;
      r_404__0_ <= r_n_404__0_;
    end 
    if(N3989) begin
      r_405__63_ <= r_n_405__63_;
      r_405__62_ <= r_n_405__62_;
      r_405__61_ <= r_n_405__61_;
      r_405__60_ <= r_n_405__60_;
      r_405__59_ <= r_n_405__59_;
      r_405__58_ <= r_n_405__58_;
      r_405__57_ <= r_n_405__57_;
      r_405__56_ <= r_n_405__56_;
      r_405__55_ <= r_n_405__55_;
      r_405__54_ <= r_n_405__54_;
      r_405__53_ <= r_n_405__53_;
      r_405__52_ <= r_n_405__52_;
      r_405__51_ <= r_n_405__51_;
      r_405__50_ <= r_n_405__50_;
      r_405__49_ <= r_n_405__49_;
      r_405__48_ <= r_n_405__48_;
      r_405__47_ <= r_n_405__47_;
      r_405__46_ <= r_n_405__46_;
      r_405__45_ <= r_n_405__45_;
      r_405__44_ <= r_n_405__44_;
      r_405__43_ <= r_n_405__43_;
      r_405__42_ <= r_n_405__42_;
      r_405__41_ <= r_n_405__41_;
      r_405__40_ <= r_n_405__40_;
      r_405__39_ <= r_n_405__39_;
      r_405__38_ <= r_n_405__38_;
      r_405__37_ <= r_n_405__37_;
      r_405__36_ <= r_n_405__36_;
      r_405__35_ <= r_n_405__35_;
      r_405__34_ <= r_n_405__34_;
      r_405__33_ <= r_n_405__33_;
      r_405__32_ <= r_n_405__32_;
      r_405__31_ <= r_n_405__31_;
      r_405__30_ <= r_n_405__30_;
      r_405__29_ <= r_n_405__29_;
      r_405__28_ <= r_n_405__28_;
      r_405__27_ <= r_n_405__27_;
      r_405__26_ <= r_n_405__26_;
      r_405__25_ <= r_n_405__25_;
      r_405__24_ <= r_n_405__24_;
      r_405__23_ <= r_n_405__23_;
      r_405__22_ <= r_n_405__22_;
      r_405__21_ <= r_n_405__21_;
      r_405__20_ <= r_n_405__20_;
      r_405__19_ <= r_n_405__19_;
      r_405__18_ <= r_n_405__18_;
      r_405__17_ <= r_n_405__17_;
      r_405__16_ <= r_n_405__16_;
      r_405__15_ <= r_n_405__15_;
      r_405__14_ <= r_n_405__14_;
      r_405__13_ <= r_n_405__13_;
      r_405__12_ <= r_n_405__12_;
      r_405__11_ <= r_n_405__11_;
      r_405__10_ <= r_n_405__10_;
      r_405__9_ <= r_n_405__9_;
      r_405__8_ <= r_n_405__8_;
      r_405__7_ <= r_n_405__7_;
      r_405__6_ <= r_n_405__6_;
      r_405__5_ <= r_n_405__5_;
      r_405__4_ <= r_n_405__4_;
      r_405__3_ <= r_n_405__3_;
      r_405__2_ <= r_n_405__2_;
      r_405__1_ <= r_n_405__1_;
      r_405__0_ <= r_n_405__0_;
    end 
    if(N3990) begin
      r_406__63_ <= r_n_406__63_;
      r_406__62_ <= r_n_406__62_;
      r_406__61_ <= r_n_406__61_;
      r_406__60_ <= r_n_406__60_;
      r_406__59_ <= r_n_406__59_;
      r_406__58_ <= r_n_406__58_;
      r_406__57_ <= r_n_406__57_;
      r_406__56_ <= r_n_406__56_;
      r_406__55_ <= r_n_406__55_;
      r_406__54_ <= r_n_406__54_;
      r_406__53_ <= r_n_406__53_;
      r_406__52_ <= r_n_406__52_;
      r_406__51_ <= r_n_406__51_;
      r_406__50_ <= r_n_406__50_;
      r_406__49_ <= r_n_406__49_;
      r_406__48_ <= r_n_406__48_;
      r_406__47_ <= r_n_406__47_;
      r_406__46_ <= r_n_406__46_;
      r_406__45_ <= r_n_406__45_;
      r_406__44_ <= r_n_406__44_;
      r_406__43_ <= r_n_406__43_;
      r_406__42_ <= r_n_406__42_;
      r_406__41_ <= r_n_406__41_;
      r_406__40_ <= r_n_406__40_;
      r_406__39_ <= r_n_406__39_;
      r_406__38_ <= r_n_406__38_;
      r_406__37_ <= r_n_406__37_;
      r_406__36_ <= r_n_406__36_;
      r_406__35_ <= r_n_406__35_;
      r_406__34_ <= r_n_406__34_;
      r_406__33_ <= r_n_406__33_;
      r_406__32_ <= r_n_406__32_;
      r_406__31_ <= r_n_406__31_;
      r_406__30_ <= r_n_406__30_;
      r_406__29_ <= r_n_406__29_;
      r_406__28_ <= r_n_406__28_;
      r_406__27_ <= r_n_406__27_;
      r_406__26_ <= r_n_406__26_;
      r_406__25_ <= r_n_406__25_;
      r_406__24_ <= r_n_406__24_;
      r_406__23_ <= r_n_406__23_;
      r_406__22_ <= r_n_406__22_;
      r_406__21_ <= r_n_406__21_;
      r_406__20_ <= r_n_406__20_;
      r_406__19_ <= r_n_406__19_;
      r_406__18_ <= r_n_406__18_;
      r_406__17_ <= r_n_406__17_;
      r_406__16_ <= r_n_406__16_;
      r_406__15_ <= r_n_406__15_;
      r_406__14_ <= r_n_406__14_;
      r_406__13_ <= r_n_406__13_;
      r_406__12_ <= r_n_406__12_;
      r_406__11_ <= r_n_406__11_;
      r_406__10_ <= r_n_406__10_;
      r_406__9_ <= r_n_406__9_;
      r_406__8_ <= r_n_406__8_;
      r_406__7_ <= r_n_406__7_;
      r_406__6_ <= r_n_406__6_;
      r_406__5_ <= r_n_406__5_;
      r_406__4_ <= r_n_406__4_;
      r_406__3_ <= r_n_406__3_;
      r_406__2_ <= r_n_406__2_;
      r_406__1_ <= r_n_406__1_;
      r_406__0_ <= r_n_406__0_;
    end 
    if(N3991) begin
      r_407__63_ <= r_n_407__63_;
      r_407__62_ <= r_n_407__62_;
      r_407__61_ <= r_n_407__61_;
      r_407__60_ <= r_n_407__60_;
      r_407__59_ <= r_n_407__59_;
      r_407__58_ <= r_n_407__58_;
      r_407__57_ <= r_n_407__57_;
      r_407__56_ <= r_n_407__56_;
      r_407__55_ <= r_n_407__55_;
      r_407__54_ <= r_n_407__54_;
      r_407__53_ <= r_n_407__53_;
      r_407__52_ <= r_n_407__52_;
      r_407__51_ <= r_n_407__51_;
      r_407__50_ <= r_n_407__50_;
      r_407__49_ <= r_n_407__49_;
      r_407__48_ <= r_n_407__48_;
      r_407__47_ <= r_n_407__47_;
      r_407__46_ <= r_n_407__46_;
      r_407__45_ <= r_n_407__45_;
      r_407__44_ <= r_n_407__44_;
      r_407__43_ <= r_n_407__43_;
      r_407__42_ <= r_n_407__42_;
      r_407__41_ <= r_n_407__41_;
      r_407__40_ <= r_n_407__40_;
      r_407__39_ <= r_n_407__39_;
      r_407__38_ <= r_n_407__38_;
      r_407__37_ <= r_n_407__37_;
      r_407__36_ <= r_n_407__36_;
      r_407__35_ <= r_n_407__35_;
      r_407__34_ <= r_n_407__34_;
      r_407__33_ <= r_n_407__33_;
      r_407__32_ <= r_n_407__32_;
      r_407__31_ <= r_n_407__31_;
      r_407__30_ <= r_n_407__30_;
      r_407__29_ <= r_n_407__29_;
      r_407__28_ <= r_n_407__28_;
      r_407__27_ <= r_n_407__27_;
      r_407__26_ <= r_n_407__26_;
      r_407__25_ <= r_n_407__25_;
      r_407__24_ <= r_n_407__24_;
      r_407__23_ <= r_n_407__23_;
      r_407__22_ <= r_n_407__22_;
      r_407__21_ <= r_n_407__21_;
      r_407__20_ <= r_n_407__20_;
      r_407__19_ <= r_n_407__19_;
      r_407__18_ <= r_n_407__18_;
      r_407__17_ <= r_n_407__17_;
      r_407__16_ <= r_n_407__16_;
      r_407__15_ <= r_n_407__15_;
      r_407__14_ <= r_n_407__14_;
      r_407__13_ <= r_n_407__13_;
      r_407__12_ <= r_n_407__12_;
      r_407__11_ <= r_n_407__11_;
      r_407__10_ <= r_n_407__10_;
      r_407__9_ <= r_n_407__9_;
      r_407__8_ <= r_n_407__8_;
      r_407__7_ <= r_n_407__7_;
      r_407__6_ <= r_n_407__6_;
      r_407__5_ <= r_n_407__5_;
      r_407__4_ <= r_n_407__4_;
      r_407__3_ <= r_n_407__3_;
      r_407__2_ <= r_n_407__2_;
      r_407__1_ <= r_n_407__1_;
      r_407__0_ <= r_n_407__0_;
    end 
    if(N3992) begin
      r_408__63_ <= r_n_408__63_;
      r_408__62_ <= r_n_408__62_;
      r_408__61_ <= r_n_408__61_;
      r_408__60_ <= r_n_408__60_;
      r_408__59_ <= r_n_408__59_;
      r_408__58_ <= r_n_408__58_;
      r_408__57_ <= r_n_408__57_;
      r_408__56_ <= r_n_408__56_;
      r_408__55_ <= r_n_408__55_;
      r_408__54_ <= r_n_408__54_;
      r_408__53_ <= r_n_408__53_;
      r_408__52_ <= r_n_408__52_;
      r_408__51_ <= r_n_408__51_;
      r_408__50_ <= r_n_408__50_;
      r_408__49_ <= r_n_408__49_;
      r_408__48_ <= r_n_408__48_;
      r_408__47_ <= r_n_408__47_;
      r_408__46_ <= r_n_408__46_;
      r_408__45_ <= r_n_408__45_;
      r_408__44_ <= r_n_408__44_;
      r_408__43_ <= r_n_408__43_;
      r_408__42_ <= r_n_408__42_;
      r_408__41_ <= r_n_408__41_;
      r_408__40_ <= r_n_408__40_;
      r_408__39_ <= r_n_408__39_;
      r_408__38_ <= r_n_408__38_;
      r_408__37_ <= r_n_408__37_;
      r_408__36_ <= r_n_408__36_;
      r_408__35_ <= r_n_408__35_;
      r_408__34_ <= r_n_408__34_;
      r_408__33_ <= r_n_408__33_;
      r_408__32_ <= r_n_408__32_;
      r_408__31_ <= r_n_408__31_;
      r_408__30_ <= r_n_408__30_;
      r_408__29_ <= r_n_408__29_;
      r_408__28_ <= r_n_408__28_;
      r_408__27_ <= r_n_408__27_;
      r_408__26_ <= r_n_408__26_;
      r_408__25_ <= r_n_408__25_;
      r_408__24_ <= r_n_408__24_;
      r_408__23_ <= r_n_408__23_;
      r_408__22_ <= r_n_408__22_;
      r_408__21_ <= r_n_408__21_;
      r_408__20_ <= r_n_408__20_;
      r_408__19_ <= r_n_408__19_;
      r_408__18_ <= r_n_408__18_;
      r_408__17_ <= r_n_408__17_;
      r_408__16_ <= r_n_408__16_;
      r_408__15_ <= r_n_408__15_;
      r_408__14_ <= r_n_408__14_;
      r_408__13_ <= r_n_408__13_;
      r_408__12_ <= r_n_408__12_;
      r_408__11_ <= r_n_408__11_;
      r_408__10_ <= r_n_408__10_;
      r_408__9_ <= r_n_408__9_;
      r_408__8_ <= r_n_408__8_;
      r_408__7_ <= r_n_408__7_;
      r_408__6_ <= r_n_408__6_;
      r_408__5_ <= r_n_408__5_;
      r_408__4_ <= r_n_408__4_;
      r_408__3_ <= r_n_408__3_;
      r_408__2_ <= r_n_408__2_;
      r_408__1_ <= r_n_408__1_;
      r_408__0_ <= r_n_408__0_;
    end 
    if(N3993) begin
      r_409__63_ <= r_n_409__63_;
      r_409__62_ <= r_n_409__62_;
      r_409__61_ <= r_n_409__61_;
      r_409__60_ <= r_n_409__60_;
      r_409__59_ <= r_n_409__59_;
      r_409__58_ <= r_n_409__58_;
      r_409__57_ <= r_n_409__57_;
      r_409__56_ <= r_n_409__56_;
      r_409__55_ <= r_n_409__55_;
      r_409__54_ <= r_n_409__54_;
      r_409__53_ <= r_n_409__53_;
      r_409__52_ <= r_n_409__52_;
      r_409__51_ <= r_n_409__51_;
      r_409__50_ <= r_n_409__50_;
      r_409__49_ <= r_n_409__49_;
      r_409__48_ <= r_n_409__48_;
      r_409__47_ <= r_n_409__47_;
      r_409__46_ <= r_n_409__46_;
      r_409__45_ <= r_n_409__45_;
      r_409__44_ <= r_n_409__44_;
      r_409__43_ <= r_n_409__43_;
      r_409__42_ <= r_n_409__42_;
      r_409__41_ <= r_n_409__41_;
      r_409__40_ <= r_n_409__40_;
      r_409__39_ <= r_n_409__39_;
      r_409__38_ <= r_n_409__38_;
      r_409__37_ <= r_n_409__37_;
      r_409__36_ <= r_n_409__36_;
      r_409__35_ <= r_n_409__35_;
      r_409__34_ <= r_n_409__34_;
      r_409__33_ <= r_n_409__33_;
      r_409__32_ <= r_n_409__32_;
      r_409__31_ <= r_n_409__31_;
      r_409__30_ <= r_n_409__30_;
      r_409__29_ <= r_n_409__29_;
      r_409__28_ <= r_n_409__28_;
      r_409__27_ <= r_n_409__27_;
      r_409__26_ <= r_n_409__26_;
      r_409__25_ <= r_n_409__25_;
      r_409__24_ <= r_n_409__24_;
      r_409__23_ <= r_n_409__23_;
      r_409__22_ <= r_n_409__22_;
      r_409__21_ <= r_n_409__21_;
      r_409__20_ <= r_n_409__20_;
      r_409__19_ <= r_n_409__19_;
      r_409__18_ <= r_n_409__18_;
      r_409__17_ <= r_n_409__17_;
      r_409__16_ <= r_n_409__16_;
      r_409__15_ <= r_n_409__15_;
      r_409__14_ <= r_n_409__14_;
      r_409__13_ <= r_n_409__13_;
      r_409__12_ <= r_n_409__12_;
      r_409__11_ <= r_n_409__11_;
      r_409__10_ <= r_n_409__10_;
      r_409__9_ <= r_n_409__9_;
      r_409__8_ <= r_n_409__8_;
      r_409__7_ <= r_n_409__7_;
      r_409__6_ <= r_n_409__6_;
      r_409__5_ <= r_n_409__5_;
      r_409__4_ <= r_n_409__4_;
      r_409__3_ <= r_n_409__3_;
      r_409__2_ <= r_n_409__2_;
      r_409__1_ <= r_n_409__1_;
      r_409__0_ <= r_n_409__0_;
    end 
    if(N3994) begin
      r_410__63_ <= r_n_410__63_;
      r_410__62_ <= r_n_410__62_;
      r_410__61_ <= r_n_410__61_;
      r_410__60_ <= r_n_410__60_;
      r_410__59_ <= r_n_410__59_;
      r_410__58_ <= r_n_410__58_;
      r_410__57_ <= r_n_410__57_;
      r_410__56_ <= r_n_410__56_;
      r_410__55_ <= r_n_410__55_;
      r_410__54_ <= r_n_410__54_;
      r_410__53_ <= r_n_410__53_;
      r_410__52_ <= r_n_410__52_;
      r_410__51_ <= r_n_410__51_;
      r_410__50_ <= r_n_410__50_;
      r_410__49_ <= r_n_410__49_;
      r_410__48_ <= r_n_410__48_;
      r_410__47_ <= r_n_410__47_;
      r_410__46_ <= r_n_410__46_;
      r_410__45_ <= r_n_410__45_;
      r_410__44_ <= r_n_410__44_;
      r_410__43_ <= r_n_410__43_;
      r_410__42_ <= r_n_410__42_;
      r_410__41_ <= r_n_410__41_;
      r_410__40_ <= r_n_410__40_;
      r_410__39_ <= r_n_410__39_;
      r_410__38_ <= r_n_410__38_;
      r_410__37_ <= r_n_410__37_;
      r_410__36_ <= r_n_410__36_;
      r_410__35_ <= r_n_410__35_;
      r_410__34_ <= r_n_410__34_;
      r_410__33_ <= r_n_410__33_;
      r_410__32_ <= r_n_410__32_;
      r_410__31_ <= r_n_410__31_;
      r_410__30_ <= r_n_410__30_;
      r_410__29_ <= r_n_410__29_;
      r_410__28_ <= r_n_410__28_;
      r_410__27_ <= r_n_410__27_;
      r_410__26_ <= r_n_410__26_;
      r_410__25_ <= r_n_410__25_;
      r_410__24_ <= r_n_410__24_;
      r_410__23_ <= r_n_410__23_;
      r_410__22_ <= r_n_410__22_;
      r_410__21_ <= r_n_410__21_;
      r_410__20_ <= r_n_410__20_;
      r_410__19_ <= r_n_410__19_;
      r_410__18_ <= r_n_410__18_;
      r_410__17_ <= r_n_410__17_;
      r_410__16_ <= r_n_410__16_;
      r_410__15_ <= r_n_410__15_;
      r_410__14_ <= r_n_410__14_;
      r_410__13_ <= r_n_410__13_;
      r_410__12_ <= r_n_410__12_;
      r_410__11_ <= r_n_410__11_;
      r_410__10_ <= r_n_410__10_;
      r_410__9_ <= r_n_410__9_;
      r_410__8_ <= r_n_410__8_;
      r_410__7_ <= r_n_410__7_;
      r_410__6_ <= r_n_410__6_;
      r_410__5_ <= r_n_410__5_;
      r_410__4_ <= r_n_410__4_;
      r_410__3_ <= r_n_410__3_;
      r_410__2_ <= r_n_410__2_;
      r_410__1_ <= r_n_410__1_;
      r_410__0_ <= r_n_410__0_;
    end 
    if(N3995) begin
      r_411__63_ <= r_n_411__63_;
      r_411__62_ <= r_n_411__62_;
      r_411__61_ <= r_n_411__61_;
      r_411__60_ <= r_n_411__60_;
      r_411__59_ <= r_n_411__59_;
      r_411__58_ <= r_n_411__58_;
      r_411__57_ <= r_n_411__57_;
      r_411__56_ <= r_n_411__56_;
      r_411__55_ <= r_n_411__55_;
      r_411__54_ <= r_n_411__54_;
      r_411__53_ <= r_n_411__53_;
      r_411__52_ <= r_n_411__52_;
      r_411__51_ <= r_n_411__51_;
      r_411__50_ <= r_n_411__50_;
      r_411__49_ <= r_n_411__49_;
      r_411__48_ <= r_n_411__48_;
      r_411__47_ <= r_n_411__47_;
      r_411__46_ <= r_n_411__46_;
      r_411__45_ <= r_n_411__45_;
      r_411__44_ <= r_n_411__44_;
      r_411__43_ <= r_n_411__43_;
      r_411__42_ <= r_n_411__42_;
      r_411__41_ <= r_n_411__41_;
      r_411__40_ <= r_n_411__40_;
      r_411__39_ <= r_n_411__39_;
      r_411__38_ <= r_n_411__38_;
      r_411__37_ <= r_n_411__37_;
      r_411__36_ <= r_n_411__36_;
      r_411__35_ <= r_n_411__35_;
      r_411__34_ <= r_n_411__34_;
      r_411__33_ <= r_n_411__33_;
      r_411__32_ <= r_n_411__32_;
      r_411__31_ <= r_n_411__31_;
      r_411__30_ <= r_n_411__30_;
      r_411__29_ <= r_n_411__29_;
      r_411__28_ <= r_n_411__28_;
      r_411__27_ <= r_n_411__27_;
      r_411__26_ <= r_n_411__26_;
      r_411__25_ <= r_n_411__25_;
      r_411__24_ <= r_n_411__24_;
      r_411__23_ <= r_n_411__23_;
      r_411__22_ <= r_n_411__22_;
      r_411__21_ <= r_n_411__21_;
      r_411__20_ <= r_n_411__20_;
      r_411__19_ <= r_n_411__19_;
      r_411__18_ <= r_n_411__18_;
      r_411__17_ <= r_n_411__17_;
      r_411__16_ <= r_n_411__16_;
      r_411__15_ <= r_n_411__15_;
      r_411__14_ <= r_n_411__14_;
      r_411__13_ <= r_n_411__13_;
      r_411__12_ <= r_n_411__12_;
      r_411__11_ <= r_n_411__11_;
      r_411__10_ <= r_n_411__10_;
      r_411__9_ <= r_n_411__9_;
      r_411__8_ <= r_n_411__8_;
      r_411__7_ <= r_n_411__7_;
      r_411__6_ <= r_n_411__6_;
      r_411__5_ <= r_n_411__5_;
      r_411__4_ <= r_n_411__4_;
      r_411__3_ <= r_n_411__3_;
      r_411__2_ <= r_n_411__2_;
      r_411__1_ <= r_n_411__1_;
      r_411__0_ <= r_n_411__0_;
    end 
    if(N3996) begin
      r_412__63_ <= r_n_412__63_;
      r_412__62_ <= r_n_412__62_;
      r_412__61_ <= r_n_412__61_;
      r_412__60_ <= r_n_412__60_;
      r_412__59_ <= r_n_412__59_;
      r_412__58_ <= r_n_412__58_;
      r_412__57_ <= r_n_412__57_;
      r_412__56_ <= r_n_412__56_;
      r_412__55_ <= r_n_412__55_;
      r_412__54_ <= r_n_412__54_;
      r_412__53_ <= r_n_412__53_;
      r_412__52_ <= r_n_412__52_;
      r_412__51_ <= r_n_412__51_;
      r_412__50_ <= r_n_412__50_;
      r_412__49_ <= r_n_412__49_;
      r_412__48_ <= r_n_412__48_;
      r_412__47_ <= r_n_412__47_;
      r_412__46_ <= r_n_412__46_;
      r_412__45_ <= r_n_412__45_;
      r_412__44_ <= r_n_412__44_;
      r_412__43_ <= r_n_412__43_;
      r_412__42_ <= r_n_412__42_;
      r_412__41_ <= r_n_412__41_;
      r_412__40_ <= r_n_412__40_;
      r_412__39_ <= r_n_412__39_;
      r_412__38_ <= r_n_412__38_;
      r_412__37_ <= r_n_412__37_;
      r_412__36_ <= r_n_412__36_;
      r_412__35_ <= r_n_412__35_;
      r_412__34_ <= r_n_412__34_;
      r_412__33_ <= r_n_412__33_;
      r_412__32_ <= r_n_412__32_;
      r_412__31_ <= r_n_412__31_;
      r_412__30_ <= r_n_412__30_;
      r_412__29_ <= r_n_412__29_;
      r_412__28_ <= r_n_412__28_;
      r_412__27_ <= r_n_412__27_;
      r_412__26_ <= r_n_412__26_;
      r_412__25_ <= r_n_412__25_;
      r_412__24_ <= r_n_412__24_;
      r_412__23_ <= r_n_412__23_;
      r_412__22_ <= r_n_412__22_;
      r_412__21_ <= r_n_412__21_;
      r_412__20_ <= r_n_412__20_;
      r_412__19_ <= r_n_412__19_;
      r_412__18_ <= r_n_412__18_;
      r_412__17_ <= r_n_412__17_;
      r_412__16_ <= r_n_412__16_;
      r_412__15_ <= r_n_412__15_;
      r_412__14_ <= r_n_412__14_;
      r_412__13_ <= r_n_412__13_;
      r_412__12_ <= r_n_412__12_;
      r_412__11_ <= r_n_412__11_;
      r_412__10_ <= r_n_412__10_;
      r_412__9_ <= r_n_412__9_;
      r_412__8_ <= r_n_412__8_;
      r_412__7_ <= r_n_412__7_;
      r_412__6_ <= r_n_412__6_;
      r_412__5_ <= r_n_412__5_;
      r_412__4_ <= r_n_412__4_;
      r_412__3_ <= r_n_412__3_;
      r_412__2_ <= r_n_412__2_;
      r_412__1_ <= r_n_412__1_;
      r_412__0_ <= r_n_412__0_;
    end 
    if(N3997) begin
      r_413__63_ <= r_n_413__63_;
      r_413__62_ <= r_n_413__62_;
      r_413__61_ <= r_n_413__61_;
      r_413__60_ <= r_n_413__60_;
      r_413__59_ <= r_n_413__59_;
      r_413__58_ <= r_n_413__58_;
      r_413__57_ <= r_n_413__57_;
      r_413__56_ <= r_n_413__56_;
      r_413__55_ <= r_n_413__55_;
      r_413__54_ <= r_n_413__54_;
      r_413__53_ <= r_n_413__53_;
      r_413__52_ <= r_n_413__52_;
      r_413__51_ <= r_n_413__51_;
      r_413__50_ <= r_n_413__50_;
      r_413__49_ <= r_n_413__49_;
      r_413__48_ <= r_n_413__48_;
      r_413__47_ <= r_n_413__47_;
      r_413__46_ <= r_n_413__46_;
      r_413__45_ <= r_n_413__45_;
      r_413__44_ <= r_n_413__44_;
      r_413__43_ <= r_n_413__43_;
      r_413__42_ <= r_n_413__42_;
      r_413__41_ <= r_n_413__41_;
      r_413__40_ <= r_n_413__40_;
      r_413__39_ <= r_n_413__39_;
      r_413__38_ <= r_n_413__38_;
      r_413__37_ <= r_n_413__37_;
      r_413__36_ <= r_n_413__36_;
      r_413__35_ <= r_n_413__35_;
      r_413__34_ <= r_n_413__34_;
      r_413__33_ <= r_n_413__33_;
      r_413__32_ <= r_n_413__32_;
      r_413__31_ <= r_n_413__31_;
      r_413__30_ <= r_n_413__30_;
      r_413__29_ <= r_n_413__29_;
      r_413__28_ <= r_n_413__28_;
      r_413__27_ <= r_n_413__27_;
      r_413__26_ <= r_n_413__26_;
      r_413__25_ <= r_n_413__25_;
      r_413__24_ <= r_n_413__24_;
      r_413__23_ <= r_n_413__23_;
      r_413__22_ <= r_n_413__22_;
      r_413__21_ <= r_n_413__21_;
      r_413__20_ <= r_n_413__20_;
      r_413__19_ <= r_n_413__19_;
      r_413__18_ <= r_n_413__18_;
      r_413__17_ <= r_n_413__17_;
      r_413__16_ <= r_n_413__16_;
      r_413__15_ <= r_n_413__15_;
      r_413__14_ <= r_n_413__14_;
      r_413__13_ <= r_n_413__13_;
      r_413__12_ <= r_n_413__12_;
      r_413__11_ <= r_n_413__11_;
      r_413__10_ <= r_n_413__10_;
      r_413__9_ <= r_n_413__9_;
      r_413__8_ <= r_n_413__8_;
      r_413__7_ <= r_n_413__7_;
      r_413__6_ <= r_n_413__6_;
      r_413__5_ <= r_n_413__5_;
      r_413__4_ <= r_n_413__4_;
      r_413__3_ <= r_n_413__3_;
      r_413__2_ <= r_n_413__2_;
      r_413__1_ <= r_n_413__1_;
      r_413__0_ <= r_n_413__0_;
    end 
    if(N3998) begin
      r_414__63_ <= r_n_414__63_;
      r_414__62_ <= r_n_414__62_;
      r_414__61_ <= r_n_414__61_;
      r_414__60_ <= r_n_414__60_;
      r_414__59_ <= r_n_414__59_;
      r_414__58_ <= r_n_414__58_;
      r_414__57_ <= r_n_414__57_;
      r_414__56_ <= r_n_414__56_;
      r_414__55_ <= r_n_414__55_;
      r_414__54_ <= r_n_414__54_;
      r_414__53_ <= r_n_414__53_;
      r_414__52_ <= r_n_414__52_;
      r_414__51_ <= r_n_414__51_;
      r_414__50_ <= r_n_414__50_;
      r_414__49_ <= r_n_414__49_;
      r_414__48_ <= r_n_414__48_;
      r_414__47_ <= r_n_414__47_;
      r_414__46_ <= r_n_414__46_;
      r_414__45_ <= r_n_414__45_;
      r_414__44_ <= r_n_414__44_;
      r_414__43_ <= r_n_414__43_;
      r_414__42_ <= r_n_414__42_;
      r_414__41_ <= r_n_414__41_;
      r_414__40_ <= r_n_414__40_;
      r_414__39_ <= r_n_414__39_;
      r_414__38_ <= r_n_414__38_;
      r_414__37_ <= r_n_414__37_;
      r_414__36_ <= r_n_414__36_;
      r_414__35_ <= r_n_414__35_;
      r_414__34_ <= r_n_414__34_;
      r_414__33_ <= r_n_414__33_;
      r_414__32_ <= r_n_414__32_;
      r_414__31_ <= r_n_414__31_;
      r_414__30_ <= r_n_414__30_;
      r_414__29_ <= r_n_414__29_;
      r_414__28_ <= r_n_414__28_;
      r_414__27_ <= r_n_414__27_;
      r_414__26_ <= r_n_414__26_;
      r_414__25_ <= r_n_414__25_;
      r_414__24_ <= r_n_414__24_;
      r_414__23_ <= r_n_414__23_;
      r_414__22_ <= r_n_414__22_;
      r_414__21_ <= r_n_414__21_;
      r_414__20_ <= r_n_414__20_;
      r_414__19_ <= r_n_414__19_;
      r_414__18_ <= r_n_414__18_;
      r_414__17_ <= r_n_414__17_;
      r_414__16_ <= r_n_414__16_;
      r_414__15_ <= r_n_414__15_;
      r_414__14_ <= r_n_414__14_;
      r_414__13_ <= r_n_414__13_;
      r_414__12_ <= r_n_414__12_;
      r_414__11_ <= r_n_414__11_;
      r_414__10_ <= r_n_414__10_;
      r_414__9_ <= r_n_414__9_;
      r_414__8_ <= r_n_414__8_;
      r_414__7_ <= r_n_414__7_;
      r_414__6_ <= r_n_414__6_;
      r_414__5_ <= r_n_414__5_;
      r_414__4_ <= r_n_414__4_;
      r_414__3_ <= r_n_414__3_;
      r_414__2_ <= r_n_414__2_;
      r_414__1_ <= r_n_414__1_;
      r_414__0_ <= r_n_414__0_;
    end 
    if(N3999) begin
      r_415__63_ <= r_n_415__63_;
      r_415__62_ <= r_n_415__62_;
      r_415__61_ <= r_n_415__61_;
      r_415__60_ <= r_n_415__60_;
      r_415__59_ <= r_n_415__59_;
      r_415__58_ <= r_n_415__58_;
      r_415__57_ <= r_n_415__57_;
      r_415__56_ <= r_n_415__56_;
      r_415__55_ <= r_n_415__55_;
      r_415__54_ <= r_n_415__54_;
      r_415__53_ <= r_n_415__53_;
      r_415__52_ <= r_n_415__52_;
      r_415__51_ <= r_n_415__51_;
      r_415__50_ <= r_n_415__50_;
      r_415__49_ <= r_n_415__49_;
      r_415__48_ <= r_n_415__48_;
      r_415__47_ <= r_n_415__47_;
      r_415__46_ <= r_n_415__46_;
      r_415__45_ <= r_n_415__45_;
      r_415__44_ <= r_n_415__44_;
      r_415__43_ <= r_n_415__43_;
      r_415__42_ <= r_n_415__42_;
      r_415__41_ <= r_n_415__41_;
      r_415__40_ <= r_n_415__40_;
      r_415__39_ <= r_n_415__39_;
      r_415__38_ <= r_n_415__38_;
      r_415__37_ <= r_n_415__37_;
      r_415__36_ <= r_n_415__36_;
      r_415__35_ <= r_n_415__35_;
      r_415__34_ <= r_n_415__34_;
      r_415__33_ <= r_n_415__33_;
      r_415__32_ <= r_n_415__32_;
      r_415__31_ <= r_n_415__31_;
      r_415__30_ <= r_n_415__30_;
      r_415__29_ <= r_n_415__29_;
      r_415__28_ <= r_n_415__28_;
      r_415__27_ <= r_n_415__27_;
      r_415__26_ <= r_n_415__26_;
      r_415__25_ <= r_n_415__25_;
      r_415__24_ <= r_n_415__24_;
      r_415__23_ <= r_n_415__23_;
      r_415__22_ <= r_n_415__22_;
      r_415__21_ <= r_n_415__21_;
      r_415__20_ <= r_n_415__20_;
      r_415__19_ <= r_n_415__19_;
      r_415__18_ <= r_n_415__18_;
      r_415__17_ <= r_n_415__17_;
      r_415__16_ <= r_n_415__16_;
      r_415__15_ <= r_n_415__15_;
      r_415__14_ <= r_n_415__14_;
      r_415__13_ <= r_n_415__13_;
      r_415__12_ <= r_n_415__12_;
      r_415__11_ <= r_n_415__11_;
      r_415__10_ <= r_n_415__10_;
      r_415__9_ <= r_n_415__9_;
      r_415__8_ <= r_n_415__8_;
      r_415__7_ <= r_n_415__7_;
      r_415__6_ <= r_n_415__6_;
      r_415__5_ <= r_n_415__5_;
      r_415__4_ <= r_n_415__4_;
      r_415__3_ <= r_n_415__3_;
      r_415__2_ <= r_n_415__2_;
      r_415__1_ <= r_n_415__1_;
      r_415__0_ <= r_n_415__0_;
    end 
    if(N4000) begin
      r_416__63_ <= r_n_416__63_;
      r_416__62_ <= r_n_416__62_;
      r_416__61_ <= r_n_416__61_;
      r_416__60_ <= r_n_416__60_;
      r_416__59_ <= r_n_416__59_;
      r_416__58_ <= r_n_416__58_;
      r_416__57_ <= r_n_416__57_;
      r_416__56_ <= r_n_416__56_;
      r_416__55_ <= r_n_416__55_;
      r_416__54_ <= r_n_416__54_;
      r_416__53_ <= r_n_416__53_;
      r_416__52_ <= r_n_416__52_;
      r_416__51_ <= r_n_416__51_;
      r_416__50_ <= r_n_416__50_;
      r_416__49_ <= r_n_416__49_;
      r_416__48_ <= r_n_416__48_;
      r_416__47_ <= r_n_416__47_;
      r_416__46_ <= r_n_416__46_;
      r_416__45_ <= r_n_416__45_;
      r_416__44_ <= r_n_416__44_;
      r_416__43_ <= r_n_416__43_;
      r_416__42_ <= r_n_416__42_;
      r_416__41_ <= r_n_416__41_;
      r_416__40_ <= r_n_416__40_;
      r_416__39_ <= r_n_416__39_;
      r_416__38_ <= r_n_416__38_;
      r_416__37_ <= r_n_416__37_;
      r_416__36_ <= r_n_416__36_;
      r_416__35_ <= r_n_416__35_;
      r_416__34_ <= r_n_416__34_;
      r_416__33_ <= r_n_416__33_;
      r_416__32_ <= r_n_416__32_;
      r_416__31_ <= r_n_416__31_;
      r_416__30_ <= r_n_416__30_;
      r_416__29_ <= r_n_416__29_;
      r_416__28_ <= r_n_416__28_;
      r_416__27_ <= r_n_416__27_;
      r_416__26_ <= r_n_416__26_;
      r_416__25_ <= r_n_416__25_;
      r_416__24_ <= r_n_416__24_;
      r_416__23_ <= r_n_416__23_;
      r_416__22_ <= r_n_416__22_;
      r_416__21_ <= r_n_416__21_;
      r_416__20_ <= r_n_416__20_;
      r_416__19_ <= r_n_416__19_;
      r_416__18_ <= r_n_416__18_;
      r_416__17_ <= r_n_416__17_;
      r_416__16_ <= r_n_416__16_;
      r_416__15_ <= r_n_416__15_;
      r_416__14_ <= r_n_416__14_;
      r_416__13_ <= r_n_416__13_;
      r_416__12_ <= r_n_416__12_;
      r_416__11_ <= r_n_416__11_;
      r_416__10_ <= r_n_416__10_;
      r_416__9_ <= r_n_416__9_;
      r_416__8_ <= r_n_416__8_;
      r_416__7_ <= r_n_416__7_;
      r_416__6_ <= r_n_416__6_;
      r_416__5_ <= r_n_416__5_;
      r_416__4_ <= r_n_416__4_;
      r_416__3_ <= r_n_416__3_;
      r_416__2_ <= r_n_416__2_;
      r_416__1_ <= r_n_416__1_;
      r_416__0_ <= r_n_416__0_;
    end 
    if(N4001) begin
      r_417__63_ <= r_n_417__63_;
      r_417__62_ <= r_n_417__62_;
      r_417__61_ <= r_n_417__61_;
      r_417__60_ <= r_n_417__60_;
      r_417__59_ <= r_n_417__59_;
      r_417__58_ <= r_n_417__58_;
      r_417__57_ <= r_n_417__57_;
      r_417__56_ <= r_n_417__56_;
      r_417__55_ <= r_n_417__55_;
      r_417__54_ <= r_n_417__54_;
      r_417__53_ <= r_n_417__53_;
      r_417__52_ <= r_n_417__52_;
      r_417__51_ <= r_n_417__51_;
      r_417__50_ <= r_n_417__50_;
      r_417__49_ <= r_n_417__49_;
      r_417__48_ <= r_n_417__48_;
      r_417__47_ <= r_n_417__47_;
      r_417__46_ <= r_n_417__46_;
      r_417__45_ <= r_n_417__45_;
      r_417__44_ <= r_n_417__44_;
      r_417__43_ <= r_n_417__43_;
      r_417__42_ <= r_n_417__42_;
      r_417__41_ <= r_n_417__41_;
      r_417__40_ <= r_n_417__40_;
      r_417__39_ <= r_n_417__39_;
      r_417__38_ <= r_n_417__38_;
      r_417__37_ <= r_n_417__37_;
      r_417__36_ <= r_n_417__36_;
      r_417__35_ <= r_n_417__35_;
      r_417__34_ <= r_n_417__34_;
      r_417__33_ <= r_n_417__33_;
      r_417__32_ <= r_n_417__32_;
      r_417__31_ <= r_n_417__31_;
      r_417__30_ <= r_n_417__30_;
      r_417__29_ <= r_n_417__29_;
      r_417__28_ <= r_n_417__28_;
      r_417__27_ <= r_n_417__27_;
      r_417__26_ <= r_n_417__26_;
      r_417__25_ <= r_n_417__25_;
      r_417__24_ <= r_n_417__24_;
      r_417__23_ <= r_n_417__23_;
      r_417__22_ <= r_n_417__22_;
      r_417__21_ <= r_n_417__21_;
      r_417__20_ <= r_n_417__20_;
      r_417__19_ <= r_n_417__19_;
      r_417__18_ <= r_n_417__18_;
      r_417__17_ <= r_n_417__17_;
      r_417__16_ <= r_n_417__16_;
      r_417__15_ <= r_n_417__15_;
      r_417__14_ <= r_n_417__14_;
      r_417__13_ <= r_n_417__13_;
      r_417__12_ <= r_n_417__12_;
      r_417__11_ <= r_n_417__11_;
      r_417__10_ <= r_n_417__10_;
      r_417__9_ <= r_n_417__9_;
      r_417__8_ <= r_n_417__8_;
      r_417__7_ <= r_n_417__7_;
      r_417__6_ <= r_n_417__6_;
      r_417__5_ <= r_n_417__5_;
      r_417__4_ <= r_n_417__4_;
      r_417__3_ <= r_n_417__3_;
      r_417__2_ <= r_n_417__2_;
      r_417__1_ <= r_n_417__1_;
      r_417__0_ <= r_n_417__0_;
    end 
    if(N4002) begin
      r_418__63_ <= r_n_418__63_;
      r_418__62_ <= r_n_418__62_;
      r_418__61_ <= r_n_418__61_;
      r_418__60_ <= r_n_418__60_;
      r_418__59_ <= r_n_418__59_;
      r_418__58_ <= r_n_418__58_;
      r_418__57_ <= r_n_418__57_;
      r_418__56_ <= r_n_418__56_;
      r_418__55_ <= r_n_418__55_;
      r_418__54_ <= r_n_418__54_;
      r_418__53_ <= r_n_418__53_;
      r_418__52_ <= r_n_418__52_;
      r_418__51_ <= r_n_418__51_;
      r_418__50_ <= r_n_418__50_;
      r_418__49_ <= r_n_418__49_;
      r_418__48_ <= r_n_418__48_;
      r_418__47_ <= r_n_418__47_;
      r_418__46_ <= r_n_418__46_;
      r_418__45_ <= r_n_418__45_;
      r_418__44_ <= r_n_418__44_;
      r_418__43_ <= r_n_418__43_;
      r_418__42_ <= r_n_418__42_;
      r_418__41_ <= r_n_418__41_;
      r_418__40_ <= r_n_418__40_;
      r_418__39_ <= r_n_418__39_;
      r_418__38_ <= r_n_418__38_;
      r_418__37_ <= r_n_418__37_;
      r_418__36_ <= r_n_418__36_;
      r_418__35_ <= r_n_418__35_;
      r_418__34_ <= r_n_418__34_;
      r_418__33_ <= r_n_418__33_;
      r_418__32_ <= r_n_418__32_;
      r_418__31_ <= r_n_418__31_;
      r_418__30_ <= r_n_418__30_;
      r_418__29_ <= r_n_418__29_;
      r_418__28_ <= r_n_418__28_;
      r_418__27_ <= r_n_418__27_;
      r_418__26_ <= r_n_418__26_;
      r_418__25_ <= r_n_418__25_;
      r_418__24_ <= r_n_418__24_;
      r_418__23_ <= r_n_418__23_;
      r_418__22_ <= r_n_418__22_;
      r_418__21_ <= r_n_418__21_;
      r_418__20_ <= r_n_418__20_;
      r_418__19_ <= r_n_418__19_;
      r_418__18_ <= r_n_418__18_;
      r_418__17_ <= r_n_418__17_;
      r_418__16_ <= r_n_418__16_;
      r_418__15_ <= r_n_418__15_;
      r_418__14_ <= r_n_418__14_;
      r_418__13_ <= r_n_418__13_;
      r_418__12_ <= r_n_418__12_;
      r_418__11_ <= r_n_418__11_;
      r_418__10_ <= r_n_418__10_;
      r_418__9_ <= r_n_418__9_;
      r_418__8_ <= r_n_418__8_;
      r_418__7_ <= r_n_418__7_;
      r_418__6_ <= r_n_418__6_;
      r_418__5_ <= r_n_418__5_;
      r_418__4_ <= r_n_418__4_;
      r_418__3_ <= r_n_418__3_;
      r_418__2_ <= r_n_418__2_;
      r_418__1_ <= r_n_418__1_;
      r_418__0_ <= r_n_418__0_;
    end 
    if(N4003) begin
      r_419__63_ <= r_n_419__63_;
      r_419__62_ <= r_n_419__62_;
      r_419__61_ <= r_n_419__61_;
      r_419__60_ <= r_n_419__60_;
      r_419__59_ <= r_n_419__59_;
      r_419__58_ <= r_n_419__58_;
      r_419__57_ <= r_n_419__57_;
      r_419__56_ <= r_n_419__56_;
      r_419__55_ <= r_n_419__55_;
      r_419__54_ <= r_n_419__54_;
      r_419__53_ <= r_n_419__53_;
      r_419__52_ <= r_n_419__52_;
      r_419__51_ <= r_n_419__51_;
      r_419__50_ <= r_n_419__50_;
      r_419__49_ <= r_n_419__49_;
      r_419__48_ <= r_n_419__48_;
      r_419__47_ <= r_n_419__47_;
      r_419__46_ <= r_n_419__46_;
      r_419__45_ <= r_n_419__45_;
      r_419__44_ <= r_n_419__44_;
      r_419__43_ <= r_n_419__43_;
      r_419__42_ <= r_n_419__42_;
      r_419__41_ <= r_n_419__41_;
      r_419__40_ <= r_n_419__40_;
      r_419__39_ <= r_n_419__39_;
      r_419__38_ <= r_n_419__38_;
      r_419__37_ <= r_n_419__37_;
      r_419__36_ <= r_n_419__36_;
      r_419__35_ <= r_n_419__35_;
      r_419__34_ <= r_n_419__34_;
      r_419__33_ <= r_n_419__33_;
      r_419__32_ <= r_n_419__32_;
      r_419__31_ <= r_n_419__31_;
      r_419__30_ <= r_n_419__30_;
      r_419__29_ <= r_n_419__29_;
      r_419__28_ <= r_n_419__28_;
      r_419__27_ <= r_n_419__27_;
      r_419__26_ <= r_n_419__26_;
      r_419__25_ <= r_n_419__25_;
      r_419__24_ <= r_n_419__24_;
      r_419__23_ <= r_n_419__23_;
      r_419__22_ <= r_n_419__22_;
      r_419__21_ <= r_n_419__21_;
      r_419__20_ <= r_n_419__20_;
      r_419__19_ <= r_n_419__19_;
      r_419__18_ <= r_n_419__18_;
      r_419__17_ <= r_n_419__17_;
      r_419__16_ <= r_n_419__16_;
      r_419__15_ <= r_n_419__15_;
      r_419__14_ <= r_n_419__14_;
      r_419__13_ <= r_n_419__13_;
      r_419__12_ <= r_n_419__12_;
      r_419__11_ <= r_n_419__11_;
      r_419__10_ <= r_n_419__10_;
      r_419__9_ <= r_n_419__9_;
      r_419__8_ <= r_n_419__8_;
      r_419__7_ <= r_n_419__7_;
      r_419__6_ <= r_n_419__6_;
      r_419__5_ <= r_n_419__5_;
      r_419__4_ <= r_n_419__4_;
      r_419__3_ <= r_n_419__3_;
      r_419__2_ <= r_n_419__2_;
      r_419__1_ <= r_n_419__1_;
      r_419__0_ <= r_n_419__0_;
    end 
    if(N4004) begin
      r_420__63_ <= r_n_420__63_;
      r_420__62_ <= r_n_420__62_;
      r_420__61_ <= r_n_420__61_;
      r_420__60_ <= r_n_420__60_;
      r_420__59_ <= r_n_420__59_;
      r_420__58_ <= r_n_420__58_;
      r_420__57_ <= r_n_420__57_;
      r_420__56_ <= r_n_420__56_;
      r_420__55_ <= r_n_420__55_;
      r_420__54_ <= r_n_420__54_;
      r_420__53_ <= r_n_420__53_;
      r_420__52_ <= r_n_420__52_;
      r_420__51_ <= r_n_420__51_;
      r_420__50_ <= r_n_420__50_;
      r_420__49_ <= r_n_420__49_;
      r_420__48_ <= r_n_420__48_;
      r_420__47_ <= r_n_420__47_;
      r_420__46_ <= r_n_420__46_;
      r_420__45_ <= r_n_420__45_;
      r_420__44_ <= r_n_420__44_;
      r_420__43_ <= r_n_420__43_;
      r_420__42_ <= r_n_420__42_;
      r_420__41_ <= r_n_420__41_;
      r_420__40_ <= r_n_420__40_;
      r_420__39_ <= r_n_420__39_;
      r_420__38_ <= r_n_420__38_;
      r_420__37_ <= r_n_420__37_;
      r_420__36_ <= r_n_420__36_;
      r_420__35_ <= r_n_420__35_;
      r_420__34_ <= r_n_420__34_;
      r_420__33_ <= r_n_420__33_;
      r_420__32_ <= r_n_420__32_;
      r_420__31_ <= r_n_420__31_;
      r_420__30_ <= r_n_420__30_;
      r_420__29_ <= r_n_420__29_;
      r_420__28_ <= r_n_420__28_;
      r_420__27_ <= r_n_420__27_;
      r_420__26_ <= r_n_420__26_;
      r_420__25_ <= r_n_420__25_;
      r_420__24_ <= r_n_420__24_;
      r_420__23_ <= r_n_420__23_;
      r_420__22_ <= r_n_420__22_;
      r_420__21_ <= r_n_420__21_;
      r_420__20_ <= r_n_420__20_;
      r_420__19_ <= r_n_420__19_;
      r_420__18_ <= r_n_420__18_;
      r_420__17_ <= r_n_420__17_;
      r_420__16_ <= r_n_420__16_;
      r_420__15_ <= r_n_420__15_;
      r_420__14_ <= r_n_420__14_;
      r_420__13_ <= r_n_420__13_;
      r_420__12_ <= r_n_420__12_;
      r_420__11_ <= r_n_420__11_;
      r_420__10_ <= r_n_420__10_;
      r_420__9_ <= r_n_420__9_;
      r_420__8_ <= r_n_420__8_;
      r_420__7_ <= r_n_420__7_;
      r_420__6_ <= r_n_420__6_;
      r_420__5_ <= r_n_420__5_;
      r_420__4_ <= r_n_420__4_;
      r_420__3_ <= r_n_420__3_;
      r_420__2_ <= r_n_420__2_;
      r_420__1_ <= r_n_420__1_;
      r_420__0_ <= r_n_420__0_;
    end 
    if(N4005) begin
      r_421__63_ <= r_n_421__63_;
      r_421__62_ <= r_n_421__62_;
      r_421__61_ <= r_n_421__61_;
      r_421__60_ <= r_n_421__60_;
      r_421__59_ <= r_n_421__59_;
      r_421__58_ <= r_n_421__58_;
      r_421__57_ <= r_n_421__57_;
      r_421__56_ <= r_n_421__56_;
      r_421__55_ <= r_n_421__55_;
      r_421__54_ <= r_n_421__54_;
      r_421__53_ <= r_n_421__53_;
      r_421__52_ <= r_n_421__52_;
      r_421__51_ <= r_n_421__51_;
      r_421__50_ <= r_n_421__50_;
      r_421__49_ <= r_n_421__49_;
      r_421__48_ <= r_n_421__48_;
      r_421__47_ <= r_n_421__47_;
      r_421__46_ <= r_n_421__46_;
      r_421__45_ <= r_n_421__45_;
      r_421__44_ <= r_n_421__44_;
      r_421__43_ <= r_n_421__43_;
      r_421__42_ <= r_n_421__42_;
      r_421__41_ <= r_n_421__41_;
      r_421__40_ <= r_n_421__40_;
      r_421__39_ <= r_n_421__39_;
      r_421__38_ <= r_n_421__38_;
      r_421__37_ <= r_n_421__37_;
      r_421__36_ <= r_n_421__36_;
      r_421__35_ <= r_n_421__35_;
      r_421__34_ <= r_n_421__34_;
      r_421__33_ <= r_n_421__33_;
      r_421__32_ <= r_n_421__32_;
      r_421__31_ <= r_n_421__31_;
      r_421__30_ <= r_n_421__30_;
      r_421__29_ <= r_n_421__29_;
      r_421__28_ <= r_n_421__28_;
      r_421__27_ <= r_n_421__27_;
      r_421__26_ <= r_n_421__26_;
      r_421__25_ <= r_n_421__25_;
      r_421__24_ <= r_n_421__24_;
      r_421__23_ <= r_n_421__23_;
      r_421__22_ <= r_n_421__22_;
      r_421__21_ <= r_n_421__21_;
      r_421__20_ <= r_n_421__20_;
      r_421__19_ <= r_n_421__19_;
      r_421__18_ <= r_n_421__18_;
      r_421__17_ <= r_n_421__17_;
      r_421__16_ <= r_n_421__16_;
      r_421__15_ <= r_n_421__15_;
      r_421__14_ <= r_n_421__14_;
      r_421__13_ <= r_n_421__13_;
      r_421__12_ <= r_n_421__12_;
      r_421__11_ <= r_n_421__11_;
      r_421__10_ <= r_n_421__10_;
      r_421__9_ <= r_n_421__9_;
      r_421__8_ <= r_n_421__8_;
      r_421__7_ <= r_n_421__7_;
      r_421__6_ <= r_n_421__6_;
      r_421__5_ <= r_n_421__5_;
      r_421__4_ <= r_n_421__4_;
      r_421__3_ <= r_n_421__3_;
      r_421__2_ <= r_n_421__2_;
      r_421__1_ <= r_n_421__1_;
      r_421__0_ <= r_n_421__0_;
    end 
    if(N4006) begin
      r_422__63_ <= r_n_422__63_;
      r_422__62_ <= r_n_422__62_;
      r_422__61_ <= r_n_422__61_;
      r_422__60_ <= r_n_422__60_;
      r_422__59_ <= r_n_422__59_;
      r_422__58_ <= r_n_422__58_;
      r_422__57_ <= r_n_422__57_;
      r_422__56_ <= r_n_422__56_;
      r_422__55_ <= r_n_422__55_;
      r_422__54_ <= r_n_422__54_;
      r_422__53_ <= r_n_422__53_;
      r_422__52_ <= r_n_422__52_;
      r_422__51_ <= r_n_422__51_;
      r_422__50_ <= r_n_422__50_;
      r_422__49_ <= r_n_422__49_;
      r_422__48_ <= r_n_422__48_;
      r_422__47_ <= r_n_422__47_;
      r_422__46_ <= r_n_422__46_;
      r_422__45_ <= r_n_422__45_;
      r_422__44_ <= r_n_422__44_;
      r_422__43_ <= r_n_422__43_;
      r_422__42_ <= r_n_422__42_;
      r_422__41_ <= r_n_422__41_;
      r_422__40_ <= r_n_422__40_;
      r_422__39_ <= r_n_422__39_;
      r_422__38_ <= r_n_422__38_;
      r_422__37_ <= r_n_422__37_;
      r_422__36_ <= r_n_422__36_;
      r_422__35_ <= r_n_422__35_;
      r_422__34_ <= r_n_422__34_;
      r_422__33_ <= r_n_422__33_;
      r_422__32_ <= r_n_422__32_;
      r_422__31_ <= r_n_422__31_;
      r_422__30_ <= r_n_422__30_;
      r_422__29_ <= r_n_422__29_;
      r_422__28_ <= r_n_422__28_;
      r_422__27_ <= r_n_422__27_;
      r_422__26_ <= r_n_422__26_;
      r_422__25_ <= r_n_422__25_;
      r_422__24_ <= r_n_422__24_;
      r_422__23_ <= r_n_422__23_;
      r_422__22_ <= r_n_422__22_;
      r_422__21_ <= r_n_422__21_;
      r_422__20_ <= r_n_422__20_;
      r_422__19_ <= r_n_422__19_;
      r_422__18_ <= r_n_422__18_;
      r_422__17_ <= r_n_422__17_;
      r_422__16_ <= r_n_422__16_;
      r_422__15_ <= r_n_422__15_;
      r_422__14_ <= r_n_422__14_;
      r_422__13_ <= r_n_422__13_;
      r_422__12_ <= r_n_422__12_;
      r_422__11_ <= r_n_422__11_;
      r_422__10_ <= r_n_422__10_;
      r_422__9_ <= r_n_422__9_;
      r_422__8_ <= r_n_422__8_;
      r_422__7_ <= r_n_422__7_;
      r_422__6_ <= r_n_422__6_;
      r_422__5_ <= r_n_422__5_;
      r_422__4_ <= r_n_422__4_;
      r_422__3_ <= r_n_422__3_;
      r_422__2_ <= r_n_422__2_;
      r_422__1_ <= r_n_422__1_;
      r_422__0_ <= r_n_422__0_;
    end 
    if(N4007) begin
      r_423__63_ <= r_n_423__63_;
      r_423__62_ <= r_n_423__62_;
      r_423__61_ <= r_n_423__61_;
      r_423__60_ <= r_n_423__60_;
      r_423__59_ <= r_n_423__59_;
      r_423__58_ <= r_n_423__58_;
      r_423__57_ <= r_n_423__57_;
      r_423__56_ <= r_n_423__56_;
      r_423__55_ <= r_n_423__55_;
      r_423__54_ <= r_n_423__54_;
      r_423__53_ <= r_n_423__53_;
      r_423__52_ <= r_n_423__52_;
      r_423__51_ <= r_n_423__51_;
      r_423__50_ <= r_n_423__50_;
      r_423__49_ <= r_n_423__49_;
      r_423__48_ <= r_n_423__48_;
      r_423__47_ <= r_n_423__47_;
      r_423__46_ <= r_n_423__46_;
      r_423__45_ <= r_n_423__45_;
      r_423__44_ <= r_n_423__44_;
      r_423__43_ <= r_n_423__43_;
      r_423__42_ <= r_n_423__42_;
      r_423__41_ <= r_n_423__41_;
      r_423__40_ <= r_n_423__40_;
      r_423__39_ <= r_n_423__39_;
      r_423__38_ <= r_n_423__38_;
      r_423__37_ <= r_n_423__37_;
      r_423__36_ <= r_n_423__36_;
      r_423__35_ <= r_n_423__35_;
      r_423__34_ <= r_n_423__34_;
      r_423__33_ <= r_n_423__33_;
      r_423__32_ <= r_n_423__32_;
      r_423__31_ <= r_n_423__31_;
      r_423__30_ <= r_n_423__30_;
      r_423__29_ <= r_n_423__29_;
      r_423__28_ <= r_n_423__28_;
      r_423__27_ <= r_n_423__27_;
      r_423__26_ <= r_n_423__26_;
      r_423__25_ <= r_n_423__25_;
      r_423__24_ <= r_n_423__24_;
      r_423__23_ <= r_n_423__23_;
      r_423__22_ <= r_n_423__22_;
      r_423__21_ <= r_n_423__21_;
      r_423__20_ <= r_n_423__20_;
      r_423__19_ <= r_n_423__19_;
      r_423__18_ <= r_n_423__18_;
      r_423__17_ <= r_n_423__17_;
      r_423__16_ <= r_n_423__16_;
      r_423__15_ <= r_n_423__15_;
      r_423__14_ <= r_n_423__14_;
      r_423__13_ <= r_n_423__13_;
      r_423__12_ <= r_n_423__12_;
      r_423__11_ <= r_n_423__11_;
      r_423__10_ <= r_n_423__10_;
      r_423__9_ <= r_n_423__9_;
      r_423__8_ <= r_n_423__8_;
      r_423__7_ <= r_n_423__7_;
      r_423__6_ <= r_n_423__6_;
      r_423__5_ <= r_n_423__5_;
      r_423__4_ <= r_n_423__4_;
      r_423__3_ <= r_n_423__3_;
      r_423__2_ <= r_n_423__2_;
      r_423__1_ <= r_n_423__1_;
      r_423__0_ <= r_n_423__0_;
    end 
    if(N4008) begin
      r_424__63_ <= r_n_424__63_;
      r_424__62_ <= r_n_424__62_;
      r_424__61_ <= r_n_424__61_;
      r_424__60_ <= r_n_424__60_;
      r_424__59_ <= r_n_424__59_;
      r_424__58_ <= r_n_424__58_;
      r_424__57_ <= r_n_424__57_;
      r_424__56_ <= r_n_424__56_;
      r_424__55_ <= r_n_424__55_;
      r_424__54_ <= r_n_424__54_;
      r_424__53_ <= r_n_424__53_;
      r_424__52_ <= r_n_424__52_;
      r_424__51_ <= r_n_424__51_;
      r_424__50_ <= r_n_424__50_;
      r_424__49_ <= r_n_424__49_;
      r_424__48_ <= r_n_424__48_;
      r_424__47_ <= r_n_424__47_;
      r_424__46_ <= r_n_424__46_;
      r_424__45_ <= r_n_424__45_;
      r_424__44_ <= r_n_424__44_;
      r_424__43_ <= r_n_424__43_;
      r_424__42_ <= r_n_424__42_;
      r_424__41_ <= r_n_424__41_;
      r_424__40_ <= r_n_424__40_;
      r_424__39_ <= r_n_424__39_;
      r_424__38_ <= r_n_424__38_;
      r_424__37_ <= r_n_424__37_;
      r_424__36_ <= r_n_424__36_;
      r_424__35_ <= r_n_424__35_;
      r_424__34_ <= r_n_424__34_;
      r_424__33_ <= r_n_424__33_;
      r_424__32_ <= r_n_424__32_;
      r_424__31_ <= r_n_424__31_;
      r_424__30_ <= r_n_424__30_;
      r_424__29_ <= r_n_424__29_;
      r_424__28_ <= r_n_424__28_;
      r_424__27_ <= r_n_424__27_;
      r_424__26_ <= r_n_424__26_;
      r_424__25_ <= r_n_424__25_;
      r_424__24_ <= r_n_424__24_;
      r_424__23_ <= r_n_424__23_;
      r_424__22_ <= r_n_424__22_;
      r_424__21_ <= r_n_424__21_;
      r_424__20_ <= r_n_424__20_;
      r_424__19_ <= r_n_424__19_;
      r_424__18_ <= r_n_424__18_;
      r_424__17_ <= r_n_424__17_;
      r_424__16_ <= r_n_424__16_;
      r_424__15_ <= r_n_424__15_;
      r_424__14_ <= r_n_424__14_;
      r_424__13_ <= r_n_424__13_;
      r_424__12_ <= r_n_424__12_;
      r_424__11_ <= r_n_424__11_;
      r_424__10_ <= r_n_424__10_;
      r_424__9_ <= r_n_424__9_;
      r_424__8_ <= r_n_424__8_;
      r_424__7_ <= r_n_424__7_;
      r_424__6_ <= r_n_424__6_;
      r_424__5_ <= r_n_424__5_;
      r_424__4_ <= r_n_424__4_;
      r_424__3_ <= r_n_424__3_;
      r_424__2_ <= r_n_424__2_;
      r_424__1_ <= r_n_424__1_;
      r_424__0_ <= r_n_424__0_;
    end 
    if(N4009) begin
      r_425__63_ <= r_n_425__63_;
      r_425__62_ <= r_n_425__62_;
      r_425__61_ <= r_n_425__61_;
      r_425__60_ <= r_n_425__60_;
      r_425__59_ <= r_n_425__59_;
      r_425__58_ <= r_n_425__58_;
      r_425__57_ <= r_n_425__57_;
      r_425__56_ <= r_n_425__56_;
      r_425__55_ <= r_n_425__55_;
      r_425__54_ <= r_n_425__54_;
      r_425__53_ <= r_n_425__53_;
      r_425__52_ <= r_n_425__52_;
      r_425__51_ <= r_n_425__51_;
      r_425__50_ <= r_n_425__50_;
      r_425__49_ <= r_n_425__49_;
      r_425__48_ <= r_n_425__48_;
      r_425__47_ <= r_n_425__47_;
      r_425__46_ <= r_n_425__46_;
      r_425__45_ <= r_n_425__45_;
      r_425__44_ <= r_n_425__44_;
      r_425__43_ <= r_n_425__43_;
      r_425__42_ <= r_n_425__42_;
      r_425__41_ <= r_n_425__41_;
      r_425__40_ <= r_n_425__40_;
      r_425__39_ <= r_n_425__39_;
      r_425__38_ <= r_n_425__38_;
      r_425__37_ <= r_n_425__37_;
      r_425__36_ <= r_n_425__36_;
      r_425__35_ <= r_n_425__35_;
      r_425__34_ <= r_n_425__34_;
      r_425__33_ <= r_n_425__33_;
      r_425__32_ <= r_n_425__32_;
      r_425__31_ <= r_n_425__31_;
      r_425__30_ <= r_n_425__30_;
      r_425__29_ <= r_n_425__29_;
      r_425__28_ <= r_n_425__28_;
      r_425__27_ <= r_n_425__27_;
      r_425__26_ <= r_n_425__26_;
      r_425__25_ <= r_n_425__25_;
      r_425__24_ <= r_n_425__24_;
      r_425__23_ <= r_n_425__23_;
      r_425__22_ <= r_n_425__22_;
      r_425__21_ <= r_n_425__21_;
      r_425__20_ <= r_n_425__20_;
      r_425__19_ <= r_n_425__19_;
      r_425__18_ <= r_n_425__18_;
      r_425__17_ <= r_n_425__17_;
      r_425__16_ <= r_n_425__16_;
      r_425__15_ <= r_n_425__15_;
      r_425__14_ <= r_n_425__14_;
      r_425__13_ <= r_n_425__13_;
      r_425__12_ <= r_n_425__12_;
      r_425__11_ <= r_n_425__11_;
      r_425__10_ <= r_n_425__10_;
      r_425__9_ <= r_n_425__9_;
      r_425__8_ <= r_n_425__8_;
      r_425__7_ <= r_n_425__7_;
      r_425__6_ <= r_n_425__6_;
      r_425__5_ <= r_n_425__5_;
      r_425__4_ <= r_n_425__4_;
      r_425__3_ <= r_n_425__3_;
      r_425__2_ <= r_n_425__2_;
      r_425__1_ <= r_n_425__1_;
      r_425__0_ <= r_n_425__0_;
    end 
    if(N4010) begin
      r_426__63_ <= r_n_426__63_;
      r_426__62_ <= r_n_426__62_;
      r_426__61_ <= r_n_426__61_;
      r_426__60_ <= r_n_426__60_;
      r_426__59_ <= r_n_426__59_;
      r_426__58_ <= r_n_426__58_;
      r_426__57_ <= r_n_426__57_;
      r_426__56_ <= r_n_426__56_;
      r_426__55_ <= r_n_426__55_;
      r_426__54_ <= r_n_426__54_;
      r_426__53_ <= r_n_426__53_;
      r_426__52_ <= r_n_426__52_;
      r_426__51_ <= r_n_426__51_;
      r_426__50_ <= r_n_426__50_;
      r_426__49_ <= r_n_426__49_;
      r_426__48_ <= r_n_426__48_;
      r_426__47_ <= r_n_426__47_;
      r_426__46_ <= r_n_426__46_;
      r_426__45_ <= r_n_426__45_;
      r_426__44_ <= r_n_426__44_;
      r_426__43_ <= r_n_426__43_;
      r_426__42_ <= r_n_426__42_;
      r_426__41_ <= r_n_426__41_;
      r_426__40_ <= r_n_426__40_;
      r_426__39_ <= r_n_426__39_;
      r_426__38_ <= r_n_426__38_;
      r_426__37_ <= r_n_426__37_;
      r_426__36_ <= r_n_426__36_;
      r_426__35_ <= r_n_426__35_;
      r_426__34_ <= r_n_426__34_;
      r_426__33_ <= r_n_426__33_;
      r_426__32_ <= r_n_426__32_;
      r_426__31_ <= r_n_426__31_;
      r_426__30_ <= r_n_426__30_;
      r_426__29_ <= r_n_426__29_;
      r_426__28_ <= r_n_426__28_;
      r_426__27_ <= r_n_426__27_;
      r_426__26_ <= r_n_426__26_;
      r_426__25_ <= r_n_426__25_;
      r_426__24_ <= r_n_426__24_;
      r_426__23_ <= r_n_426__23_;
      r_426__22_ <= r_n_426__22_;
      r_426__21_ <= r_n_426__21_;
      r_426__20_ <= r_n_426__20_;
      r_426__19_ <= r_n_426__19_;
      r_426__18_ <= r_n_426__18_;
      r_426__17_ <= r_n_426__17_;
      r_426__16_ <= r_n_426__16_;
      r_426__15_ <= r_n_426__15_;
      r_426__14_ <= r_n_426__14_;
      r_426__13_ <= r_n_426__13_;
      r_426__12_ <= r_n_426__12_;
      r_426__11_ <= r_n_426__11_;
      r_426__10_ <= r_n_426__10_;
      r_426__9_ <= r_n_426__9_;
      r_426__8_ <= r_n_426__8_;
      r_426__7_ <= r_n_426__7_;
      r_426__6_ <= r_n_426__6_;
      r_426__5_ <= r_n_426__5_;
      r_426__4_ <= r_n_426__4_;
      r_426__3_ <= r_n_426__3_;
      r_426__2_ <= r_n_426__2_;
      r_426__1_ <= r_n_426__1_;
      r_426__0_ <= r_n_426__0_;
    end 
    if(N4011) begin
      r_427__63_ <= r_n_427__63_;
      r_427__62_ <= r_n_427__62_;
      r_427__61_ <= r_n_427__61_;
      r_427__60_ <= r_n_427__60_;
      r_427__59_ <= r_n_427__59_;
      r_427__58_ <= r_n_427__58_;
      r_427__57_ <= r_n_427__57_;
      r_427__56_ <= r_n_427__56_;
      r_427__55_ <= r_n_427__55_;
      r_427__54_ <= r_n_427__54_;
      r_427__53_ <= r_n_427__53_;
      r_427__52_ <= r_n_427__52_;
      r_427__51_ <= r_n_427__51_;
      r_427__50_ <= r_n_427__50_;
      r_427__49_ <= r_n_427__49_;
      r_427__48_ <= r_n_427__48_;
      r_427__47_ <= r_n_427__47_;
      r_427__46_ <= r_n_427__46_;
      r_427__45_ <= r_n_427__45_;
      r_427__44_ <= r_n_427__44_;
      r_427__43_ <= r_n_427__43_;
      r_427__42_ <= r_n_427__42_;
      r_427__41_ <= r_n_427__41_;
      r_427__40_ <= r_n_427__40_;
      r_427__39_ <= r_n_427__39_;
      r_427__38_ <= r_n_427__38_;
      r_427__37_ <= r_n_427__37_;
      r_427__36_ <= r_n_427__36_;
      r_427__35_ <= r_n_427__35_;
      r_427__34_ <= r_n_427__34_;
      r_427__33_ <= r_n_427__33_;
      r_427__32_ <= r_n_427__32_;
      r_427__31_ <= r_n_427__31_;
      r_427__30_ <= r_n_427__30_;
      r_427__29_ <= r_n_427__29_;
      r_427__28_ <= r_n_427__28_;
      r_427__27_ <= r_n_427__27_;
      r_427__26_ <= r_n_427__26_;
      r_427__25_ <= r_n_427__25_;
      r_427__24_ <= r_n_427__24_;
      r_427__23_ <= r_n_427__23_;
      r_427__22_ <= r_n_427__22_;
      r_427__21_ <= r_n_427__21_;
      r_427__20_ <= r_n_427__20_;
      r_427__19_ <= r_n_427__19_;
      r_427__18_ <= r_n_427__18_;
      r_427__17_ <= r_n_427__17_;
      r_427__16_ <= r_n_427__16_;
      r_427__15_ <= r_n_427__15_;
      r_427__14_ <= r_n_427__14_;
      r_427__13_ <= r_n_427__13_;
      r_427__12_ <= r_n_427__12_;
      r_427__11_ <= r_n_427__11_;
      r_427__10_ <= r_n_427__10_;
      r_427__9_ <= r_n_427__9_;
      r_427__8_ <= r_n_427__8_;
      r_427__7_ <= r_n_427__7_;
      r_427__6_ <= r_n_427__6_;
      r_427__5_ <= r_n_427__5_;
      r_427__4_ <= r_n_427__4_;
      r_427__3_ <= r_n_427__3_;
      r_427__2_ <= r_n_427__2_;
      r_427__1_ <= r_n_427__1_;
      r_427__0_ <= r_n_427__0_;
    end 
    if(N4012) begin
      r_428__63_ <= r_n_428__63_;
      r_428__62_ <= r_n_428__62_;
      r_428__61_ <= r_n_428__61_;
      r_428__60_ <= r_n_428__60_;
      r_428__59_ <= r_n_428__59_;
      r_428__58_ <= r_n_428__58_;
      r_428__57_ <= r_n_428__57_;
      r_428__56_ <= r_n_428__56_;
      r_428__55_ <= r_n_428__55_;
      r_428__54_ <= r_n_428__54_;
      r_428__53_ <= r_n_428__53_;
      r_428__52_ <= r_n_428__52_;
      r_428__51_ <= r_n_428__51_;
      r_428__50_ <= r_n_428__50_;
      r_428__49_ <= r_n_428__49_;
      r_428__48_ <= r_n_428__48_;
      r_428__47_ <= r_n_428__47_;
      r_428__46_ <= r_n_428__46_;
      r_428__45_ <= r_n_428__45_;
      r_428__44_ <= r_n_428__44_;
      r_428__43_ <= r_n_428__43_;
      r_428__42_ <= r_n_428__42_;
      r_428__41_ <= r_n_428__41_;
      r_428__40_ <= r_n_428__40_;
      r_428__39_ <= r_n_428__39_;
      r_428__38_ <= r_n_428__38_;
      r_428__37_ <= r_n_428__37_;
      r_428__36_ <= r_n_428__36_;
      r_428__35_ <= r_n_428__35_;
      r_428__34_ <= r_n_428__34_;
      r_428__33_ <= r_n_428__33_;
      r_428__32_ <= r_n_428__32_;
      r_428__31_ <= r_n_428__31_;
      r_428__30_ <= r_n_428__30_;
      r_428__29_ <= r_n_428__29_;
      r_428__28_ <= r_n_428__28_;
      r_428__27_ <= r_n_428__27_;
      r_428__26_ <= r_n_428__26_;
      r_428__25_ <= r_n_428__25_;
      r_428__24_ <= r_n_428__24_;
      r_428__23_ <= r_n_428__23_;
      r_428__22_ <= r_n_428__22_;
      r_428__21_ <= r_n_428__21_;
      r_428__20_ <= r_n_428__20_;
      r_428__19_ <= r_n_428__19_;
      r_428__18_ <= r_n_428__18_;
      r_428__17_ <= r_n_428__17_;
      r_428__16_ <= r_n_428__16_;
      r_428__15_ <= r_n_428__15_;
      r_428__14_ <= r_n_428__14_;
      r_428__13_ <= r_n_428__13_;
      r_428__12_ <= r_n_428__12_;
      r_428__11_ <= r_n_428__11_;
      r_428__10_ <= r_n_428__10_;
      r_428__9_ <= r_n_428__9_;
      r_428__8_ <= r_n_428__8_;
      r_428__7_ <= r_n_428__7_;
      r_428__6_ <= r_n_428__6_;
      r_428__5_ <= r_n_428__5_;
      r_428__4_ <= r_n_428__4_;
      r_428__3_ <= r_n_428__3_;
      r_428__2_ <= r_n_428__2_;
      r_428__1_ <= r_n_428__1_;
      r_428__0_ <= r_n_428__0_;
    end 
    if(N4013) begin
      r_429__63_ <= r_n_429__63_;
      r_429__62_ <= r_n_429__62_;
      r_429__61_ <= r_n_429__61_;
      r_429__60_ <= r_n_429__60_;
      r_429__59_ <= r_n_429__59_;
      r_429__58_ <= r_n_429__58_;
      r_429__57_ <= r_n_429__57_;
      r_429__56_ <= r_n_429__56_;
      r_429__55_ <= r_n_429__55_;
      r_429__54_ <= r_n_429__54_;
      r_429__53_ <= r_n_429__53_;
      r_429__52_ <= r_n_429__52_;
      r_429__51_ <= r_n_429__51_;
      r_429__50_ <= r_n_429__50_;
      r_429__49_ <= r_n_429__49_;
      r_429__48_ <= r_n_429__48_;
      r_429__47_ <= r_n_429__47_;
      r_429__46_ <= r_n_429__46_;
      r_429__45_ <= r_n_429__45_;
      r_429__44_ <= r_n_429__44_;
      r_429__43_ <= r_n_429__43_;
      r_429__42_ <= r_n_429__42_;
      r_429__41_ <= r_n_429__41_;
      r_429__40_ <= r_n_429__40_;
      r_429__39_ <= r_n_429__39_;
      r_429__38_ <= r_n_429__38_;
      r_429__37_ <= r_n_429__37_;
      r_429__36_ <= r_n_429__36_;
      r_429__35_ <= r_n_429__35_;
      r_429__34_ <= r_n_429__34_;
      r_429__33_ <= r_n_429__33_;
      r_429__32_ <= r_n_429__32_;
      r_429__31_ <= r_n_429__31_;
      r_429__30_ <= r_n_429__30_;
      r_429__29_ <= r_n_429__29_;
      r_429__28_ <= r_n_429__28_;
      r_429__27_ <= r_n_429__27_;
      r_429__26_ <= r_n_429__26_;
      r_429__25_ <= r_n_429__25_;
      r_429__24_ <= r_n_429__24_;
      r_429__23_ <= r_n_429__23_;
      r_429__22_ <= r_n_429__22_;
      r_429__21_ <= r_n_429__21_;
      r_429__20_ <= r_n_429__20_;
      r_429__19_ <= r_n_429__19_;
      r_429__18_ <= r_n_429__18_;
      r_429__17_ <= r_n_429__17_;
      r_429__16_ <= r_n_429__16_;
      r_429__15_ <= r_n_429__15_;
      r_429__14_ <= r_n_429__14_;
      r_429__13_ <= r_n_429__13_;
      r_429__12_ <= r_n_429__12_;
      r_429__11_ <= r_n_429__11_;
      r_429__10_ <= r_n_429__10_;
      r_429__9_ <= r_n_429__9_;
      r_429__8_ <= r_n_429__8_;
      r_429__7_ <= r_n_429__7_;
      r_429__6_ <= r_n_429__6_;
      r_429__5_ <= r_n_429__5_;
      r_429__4_ <= r_n_429__4_;
      r_429__3_ <= r_n_429__3_;
      r_429__2_ <= r_n_429__2_;
      r_429__1_ <= r_n_429__1_;
      r_429__0_ <= r_n_429__0_;
    end 
    if(N4014) begin
      r_430__63_ <= r_n_430__63_;
      r_430__62_ <= r_n_430__62_;
      r_430__61_ <= r_n_430__61_;
      r_430__60_ <= r_n_430__60_;
      r_430__59_ <= r_n_430__59_;
      r_430__58_ <= r_n_430__58_;
      r_430__57_ <= r_n_430__57_;
      r_430__56_ <= r_n_430__56_;
      r_430__55_ <= r_n_430__55_;
      r_430__54_ <= r_n_430__54_;
      r_430__53_ <= r_n_430__53_;
      r_430__52_ <= r_n_430__52_;
      r_430__51_ <= r_n_430__51_;
      r_430__50_ <= r_n_430__50_;
      r_430__49_ <= r_n_430__49_;
      r_430__48_ <= r_n_430__48_;
      r_430__47_ <= r_n_430__47_;
      r_430__46_ <= r_n_430__46_;
      r_430__45_ <= r_n_430__45_;
      r_430__44_ <= r_n_430__44_;
      r_430__43_ <= r_n_430__43_;
      r_430__42_ <= r_n_430__42_;
      r_430__41_ <= r_n_430__41_;
      r_430__40_ <= r_n_430__40_;
      r_430__39_ <= r_n_430__39_;
      r_430__38_ <= r_n_430__38_;
      r_430__37_ <= r_n_430__37_;
      r_430__36_ <= r_n_430__36_;
      r_430__35_ <= r_n_430__35_;
      r_430__34_ <= r_n_430__34_;
      r_430__33_ <= r_n_430__33_;
      r_430__32_ <= r_n_430__32_;
      r_430__31_ <= r_n_430__31_;
      r_430__30_ <= r_n_430__30_;
      r_430__29_ <= r_n_430__29_;
      r_430__28_ <= r_n_430__28_;
      r_430__27_ <= r_n_430__27_;
      r_430__26_ <= r_n_430__26_;
      r_430__25_ <= r_n_430__25_;
      r_430__24_ <= r_n_430__24_;
      r_430__23_ <= r_n_430__23_;
      r_430__22_ <= r_n_430__22_;
      r_430__21_ <= r_n_430__21_;
      r_430__20_ <= r_n_430__20_;
      r_430__19_ <= r_n_430__19_;
      r_430__18_ <= r_n_430__18_;
      r_430__17_ <= r_n_430__17_;
      r_430__16_ <= r_n_430__16_;
      r_430__15_ <= r_n_430__15_;
      r_430__14_ <= r_n_430__14_;
      r_430__13_ <= r_n_430__13_;
      r_430__12_ <= r_n_430__12_;
      r_430__11_ <= r_n_430__11_;
      r_430__10_ <= r_n_430__10_;
      r_430__9_ <= r_n_430__9_;
      r_430__8_ <= r_n_430__8_;
      r_430__7_ <= r_n_430__7_;
      r_430__6_ <= r_n_430__6_;
      r_430__5_ <= r_n_430__5_;
      r_430__4_ <= r_n_430__4_;
      r_430__3_ <= r_n_430__3_;
      r_430__2_ <= r_n_430__2_;
      r_430__1_ <= r_n_430__1_;
      r_430__0_ <= r_n_430__0_;
    end 
    if(N4015) begin
      r_431__63_ <= r_n_431__63_;
      r_431__62_ <= r_n_431__62_;
      r_431__61_ <= r_n_431__61_;
      r_431__60_ <= r_n_431__60_;
      r_431__59_ <= r_n_431__59_;
      r_431__58_ <= r_n_431__58_;
      r_431__57_ <= r_n_431__57_;
      r_431__56_ <= r_n_431__56_;
      r_431__55_ <= r_n_431__55_;
      r_431__54_ <= r_n_431__54_;
      r_431__53_ <= r_n_431__53_;
      r_431__52_ <= r_n_431__52_;
      r_431__51_ <= r_n_431__51_;
      r_431__50_ <= r_n_431__50_;
      r_431__49_ <= r_n_431__49_;
      r_431__48_ <= r_n_431__48_;
      r_431__47_ <= r_n_431__47_;
      r_431__46_ <= r_n_431__46_;
      r_431__45_ <= r_n_431__45_;
      r_431__44_ <= r_n_431__44_;
      r_431__43_ <= r_n_431__43_;
      r_431__42_ <= r_n_431__42_;
      r_431__41_ <= r_n_431__41_;
      r_431__40_ <= r_n_431__40_;
      r_431__39_ <= r_n_431__39_;
      r_431__38_ <= r_n_431__38_;
      r_431__37_ <= r_n_431__37_;
      r_431__36_ <= r_n_431__36_;
      r_431__35_ <= r_n_431__35_;
      r_431__34_ <= r_n_431__34_;
      r_431__33_ <= r_n_431__33_;
      r_431__32_ <= r_n_431__32_;
      r_431__31_ <= r_n_431__31_;
      r_431__30_ <= r_n_431__30_;
      r_431__29_ <= r_n_431__29_;
      r_431__28_ <= r_n_431__28_;
      r_431__27_ <= r_n_431__27_;
      r_431__26_ <= r_n_431__26_;
      r_431__25_ <= r_n_431__25_;
      r_431__24_ <= r_n_431__24_;
      r_431__23_ <= r_n_431__23_;
      r_431__22_ <= r_n_431__22_;
      r_431__21_ <= r_n_431__21_;
      r_431__20_ <= r_n_431__20_;
      r_431__19_ <= r_n_431__19_;
      r_431__18_ <= r_n_431__18_;
      r_431__17_ <= r_n_431__17_;
      r_431__16_ <= r_n_431__16_;
      r_431__15_ <= r_n_431__15_;
      r_431__14_ <= r_n_431__14_;
      r_431__13_ <= r_n_431__13_;
      r_431__12_ <= r_n_431__12_;
      r_431__11_ <= r_n_431__11_;
      r_431__10_ <= r_n_431__10_;
      r_431__9_ <= r_n_431__9_;
      r_431__8_ <= r_n_431__8_;
      r_431__7_ <= r_n_431__7_;
      r_431__6_ <= r_n_431__6_;
      r_431__5_ <= r_n_431__5_;
      r_431__4_ <= r_n_431__4_;
      r_431__3_ <= r_n_431__3_;
      r_431__2_ <= r_n_431__2_;
      r_431__1_ <= r_n_431__1_;
      r_431__0_ <= r_n_431__0_;
    end 
    if(N4016) begin
      r_432__63_ <= r_n_432__63_;
      r_432__62_ <= r_n_432__62_;
      r_432__61_ <= r_n_432__61_;
      r_432__60_ <= r_n_432__60_;
      r_432__59_ <= r_n_432__59_;
      r_432__58_ <= r_n_432__58_;
      r_432__57_ <= r_n_432__57_;
      r_432__56_ <= r_n_432__56_;
      r_432__55_ <= r_n_432__55_;
      r_432__54_ <= r_n_432__54_;
      r_432__53_ <= r_n_432__53_;
      r_432__52_ <= r_n_432__52_;
      r_432__51_ <= r_n_432__51_;
      r_432__50_ <= r_n_432__50_;
      r_432__49_ <= r_n_432__49_;
      r_432__48_ <= r_n_432__48_;
      r_432__47_ <= r_n_432__47_;
      r_432__46_ <= r_n_432__46_;
      r_432__45_ <= r_n_432__45_;
      r_432__44_ <= r_n_432__44_;
      r_432__43_ <= r_n_432__43_;
      r_432__42_ <= r_n_432__42_;
      r_432__41_ <= r_n_432__41_;
      r_432__40_ <= r_n_432__40_;
      r_432__39_ <= r_n_432__39_;
      r_432__38_ <= r_n_432__38_;
      r_432__37_ <= r_n_432__37_;
      r_432__36_ <= r_n_432__36_;
      r_432__35_ <= r_n_432__35_;
      r_432__34_ <= r_n_432__34_;
      r_432__33_ <= r_n_432__33_;
      r_432__32_ <= r_n_432__32_;
      r_432__31_ <= r_n_432__31_;
      r_432__30_ <= r_n_432__30_;
      r_432__29_ <= r_n_432__29_;
      r_432__28_ <= r_n_432__28_;
      r_432__27_ <= r_n_432__27_;
      r_432__26_ <= r_n_432__26_;
      r_432__25_ <= r_n_432__25_;
      r_432__24_ <= r_n_432__24_;
      r_432__23_ <= r_n_432__23_;
      r_432__22_ <= r_n_432__22_;
      r_432__21_ <= r_n_432__21_;
      r_432__20_ <= r_n_432__20_;
      r_432__19_ <= r_n_432__19_;
      r_432__18_ <= r_n_432__18_;
      r_432__17_ <= r_n_432__17_;
      r_432__16_ <= r_n_432__16_;
      r_432__15_ <= r_n_432__15_;
      r_432__14_ <= r_n_432__14_;
      r_432__13_ <= r_n_432__13_;
      r_432__12_ <= r_n_432__12_;
      r_432__11_ <= r_n_432__11_;
      r_432__10_ <= r_n_432__10_;
      r_432__9_ <= r_n_432__9_;
      r_432__8_ <= r_n_432__8_;
      r_432__7_ <= r_n_432__7_;
      r_432__6_ <= r_n_432__6_;
      r_432__5_ <= r_n_432__5_;
      r_432__4_ <= r_n_432__4_;
      r_432__3_ <= r_n_432__3_;
      r_432__2_ <= r_n_432__2_;
      r_432__1_ <= r_n_432__1_;
      r_432__0_ <= r_n_432__0_;
    end 
    if(N4017) begin
      r_433__63_ <= r_n_433__63_;
      r_433__62_ <= r_n_433__62_;
      r_433__61_ <= r_n_433__61_;
      r_433__60_ <= r_n_433__60_;
      r_433__59_ <= r_n_433__59_;
      r_433__58_ <= r_n_433__58_;
      r_433__57_ <= r_n_433__57_;
      r_433__56_ <= r_n_433__56_;
      r_433__55_ <= r_n_433__55_;
      r_433__54_ <= r_n_433__54_;
      r_433__53_ <= r_n_433__53_;
      r_433__52_ <= r_n_433__52_;
      r_433__51_ <= r_n_433__51_;
      r_433__50_ <= r_n_433__50_;
      r_433__49_ <= r_n_433__49_;
      r_433__48_ <= r_n_433__48_;
      r_433__47_ <= r_n_433__47_;
      r_433__46_ <= r_n_433__46_;
      r_433__45_ <= r_n_433__45_;
      r_433__44_ <= r_n_433__44_;
      r_433__43_ <= r_n_433__43_;
      r_433__42_ <= r_n_433__42_;
      r_433__41_ <= r_n_433__41_;
      r_433__40_ <= r_n_433__40_;
      r_433__39_ <= r_n_433__39_;
      r_433__38_ <= r_n_433__38_;
      r_433__37_ <= r_n_433__37_;
      r_433__36_ <= r_n_433__36_;
      r_433__35_ <= r_n_433__35_;
      r_433__34_ <= r_n_433__34_;
      r_433__33_ <= r_n_433__33_;
      r_433__32_ <= r_n_433__32_;
      r_433__31_ <= r_n_433__31_;
      r_433__30_ <= r_n_433__30_;
      r_433__29_ <= r_n_433__29_;
      r_433__28_ <= r_n_433__28_;
      r_433__27_ <= r_n_433__27_;
      r_433__26_ <= r_n_433__26_;
      r_433__25_ <= r_n_433__25_;
      r_433__24_ <= r_n_433__24_;
      r_433__23_ <= r_n_433__23_;
      r_433__22_ <= r_n_433__22_;
      r_433__21_ <= r_n_433__21_;
      r_433__20_ <= r_n_433__20_;
      r_433__19_ <= r_n_433__19_;
      r_433__18_ <= r_n_433__18_;
      r_433__17_ <= r_n_433__17_;
      r_433__16_ <= r_n_433__16_;
      r_433__15_ <= r_n_433__15_;
      r_433__14_ <= r_n_433__14_;
      r_433__13_ <= r_n_433__13_;
      r_433__12_ <= r_n_433__12_;
      r_433__11_ <= r_n_433__11_;
      r_433__10_ <= r_n_433__10_;
      r_433__9_ <= r_n_433__9_;
      r_433__8_ <= r_n_433__8_;
      r_433__7_ <= r_n_433__7_;
      r_433__6_ <= r_n_433__6_;
      r_433__5_ <= r_n_433__5_;
      r_433__4_ <= r_n_433__4_;
      r_433__3_ <= r_n_433__3_;
      r_433__2_ <= r_n_433__2_;
      r_433__1_ <= r_n_433__1_;
      r_433__0_ <= r_n_433__0_;
    end 
    if(N4018) begin
      r_434__63_ <= r_n_434__63_;
      r_434__62_ <= r_n_434__62_;
      r_434__61_ <= r_n_434__61_;
      r_434__60_ <= r_n_434__60_;
      r_434__59_ <= r_n_434__59_;
      r_434__58_ <= r_n_434__58_;
      r_434__57_ <= r_n_434__57_;
      r_434__56_ <= r_n_434__56_;
      r_434__55_ <= r_n_434__55_;
      r_434__54_ <= r_n_434__54_;
      r_434__53_ <= r_n_434__53_;
      r_434__52_ <= r_n_434__52_;
      r_434__51_ <= r_n_434__51_;
      r_434__50_ <= r_n_434__50_;
      r_434__49_ <= r_n_434__49_;
      r_434__48_ <= r_n_434__48_;
      r_434__47_ <= r_n_434__47_;
      r_434__46_ <= r_n_434__46_;
      r_434__45_ <= r_n_434__45_;
      r_434__44_ <= r_n_434__44_;
      r_434__43_ <= r_n_434__43_;
      r_434__42_ <= r_n_434__42_;
      r_434__41_ <= r_n_434__41_;
      r_434__40_ <= r_n_434__40_;
      r_434__39_ <= r_n_434__39_;
      r_434__38_ <= r_n_434__38_;
      r_434__37_ <= r_n_434__37_;
      r_434__36_ <= r_n_434__36_;
      r_434__35_ <= r_n_434__35_;
      r_434__34_ <= r_n_434__34_;
      r_434__33_ <= r_n_434__33_;
      r_434__32_ <= r_n_434__32_;
      r_434__31_ <= r_n_434__31_;
      r_434__30_ <= r_n_434__30_;
      r_434__29_ <= r_n_434__29_;
      r_434__28_ <= r_n_434__28_;
      r_434__27_ <= r_n_434__27_;
      r_434__26_ <= r_n_434__26_;
      r_434__25_ <= r_n_434__25_;
      r_434__24_ <= r_n_434__24_;
      r_434__23_ <= r_n_434__23_;
      r_434__22_ <= r_n_434__22_;
      r_434__21_ <= r_n_434__21_;
      r_434__20_ <= r_n_434__20_;
      r_434__19_ <= r_n_434__19_;
      r_434__18_ <= r_n_434__18_;
      r_434__17_ <= r_n_434__17_;
      r_434__16_ <= r_n_434__16_;
      r_434__15_ <= r_n_434__15_;
      r_434__14_ <= r_n_434__14_;
      r_434__13_ <= r_n_434__13_;
      r_434__12_ <= r_n_434__12_;
      r_434__11_ <= r_n_434__11_;
      r_434__10_ <= r_n_434__10_;
      r_434__9_ <= r_n_434__9_;
      r_434__8_ <= r_n_434__8_;
      r_434__7_ <= r_n_434__7_;
      r_434__6_ <= r_n_434__6_;
      r_434__5_ <= r_n_434__5_;
      r_434__4_ <= r_n_434__4_;
      r_434__3_ <= r_n_434__3_;
      r_434__2_ <= r_n_434__2_;
      r_434__1_ <= r_n_434__1_;
      r_434__0_ <= r_n_434__0_;
    end 
    if(N4019) begin
      r_435__63_ <= r_n_435__63_;
      r_435__62_ <= r_n_435__62_;
      r_435__61_ <= r_n_435__61_;
      r_435__60_ <= r_n_435__60_;
      r_435__59_ <= r_n_435__59_;
      r_435__58_ <= r_n_435__58_;
      r_435__57_ <= r_n_435__57_;
      r_435__56_ <= r_n_435__56_;
      r_435__55_ <= r_n_435__55_;
      r_435__54_ <= r_n_435__54_;
      r_435__53_ <= r_n_435__53_;
      r_435__52_ <= r_n_435__52_;
      r_435__51_ <= r_n_435__51_;
      r_435__50_ <= r_n_435__50_;
      r_435__49_ <= r_n_435__49_;
      r_435__48_ <= r_n_435__48_;
      r_435__47_ <= r_n_435__47_;
      r_435__46_ <= r_n_435__46_;
      r_435__45_ <= r_n_435__45_;
      r_435__44_ <= r_n_435__44_;
      r_435__43_ <= r_n_435__43_;
      r_435__42_ <= r_n_435__42_;
      r_435__41_ <= r_n_435__41_;
      r_435__40_ <= r_n_435__40_;
      r_435__39_ <= r_n_435__39_;
      r_435__38_ <= r_n_435__38_;
      r_435__37_ <= r_n_435__37_;
      r_435__36_ <= r_n_435__36_;
      r_435__35_ <= r_n_435__35_;
      r_435__34_ <= r_n_435__34_;
      r_435__33_ <= r_n_435__33_;
      r_435__32_ <= r_n_435__32_;
      r_435__31_ <= r_n_435__31_;
      r_435__30_ <= r_n_435__30_;
      r_435__29_ <= r_n_435__29_;
      r_435__28_ <= r_n_435__28_;
      r_435__27_ <= r_n_435__27_;
      r_435__26_ <= r_n_435__26_;
      r_435__25_ <= r_n_435__25_;
      r_435__24_ <= r_n_435__24_;
      r_435__23_ <= r_n_435__23_;
      r_435__22_ <= r_n_435__22_;
      r_435__21_ <= r_n_435__21_;
      r_435__20_ <= r_n_435__20_;
      r_435__19_ <= r_n_435__19_;
      r_435__18_ <= r_n_435__18_;
      r_435__17_ <= r_n_435__17_;
      r_435__16_ <= r_n_435__16_;
      r_435__15_ <= r_n_435__15_;
      r_435__14_ <= r_n_435__14_;
      r_435__13_ <= r_n_435__13_;
      r_435__12_ <= r_n_435__12_;
      r_435__11_ <= r_n_435__11_;
      r_435__10_ <= r_n_435__10_;
      r_435__9_ <= r_n_435__9_;
      r_435__8_ <= r_n_435__8_;
      r_435__7_ <= r_n_435__7_;
      r_435__6_ <= r_n_435__6_;
      r_435__5_ <= r_n_435__5_;
      r_435__4_ <= r_n_435__4_;
      r_435__3_ <= r_n_435__3_;
      r_435__2_ <= r_n_435__2_;
      r_435__1_ <= r_n_435__1_;
      r_435__0_ <= r_n_435__0_;
    end 
    if(N4020) begin
      r_436__63_ <= r_n_436__63_;
      r_436__62_ <= r_n_436__62_;
      r_436__61_ <= r_n_436__61_;
      r_436__60_ <= r_n_436__60_;
      r_436__59_ <= r_n_436__59_;
      r_436__58_ <= r_n_436__58_;
      r_436__57_ <= r_n_436__57_;
      r_436__56_ <= r_n_436__56_;
      r_436__55_ <= r_n_436__55_;
      r_436__54_ <= r_n_436__54_;
      r_436__53_ <= r_n_436__53_;
      r_436__52_ <= r_n_436__52_;
      r_436__51_ <= r_n_436__51_;
      r_436__50_ <= r_n_436__50_;
      r_436__49_ <= r_n_436__49_;
      r_436__48_ <= r_n_436__48_;
      r_436__47_ <= r_n_436__47_;
      r_436__46_ <= r_n_436__46_;
      r_436__45_ <= r_n_436__45_;
      r_436__44_ <= r_n_436__44_;
      r_436__43_ <= r_n_436__43_;
      r_436__42_ <= r_n_436__42_;
      r_436__41_ <= r_n_436__41_;
      r_436__40_ <= r_n_436__40_;
      r_436__39_ <= r_n_436__39_;
      r_436__38_ <= r_n_436__38_;
      r_436__37_ <= r_n_436__37_;
      r_436__36_ <= r_n_436__36_;
      r_436__35_ <= r_n_436__35_;
      r_436__34_ <= r_n_436__34_;
      r_436__33_ <= r_n_436__33_;
      r_436__32_ <= r_n_436__32_;
      r_436__31_ <= r_n_436__31_;
      r_436__30_ <= r_n_436__30_;
      r_436__29_ <= r_n_436__29_;
      r_436__28_ <= r_n_436__28_;
      r_436__27_ <= r_n_436__27_;
      r_436__26_ <= r_n_436__26_;
      r_436__25_ <= r_n_436__25_;
      r_436__24_ <= r_n_436__24_;
      r_436__23_ <= r_n_436__23_;
      r_436__22_ <= r_n_436__22_;
      r_436__21_ <= r_n_436__21_;
      r_436__20_ <= r_n_436__20_;
      r_436__19_ <= r_n_436__19_;
      r_436__18_ <= r_n_436__18_;
      r_436__17_ <= r_n_436__17_;
      r_436__16_ <= r_n_436__16_;
      r_436__15_ <= r_n_436__15_;
      r_436__14_ <= r_n_436__14_;
      r_436__13_ <= r_n_436__13_;
      r_436__12_ <= r_n_436__12_;
      r_436__11_ <= r_n_436__11_;
      r_436__10_ <= r_n_436__10_;
      r_436__9_ <= r_n_436__9_;
      r_436__8_ <= r_n_436__8_;
      r_436__7_ <= r_n_436__7_;
      r_436__6_ <= r_n_436__6_;
      r_436__5_ <= r_n_436__5_;
      r_436__4_ <= r_n_436__4_;
      r_436__3_ <= r_n_436__3_;
      r_436__2_ <= r_n_436__2_;
      r_436__1_ <= r_n_436__1_;
      r_436__0_ <= r_n_436__0_;
    end 
    if(N4021) begin
      r_437__63_ <= r_n_437__63_;
      r_437__62_ <= r_n_437__62_;
      r_437__61_ <= r_n_437__61_;
      r_437__60_ <= r_n_437__60_;
      r_437__59_ <= r_n_437__59_;
      r_437__58_ <= r_n_437__58_;
      r_437__57_ <= r_n_437__57_;
      r_437__56_ <= r_n_437__56_;
      r_437__55_ <= r_n_437__55_;
      r_437__54_ <= r_n_437__54_;
      r_437__53_ <= r_n_437__53_;
      r_437__52_ <= r_n_437__52_;
      r_437__51_ <= r_n_437__51_;
      r_437__50_ <= r_n_437__50_;
      r_437__49_ <= r_n_437__49_;
      r_437__48_ <= r_n_437__48_;
      r_437__47_ <= r_n_437__47_;
      r_437__46_ <= r_n_437__46_;
      r_437__45_ <= r_n_437__45_;
      r_437__44_ <= r_n_437__44_;
      r_437__43_ <= r_n_437__43_;
      r_437__42_ <= r_n_437__42_;
      r_437__41_ <= r_n_437__41_;
      r_437__40_ <= r_n_437__40_;
      r_437__39_ <= r_n_437__39_;
      r_437__38_ <= r_n_437__38_;
      r_437__37_ <= r_n_437__37_;
      r_437__36_ <= r_n_437__36_;
      r_437__35_ <= r_n_437__35_;
      r_437__34_ <= r_n_437__34_;
      r_437__33_ <= r_n_437__33_;
      r_437__32_ <= r_n_437__32_;
      r_437__31_ <= r_n_437__31_;
      r_437__30_ <= r_n_437__30_;
      r_437__29_ <= r_n_437__29_;
      r_437__28_ <= r_n_437__28_;
      r_437__27_ <= r_n_437__27_;
      r_437__26_ <= r_n_437__26_;
      r_437__25_ <= r_n_437__25_;
      r_437__24_ <= r_n_437__24_;
      r_437__23_ <= r_n_437__23_;
      r_437__22_ <= r_n_437__22_;
      r_437__21_ <= r_n_437__21_;
      r_437__20_ <= r_n_437__20_;
      r_437__19_ <= r_n_437__19_;
      r_437__18_ <= r_n_437__18_;
      r_437__17_ <= r_n_437__17_;
      r_437__16_ <= r_n_437__16_;
      r_437__15_ <= r_n_437__15_;
      r_437__14_ <= r_n_437__14_;
      r_437__13_ <= r_n_437__13_;
      r_437__12_ <= r_n_437__12_;
      r_437__11_ <= r_n_437__11_;
      r_437__10_ <= r_n_437__10_;
      r_437__9_ <= r_n_437__9_;
      r_437__8_ <= r_n_437__8_;
      r_437__7_ <= r_n_437__7_;
      r_437__6_ <= r_n_437__6_;
      r_437__5_ <= r_n_437__5_;
      r_437__4_ <= r_n_437__4_;
      r_437__3_ <= r_n_437__3_;
      r_437__2_ <= r_n_437__2_;
      r_437__1_ <= r_n_437__1_;
      r_437__0_ <= r_n_437__0_;
    end 
    if(N4022) begin
      r_438__63_ <= r_n_438__63_;
      r_438__62_ <= r_n_438__62_;
      r_438__61_ <= r_n_438__61_;
      r_438__60_ <= r_n_438__60_;
      r_438__59_ <= r_n_438__59_;
      r_438__58_ <= r_n_438__58_;
      r_438__57_ <= r_n_438__57_;
      r_438__56_ <= r_n_438__56_;
      r_438__55_ <= r_n_438__55_;
      r_438__54_ <= r_n_438__54_;
      r_438__53_ <= r_n_438__53_;
      r_438__52_ <= r_n_438__52_;
      r_438__51_ <= r_n_438__51_;
      r_438__50_ <= r_n_438__50_;
      r_438__49_ <= r_n_438__49_;
      r_438__48_ <= r_n_438__48_;
      r_438__47_ <= r_n_438__47_;
      r_438__46_ <= r_n_438__46_;
      r_438__45_ <= r_n_438__45_;
      r_438__44_ <= r_n_438__44_;
      r_438__43_ <= r_n_438__43_;
      r_438__42_ <= r_n_438__42_;
      r_438__41_ <= r_n_438__41_;
      r_438__40_ <= r_n_438__40_;
      r_438__39_ <= r_n_438__39_;
      r_438__38_ <= r_n_438__38_;
      r_438__37_ <= r_n_438__37_;
      r_438__36_ <= r_n_438__36_;
      r_438__35_ <= r_n_438__35_;
      r_438__34_ <= r_n_438__34_;
      r_438__33_ <= r_n_438__33_;
      r_438__32_ <= r_n_438__32_;
      r_438__31_ <= r_n_438__31_;
      r_438__30_ <= r_n_438__30_;
      r_438__29_ <= r_n_438__29_;
      r_438__28_ <= r_n_438__28_;
      r_438__27_ <= r_n_438__27_;
      r_438__26_ <= r_n_438__26_;
      r_438__25_ <= r_n_438__25_;
      r_438__24_ <= r_n_438__24_;
      r_438__23_ <= r_n_438__23_;
      r_438__22_ <= r_n_438__22_;
      r_438__21_ <= r_n_438__21_;
      r_438__20_ <= r_n_438__20_;
      r_438__19_ <= r_n_438__19_;
      r_438__18_ <= r_n_438__18_;
      r_438__17_ <= r_n_438__17_;
      r_438__16_ <= r_n_438__16_;
      r_438__15_ <= r_n_438__15_;
      r_438__14_ <= r_n_438__14_;
      r_438__13_ <= r_n_438__13_;
      r_438__12_ <= r_n_438__12_;
      r_438__11_ <= r_n_438__11_;
      r_438__10_ <= r_n_438__10_;
      r_438__9_ <= r_n_438__9_;
      r_438__8_ <= r_n_438__8_;
      r_438__7_ <= r_n_438__7_;
      r_438__6_ <= r_n_438__6_;
      r_438__5_ <= r_n_438__5_;
      r_438__4_ <= r_n_438__4_;
      r_438__3_ <= r_n_438__3_;
      r_438__2_ <= r_n_438__2_;
      r_438__1_ <= r_n_438__1_;
      r_438__0_ <= r_n_438__0_;
    end 
    if(N4023) begin
      r_439__63_ <= r_n_439__63_;
      r_439__62_ <= r_n_439__62_;
      r_439__61_ <= r_n_439__61_;
      r_439__60_ <= r_n_439__60_;
      r_439__59_ <= r_n_439__59_;
      r_439__58_ <= r_n_439__58_;
      r_439__57_ <= r_n_439__57_;
      r_439__56_ <= r_n_439__56_;
      r_439__55_ <= r_n_439__55_;
      r_439__54_ <= r_n_439__54_;
      r_439__53_ <= r_n_439__53_;
      r_439__52_ <= r_n_439__52_;
      r_439__51_ <= r_n_439__51_;
      r_439__50_ <= r_n_439__50_;
      r_439__49_ <= r_n_439__49_;
      r_439__48_ <= r_n_439__48_;
      r_439__47_ <= r_n_439__47_;
      r_439__46_ <= r_n_439__46_;
      r_439__45_ <= r_n_439__45_;
      r_439__44_ <= r_n_439__44_;
      r_439__43_ <= r_n_439__43_;
      r_439__42_ <= r_n_439__42_;
      r_439__41_ <= r_n_439__41_;
      r_439__40_ <= r_n_439__40_;
      r_439__39_ <= r_n_439__39_;
      r_439__38_ <= r_n_439__38_;
      r_439__37_ <= r_n_439__37_;
      r_439__36_ <= r_n_439__36_;
      r_439__35_ <= r_n_439__35_;
      r_439__34_ <= r_n_439__34_;
      r_439__33_ <= r_n_439__33_;
      r_439__32_ <= r_n_439__32_;
      r_439__31_ <= r_n_439__31_;
      r_439__30_ <= r_n_439__30_;
      r_439__29_ <= r_n_439__29_;
      r_439__28_ <= r_n_439__28_;
      r_439__27_ <= r_n_439__27_;
      r_439__26_ <= r_n_439__26_;
      r_439__25_ <= r_n_439__25_;
      r_439__24_ <= r_n_439__24_;
      r_439__23_ <= r_n_439__23_;
      r_439__22_ <= r_n_439__22_;
      r_439__21_ <= r_n_439__21_;
      r_439__20_ <= r_n_439__20_;
      r_439__19_ <= r_n_439__19_;
      r_439__18_ <= r_n_439__18_;
      r_439__17_ <= r_n_439__17_;
      r_439__16_ <= r_n_439__16_;
      r_439__15_ <= r_n_439__15_;
      r_439__14_ <= r_n_439__14_;
      r_439__13_ <= r_n_439__13_;
      r_439__12_ <= r_n_439__12_;
      r_439__11_ <= r_n_439__11_;
      r_439__10_ <= r_n_439__10_;
      r_439__9_ <= r_n_439__9_;
      r_439__8_ <= r_n_439__8_;
      r_439__7_ <= r_n_439__7_;
      r_439__6_ <= r_n_439__6_;
      r_439__5_ <= r_n_439__5_;
      r_439__4_ <= r_n_439__4_;
      r_439__3_ <= r_n_439__3_;
      r_439__2_ <= r_n_439__2_;
      r_439__1_ <= r_n_439__1_;
      r_439__0_ <= r_n_439__0_;
    end 
    if(N4024) begin
      r_440__63_ <= r_n_440__63_;
      r_440__62_ <= r_n_440__62_;
      r_440__61_ <= r_n_440__61_;
      r_440__60_ <= r_n_440__60_;
      r_440__59_ <= r_n_440__59_;
      r_440__58_ <= r_n_440__58_;
      r_440__57_ <= r_n_440__57_;
      r_440__56_ <= r_n_440__56_;
      r_440__55_ <= r_n_440__55_;
      r_440__54_ <= r_n_440__54_;
      r_440__53_ <= r_n_440__53_;
      r_440__52_ <= r_n_440__52_;
      r_440__51_ <= r_n_440__51_;
      r_440__50_ <= r_n_440__50_;
      r_440__49_ <= r_n_440__49_;
      r_440__48_ <= r_n_440__48_;
      r_440__47_ <= r_n_440__47_;
      r_440__46_ <= r_n_440__46_;
      r_440__45_ <= r_n_440__45_;
      r_440__44_ <= r_n_440__44_;
      r_440__43_ <= r_n_440__43_;
      r_440__42_ <= r_n_440__42_;
      r_440__41_ <= r_n_440__41_;
      r_440__40_ <= r_n_440__40_;
      r_440__39_ <= r_n_440__39_;
      r_440__38_ <= r_n_440__38_;
      r_440__37_ <= r_n_440__37_;
      r_440__36_ <= r_n_440__36_;
      r_440__35_ <= r_n_440__35_;
      r_440__34_ <= r_n_440__34_;
      r_440__33_ <= r_n_440__33_;
      r_440__32_ <= r_n_440__32_;
      r_440__31_ <= r_n_440__31_;
      r_440__30_ <= r_n_440__30_;
      r_440__29_ <= r_n_440__29_;
      r_440__28_ <= r_n_440__28_;
      r_440__27_ <= r_n_440__27_;
      r_440__26_ <= r_n_440__26_;
      r_440__25_ <= r_n_440__25_;
      r_440__24_ <= r_n_440__24_;
      r_440__23_ <= r_n_440__23_;
      r_440__22_ <= r_n_440__22_;
      r_440__21_ <= r_n_440__21_;
      r_440__20_ <= r_n_440__20_;
      r_440__19_ <= r_n_440__19_;
      r_440__18_ <= r_n_440__18_;
      r_440__17_ <= r_n_440__17_;
      r_440__16_ <= r_n_440__16_;
      r_440__15_ <= r_n_440__15_;
      r_440__14_ <= r_n_440__14_;
      r_440__13_ <= r_n_440__13_;
      r_440__12_ <= r_n_440__12_;
      r_440__11_ <= r_n_440__11_;
      r_440__10_ <= r_n_440__10_;
      r_440__9_ <= r_n_440__9_;
      r_440__8_ <= r_n_440__8_;
      r_440__7_ <= r_n_440__7_;
      r_440__6_ <= r_n_440__6_;
      r_440__5_ <= r_n_440__5_;
      r_440__4_ <= r_n_440__4_;
      r_440__3_ <= r_n_440__3_;
      r_440__2_ <= r_n_440__2_;
      r_440__1_ <= r_n_440__1_;
      r_440__0_ <= r_n_440__0_;
    end 
    if(N4025) begin
      r_441__63_ <= r_n_441__63_;
      r_441__62_ <= r_n_441__62_;
      r_441__61_ <= r_n_441__61_;
      r_441__60_ <= r_n_441__60_;
      r_441__59_ <= r_n_441__59_;
      r_441__58_ <= r_n_441__58_;
      r_441__57_ <= r_n_441__57_;
      r_441__56_ <= r_n_441__56_;
      r_441__55_ <= r_n_441__55_;
      r_441__54_ <= r_n_441__54_;
      r_441__53_ <= r_n_441__53_;
      r_441__52_ <= r_n_441__52_;
      r_441__51_ <= r_n_441__51_;
      r_441__50_ <= r_n_441__50_;
      r_441__49_ <= r_n_441__49_;
      r_441__48_ <= r_n_441__48_;
      r_441__47_ <= r_n_441__47_;
      r_441__46_ <= r_n_441__46_;
      r_441__45_ <= r_n_441__45_;
      r_441__44_ <= r_n_441__44_;
      r_441__43_ <= r_n_441__43_;
      r_441__42_ <= r_n_441__42_;
      r_441__41_ <= r_n_441__41_;
      r_441__40_ <= r_n_441__40_;
      r_441__39_ <= r_n_441__39_;
      r_441__38_ <= r_n_441__38_;
      r_441__37_ <= r_n_441__37_;
      r_441__36_ <= r_n_441__36_;
      r_441__35_ <= r_n_441__35_;
      r_441__34_ <= r_n_441__34_;
      r_441__33_ <= r_n_441__33_;
      r_441__32_ <= r_n_441__32_;
      r_441__31_ <= r_n_441__31_;
      r_441__30_ <= r_n_441__30_;
      r_441__29_ <= r_n_441__29_;
      r_441__28_ <= r_n_441__28_;
      r_441__27_ <= r_n_441__27_;
      r_441__26_ <= r_n_441__26_;
      r_441__25_ <= r_n_441__25_;
      r_441__24_ <= r_n_441__24_;
      r_441__23_ <= r_n_441__23_;
      r_441__22_ <= r_n_441__22_;
      r_441__21_ <= r_n_441__21_;
      r_441__20_ <= r_n_441__20_;
      r_441__19_ <= r_n_441__19_;
      r_441__18_ <= r_n_441__18_;
      r_441__17_ <= r_n_441__17_;
      r_441__16_ <= r_n_441__16_;
      r_441__15_ <= r_n_441__15_;
      r_441__14_ <= r_n_441__14_;
      r_441__13_ <= r_n_441__13_;
      r_441__12_ <= r_n_441__12_;
      r_441__11_ <= r_n_441__11_;
      r_441__10_ <= r_n_441__10_;
      r_441__9_ <= r_n_441__9_;
      r_441__8_ <= r_n_441__8_;
      r_441__7_ <= r_n_441__7_;
      r_441__6_ <= r_n_441__6_;
      r_441__5_ <= r_n_441__5_;
      r_441__4_ <= r_n_441__4_;
      r_441__3_ <= r_n_441__3_;
      r_441__2_ <= r_n_441__2_;
      r_441__1_ <= r_n_441__1_;
      r_441__0_ <= r_n_441__0_;
    end 
    if(N4026) begin
      r_442__63_ <= r_n_442__63_;
      r_442__62_ <= r_n_442__62_;
      r_442__61_ <= r_n_442__61_;
      r_442__60_ <= r_n_442__60_;
      r_442__59_ <= r_n_442__59_;
      r_442__58_ <= r_n_442__58_;
      r_442__57_ <= r_n_442__57_;
      r_442__56_ <= r_n_442__56_;
      r_442__55_ <= r_n_442__55_;
      r_442__54_ <= r_n_442__54_;
      r_442__53_ <= r_n_442__53_;
      r_442__52_ <= r_n_442__52_;
      r_442__51_ <= r_n_442__51_;
      r_442__50_ <= r_n_442__50_;
      r_442__49_ <= r_n_442__49_;
      r_442__48_ <= r_n_442__48_;
      r_442__47_ <= r_n_442__47_;
      r_442__46_ <= r_n_442__46_;
      r_442__45_ <= r_n_442__45_;
      r_442__44_ <= r_n_442__44_;
      r_442__43_ <= r_n_442__43_;
      r_442__42_ <= r_n_442__42_;
      r_442__41_ <= r_n_442__41_;
      r_442__40_ <= r_n_442__40_;
      r_442__39_ <= r_n_442__39_;
      r_442__38_ <= r_n_442__38_;
      r_442__37_ <= r_n_442__37_;
      r_442__36_ <= r_n_442__36_;
      r_442__35_ <= r_n_442__35_;
      r_442__34_ <= r_n_442__34_;
      r_442__33_ <= r_n_442__33_;
      r_442__32_ <= r_n_442__32_;
      r_442__31_ <= r_n_442__31_;
      r_442__30_ <= r_n_442__30_;
      r_442__29_ <= r_n_442__29_;
      r_442__28_ <= r_n_442__28_;
      r_442__27_ <= r_n_442__27_;
      r_442__26_ <= r_n_442__26_;
      r_442__25_ <= r_n_442__25_;
      r_442__24_ <= r_n_442__24_;
      r_442__23_ <= r_n_442__23_;
      r_442__22_ <= r_n_442__22_;
      r_442__21_ <= r_n_442__21_;
      r_442__20_ <= r_n_442__20_;
      r_442__19_ <= r_n_442__19_;
      r_442__18_ <= r_n_442__18_;
      r_442__17_ <= r_n_442__17_;
      r_442__16_ <= r_n_442__16_;
      r_442__15_ <= r_n_442__15_;
      r_442__14_ <= r_n_442__14_;
      r_442__13_ <= r_n_442__13_;
      r_442__12_ <= r_n_442__12_;
      r_442__11_ <= r_n_442__11_;
      r_442__10_ <= r_n_442__10_;
      r_442__9_ <= r_n_442__9_;
      r_442__8_ <= r_n_442__8_;
      r_442__7_ <= r_n_442__7_;
      r_442__6_ <= r_n_442__6_;
      r_442__5_ <= r_n_442__5_;
      r_442__4_ <= r_n_442__4_;
      r_442__3_ <= r_n_442__3_;
      r_442__2_ <= r_n_442__2_;
      r_442__1_ <= r_n_442__1_;
      r_442__0_ <= r_n_442__0_;
    end 
    if(N4027) begin
      r_443__63_ <= r_n_443__63_;
      r_443__62_ <= r_n_443__62_;
      r_443__61_ <= r_n_443__61_;
      r_443__60_ <= r_n_443__60_;
      r_443__59_ <= r_n_443__59_;
      r_443__58_ <= r_n_443__58_;
      r_443__57_ <= r_n_443__57_;
      r_443__56_ <= r_n_443__56_;
      r_443__55_ <= r_n_443__55_;
      r_443__54_ <= r_n_443__54_;
      r_443__53_ <= r_n_443__53_;
      r_443__52_ <= r_n_443__52_;
      r_443__51_ <= r_n_443__51_;
      r_443__50_ <= r_n_443__50_;
      r_443__49_ <= r_n_443__49_;
      r_443__48_ <= r_n_443__48_;
      r_443__47_ <= r_n_443__47_;
      r_443__46_ <= r_n_443__46_;
      r_443__45_ <= r_n_443__45_;
      r_443__44_ <= r_n_443__44_;
      r_443__43_ <= r_n_443__43_;
      r_443__42_ <= r_n_443__42_;
      r_443__41_ <= r_n_443__41_;
      r_443__40_ <= r_n_443__40_;
      r_443__39_ <= r_n_443__39_;
      r_443__38_ <= r_n_443__38_;
      r_443__37_ <= r_n_443__37_;
      r_443__36_ <= r_n_443__36_;
      r_443__35_ <= r_n_443__35_;
      r_443__34_ <= r_n_443__34_;
      r_443__33_ <= r_n_443__33_;
      r_443__32_ <= r_n_443__32_;
      r_443__31_ <= r_n_443__31_;
      r_443__30_ <= r_n_443__30_;
      r_443__29_ <= r_n_443__29_;
      r_443__28_ <= r_n_443__28_;
      r_443__27_ <= r_n_443__27_;
      r_443__26_ <= r_n_443__26_;
      r_443__25_ <= r_n_443__25_;
      r_443__24_ <= r_n_443__24_;
      r_443__23_ <= r_n_443__23_;
      r_443__22_ <= r_n_443__22_;
      r_443__21_ <= r_n_443__21_;
      r_443__20_ <= r_n_443__20_;
      r_443__19_ <= r_n_443__19_;
      r_443__18_ <= r_n_443__18_;
      r_443__17_ <= r_n_443__17_;
      r_443__16_ <= r_n_443__16_;
      r_443__15_ <= r_n_443__15_;
      r_443__14_ <= r_n_443__14_;
      r_443__13_ <= r_n_443__13_;
      r_443__12_ <= r_n_443__12_;
      r_443__11_ <= r_n_443__11_;
      r_443__10_ <= r_n_443__10_;
      r_443__9_ <= r_n_443__9_;
      r_443__8_ <= r_n_443__8_;
      r_443__7_ <= r_n_443__7_;
      r_443__6_ <= r_n_443__6_;
      r_443__5_ <= r_n_443__5_;
      r_443__4_ <= r_n_443__4_;
      r_443__3_ <= r_n_443__3_;
      r_443__2_ <= r_n_443__2_;
      r_443__1_ <= r_n_443__1_;
      r_443__0_ <= r_n_443__0_;
    end 
    if(N4028) begin
      r_444__63_ <= r_n_444__63_;
      r_444__62_ <= r_n_444__62_;
      r_444__61_ <= r_n_444__61_;
      r_444__60_ <= r_n_444__60_;
      r_444__59_ <= r_n_444__59_;
      r_444__58_ <= r_n_444__58_;
      r_444__57_ <= r_n_444__57_;
      r_444__56_ <= r_n_444__56_;
      r_444__55_ <= r_n_444__55_;
      r_444__54_ <= r_n_444__54_;
      r_444__53_ <= r_n_444__53_;
      r_444__52_ <= r_n_444__52_;
      r_444__51_ <= r_n_444__51_;
      r_444__50_ <= r_n_444__50_;
      r_444__49_ <= r_n_444__49_;
      r_444__48_ <= r_n_444__48_;
      r_444__47_ <= r_n_444__47_;
      r_444__46_ <= r_n_444__46_;
      r_444__45_ <= r_n_444__45_;
      r_444__44_ <= r_n_444__44_;
      r_444__43_ <= r_n_444__43_;
      r_444__42_ <= r_n_444__42_;
      r_444__41_ <= r_n_444__41_;
      r_444__40_ <= r_n_444__40_;
      r_444__39_ <= r_n_444__39_;
      r_444__38_ <= r_n_444__38_;
      r_444__37_ <= r_n_444__37_;
      r_444__36_ <= r_n_444__36_;
      r_444__35_ <= r_n_444__35_;
      r_444__34_ <= r_n_444__34_;
      r_444__33_ <= r_n_444__33_;
      r_444__32_ <= r_n_444__32_;
      r_444__31_ <= r_n_444__31_;
      r_444__30_ <= r_n_444__30_;
      r_444__29_ <= r_n_444__29_;
      r_444__28_ <= r_n_444__28_;
      r_444__27_ <= r_n_444__27_;
      r_444__26_ <= r_n_444__26_;
      r_444__25_ <= r_n_444__25_;
      r_444__24_ <= r_n_444__24_;
      r_444__23_ <= r_n_444__23_;
      r_444__22_ <= r_n_444__22_;
      r_444__21_ <= r_n_444__21_;
      r_444__20_ <= r_n_444__20_;
      r_444__19_ <= r_n_444__19_;
      r_444__18_ <= r_n_444__18_;
      r_444__17_ <= r_n_444__17_;
      r_444__16_ <= r_n_444__16_;
      r_444__15_ <= r_n_444__15_;
      r_444__14_ <= r_n_444__14_;
      r_444__13_ <= r_n_444__13_;
      r_444__12_ <= r_n_444__12_;
      r_444__11_ <= r_n_444__11_;
      r_444__10_ <= r_n_444__10_;
      r_444__9_ <= r_n_444__9_;
      r_444__8_ <= r_n_444__8_;
      r_444__7_ <= r_n_444__7_;
      r_444__6_ <= r_n_444__6_;
      r_444__5_ <= r_n_444__5_;
      r_444__4_ <= r_n_444__4_;
      r_444__3_ <= r_n_444__3_;
      r_444__2_ <= r_n_444__2_;
      r_444__1_ <= r_n_444__1_;
      r_444__0_ <= r_n_444__0_;
    end 
    if(N4029) begin
      r_445__63_ <= r_n_445__63_;
      r_445__62_ <= r_n_445__62_;
      r_445__61_ <= r_n_445__61_;
      r_445__60_ <= r_n_445__60_;
      r_445__59_ <= r_n_445__59_;
      r_445__58_ <= r_n_445__58_;
      r_445__57_ <= r_n_445__57_;
      r_445__56_ <= r_n_445__56_;
      r_445__55_ <= r_n_445__55_;
      r_445__54_ <= r_n_445__54_;
      r_445__53_ <= r_n_445__53_;
      r_445__52_ <= r_n_445__52_;
      r_445__51_ <= r_n_445__51_;
      r_445__50_ <= r_n_445__50_;
      r_445__49_ <= r_n_445__49_;
      r_445__48_ <= r_n_445__48_;
      r_445__47_ <= r_n_445__47_;
      r_445__46_ <= r_n_445__46_;
      r_445__45_ <= r_n_445__45_;
      r_445__44_ <= r_n_445__44_;
      r_445__43_ <= r_n_445__43_;
      r_445__42_ <= r_n_445__42_;
      r_445__41_ <= r_n_445__41_;
      r_445__40_ <= r_n_445__40_;
      r_445__39_ <= r_n_445__39_;
      r_445__38_ <= r_n_445__38_;
      r_445__37_ <= r_n_445__37_;
      r_445__36_ <= r_n_445__36_;
      r_445__35_ <= r_n_445__35_;
      r_445__34_ <= r_n_445__34_;
      r_445__33_ <= r_n_445__33_;
      r_445__32_ <= r_n_445__32_;
      r_445__31_ <= r_n_445__31_;
      r_445__30_ <= r_n_445__30_;
      r_445__29_ <= r_n_445__29_;
      r_445__28_ <= r_n_445__28_;
      r_445__27_ <= r_n_445__27_;
      r_445__26_ <= r_n_445__26_;
      r_445__25_ <= r_n_445__25_;
      r_445__24_ <= r_n_445__24_;
      r_445__23_ <= r_n_445__23_;
      r_445__22_ <= r_n_445__22_;
      r_445__21_ <= r_n_445__21_;
      r_445__20_ <= r_n_445__20_;
      r_445__19_ <= r_n_445__19_;
      r_445__18_ <= r_n_445__18_;
      r_445__17_ <= r_n_445__17_;
      r_445__16_ <= r_n_445__16_;
      r_445__15_ <= r_n_445__15_;
      r_445__14_ <= r_n_445__14_;
      r_445__13_ <= r_n_445__13_;
      r_445__12_ <= r_n_445__12_;
      r_445__11_ <= r_n_445__11_;
      r_445__10_ <= r_n_445__10_;
      r_445__9_ <= r_n_445__9_;
      r_445__8_ <= r_n_445__8_;
      r_445__7_ <= r_n_445__7_;
      r_445__6_ <= r_n_445__6_;
      r_445__5_ <= r_n_445__5_;
      r_445__4_ <= r_n_445__4_;
      r_445__3_ <= r_n_445__3_;
      r_445__2_ <= r_n_445__2_;
      r_445__1_ <= r_n_445__1_;
      r_445__0_ <= r_n_445__0_;
    end 
    if(N4030) begin
      r_446__63_ <= r_n_446__63_;
      r_446__62_ <= r_n_446__62_;
      r_446__61_ <= r_n_446__61_;
      r_446__60_ <= r_n_446__60_;
      r_446__59_ <= r_n_446__59_;
      r_446__58_ <= r_n_446__58_;
      r_446__57_ <= r_n_446__57_;
      r_446__56_ <= r_n_446__56_;
      r_446__55_ <= r_n_446__55_;
      r_446__54_ <= r_n_446__54_;
      r_446__53_ <= r_n_446__53_;
      r_446__52_ <= r_n_446__52_;
      r_446__51_ <= r_n_446__51_;
      r_446__50_ <= r_n_446__50_;
      r_446__49_ <= r_n_446__49_;
      r_446__48_ <= r_n_446__48_;
      r_446__47_ <= r_n_446__47_;
      r_446__46_ <= r_n_446__46_;
      r_446__45_ <= r_n_446__45_;
      r_446__44_ <= r_n_446__44_;
      r_446__43_ <= r_n_446__43_;
      r_446__42_ <= r_n_446__42_;
      r_446__41_ <= r_n_446__41_;
      r_446__40_ <= r_n_446__40_;
      r_446__39_ <= r_n_446__39_;
      r_446__38_ <= r_n_446__38_;
      r_446__37_ <= r_n_446__37_;
      r_446__36_ <= r_n_446__36_;
      r_446__35_ <= r_n_446__35_;
      r_446__34_ <= r_n_446__34_;
      r_446__33_ <= r_n_446__33_;
      r_446__32_ <= r_n_446__32_;
      r_446__31_ <= r_n_446__31_;
      r_446__30_ <= r_n_446__30_;
      r_446__29_ <= r_n_446__29_;
      r_446__28_ <= r_n_446__28_;
      r_446__27_ <= r_n_446__27_;
      r_446__26_ <= r_n_446__26_;
      r_446__25_ <= r_n_446__25_;
      r_446__24_ <= r_n_446__24_;
      r_446__23_ <= r_n_446__23_;
      r_446__22_ <= r_n_446__22_;
      r_446__21_ <= r_n_446__21_;
      r_446__20_ <= r_n_446__20_;
      r_446__19_ <= r_n_446__19_;
      r_446__18_ <= r_n_446__18_;
      r_446__17_ <= r_n_446__17_;
      r_446__16_ <= r_n_446__16_;
      r_446__15_ <= r_n_446__15_;
      r_446__14_ <= r_n_446__14_;
      r_446__13_ <= r_n_446__13_;
      r_446__12_ <= r_n_446__12_;
      r_446__11_ <= r_n_446__11_;
      r_446__10_ <= r_n_446__10_;
      r_446__9_ <= r_n_446__9_;
      r_446__8_ <= r_n_446__8_;
      r_446__7_ <= r_n_446__7_;
      r_446__6_ <= r_n_446__6_;
      r_446__5_ <= r_n_446__5_;
      r_446__4_ <= r_n_446__4_;
      r_446__3_ <= r_n_446__3_;
      r_446__2_ <= r_n_446__2_;
      r_446__1_ <= r_n_446__1_;
      r_446__0_ <= r_n_446__0_;
    end 
    if(N4031) begin
      r_447__63_ <= r_n_447__63_;
      r_447__62_ <= r_n_447__62_;
      r_447__61_ <= r_n_447__61_;
      r_447__60_ <= r_n_447__60_;
      r_447__59_ <= r_n_447__59_;
      r_447__58_ <= r_n_447__58_;
      r_447__57_ <= r_n_447__57_;
      r_447__56_ <= r_n_447__56_;
      r_447__55_ <= r_n_447__55_;
      r_447__54_ <= r_n_447__54_;
      r_447__53_ <= r_n_447__53_;
      r_447__52_ <= r_n_447__52_;
      r_447__51_ <= r_n_447__51_;
      r_447__50_ <= r_n_447__50_;
      r_447__49_ <= r_n_447__49_;
      r_447__48_ <= r_n_447__48_;
      r_447__47_ <= r_n_447__47_;
      r_447__46_ <= r_n_447__46_;
      r_447__45_ <= r_n_447__45_;
      r_447__44_ <= r_n_447__44_;
      r_447__43_ <= r_n_447__43_;
      r_447__42_ <= r_n_447__42_;
      r_447__41_ <= r_n_447__41_;
      r_447__40_ <= r_n_447__40_;
      r_447__39_ <= r_n_447__39_;
      r_447__38_ <= r_n_447__38_;
      r_447__37_ <= r_n_447__37_;
      r_447__36_ <= r_n_447__36_;
      r_447__35_ <= r_n_447__35_;
      r_447__34_ <= r_n_447__34_;
      r_447__33_ <= r_n_447__33_;
      r_447__32_ <= r_n_447__32_;
      r_447__31_ <= r_n_447__31_;
      r_447__30_ <= r_n_447__30_;
      r_447__29_ <= r_n_447__29_;
      r_447__28_ <= r_n_447__28_;
      r_447__27_ <= r_n_447__27_;
      r_447__26_ <= r_n_447__26_;
      r_447__25_ <= r_n_447__25_;
      r_447__24_ <= r_n_447__24_;
      r_447__23_ <= r_n_447__23_;
      r_447__22_ <= r_n_447__22_;
      r_447__21_ <= r_n_447__21_;
      r_447__20_ <= r_n_447__20_;
      r_447__19_ <= r_n_447__19_;
      r_447__18_ <= r_n_447__18_;
      r_447__17_ <= r_n_447__17_;
      r_447__16_ <= r_n_447__16_;
      r_447__15_ <= r_n_447__15_;
      r_447__14_ <= r_n_447__14_;
      r_447__13_ <= r_n_447__13_;
      r_447__12_ <= r_n_447__12_;
      r_447__11_ <= r_n_447__11_;
      r_447__10_ <= r_n_447__10_;
      r_447__9_ <= r_n_447__9_;
      r_447__8_ <= r_n_447__8_;
      r_447__7_ <= r_n_447__7_;
      r_447__6_ <= r_n_447__6_;
      r_447__5_ <= r_n_447__5_;
      r_447__4_ <= r_n_447__4_;
      r_447__3_ <= r_n_447__3_;
      r_447__2_ <= r_n_447__2_;
      r_447__1_ <= r_n_447__1_;
      r_447__0_ <= r_n_447__0_;
    end 
    if(N4032) begin
      r_448__63_ <= r_n_448__63_;
      r_448__62_ <= r_n_448__62_;
      r_448__61_ <= r_n_448__61_;
      r_448__60_ <= r_n_448__60_;
      r_448__59_ <= r_n_448__59_;
      r_448__58_ <= r_n_448__58_;
      r_448__57_ <= r_n_448__57_;
      r_448__56_ <= r_n_448__56_;
      r_448__55_ <= r_n_448__55_;
      r_448__54_ <= r_n_448__54_;
      r_448__53_ <= r_n_448__53_;
      r_448__52_ <= r_n_448__52_;
      r_448__51_ <= r_n_448__51_;
      r_448__50_ <= r_n_448__50_;
      r_448__49_ <= r_n_448__49_;
      r_448__48_ <= r_n_448__48_;
      r_448__47_ <= r_n_448__47_;
      r_448__46_ <= r_n_448__46_;
      r_448__45_ <= r_n_448__45_;
      r_448__44_ <= r_n_448__44_;
      r_448__43_ <= r_n_448__43_;
      r_448__42_ <= r_n_448__42_;
      r_448__41_ <= r_n_448__41_;
      r_448__40_ <= r_n_448__40_;
      r_448__39_ <= r_n_448__39_;
      r_448__38_ <= r_n_448__38_;
      r_448__37_ <= r_n_448__37_;
      r_448__36_ <= r_n_448__36_;
      r_448__35_ <= r_n_448__35_;
      r_448__34_ <= r_n_448__34_;
      r_448__33_ <= r_n_448__33_;
      r_448__32_ <= r_n_448__32_;
      r_448__31_ <= r_n_448__31_;
      r_448__30_ <= r_n_448__30_;
      r_448__29_ <= r_n_448__29_;
      r_448__28_ <= r_n_448__28_;
      r_448__27_ <= r_n_448__27_;
      r_448__26_ <= r_n_448__26_;
      r_448__25_ <= r_n_448__25_;
      r_448__24_ <= r_n_448__24_;
      r_448__23_ <= r_n_448__23_;
      r_448__22_ <= r_n_448__22_;
      r_448__21_ <= r_n_448__21_;
      r_448__20_ <= r_n_448__20_;
      r_448__19_ <= r_n_448__19_;
      r_448__18_ <= r_n_448__18_;
      r_448__17_ <= r_n_448__17_;
      r_448__16_ <= r_n_448__16_;
      r_448__15_ <= r_n_448__15_;
      r_448__14_ <= r_n_448__14_;
      r_448__13_ <= r_n_448__13_;
      r_448__12_ <= r_n_448__12_;
      r_448__11_ <= r_n_448__11_;
      r_448__10_ <= r_n_448__10_;
      r_448__9_ <= r_n_448__9_;
      r_448__8_ <= r_n_448__8_;
      r_448__7_ <= r_n_448__7_;
      r_448__6_ <= r_n_448__6_;
      r_448__5_ <= r_n_448__5_;
      r_448__4_ <= r_n_448__4_;
      r_448__3_ <= r_n_448__3_;
      r_448__2_ <= r_n_448__2_;
      r_448__1_ <= r_n_448__1_;
      r_448__0_ <= r_n_448__0_;
    end 
    if(N4033) begin
      r_449__63_ <= r_n_449__63_;
      r_449__62_ <= r_n_449__62_;
      r_449__61_ <= r_n_449__61_;
      r_449__60_ <= r_n_449__60_;
      r_449__59_ <= r_n_449__59_;
      r_449__58_ <= r_n_449__58_;
      r_449__57_ <= r_n_449__57_;
      r_449__56_ <= r_n_449__56_;
      r_449__55_ <= r_n_449__55_;
      r_449__54_ <= r_n_449__54_;
      r_449__53_ <= r_n_449__53_;
      r_449__52_ <= r_n_449__52_;
      r_449__51_ <= r_n_449__51_;
      r_449__50_ <= r_n_449__50_;
      r_449__49_ <= r_n_449__49_;
      r_449__48_ <= r_n_449__48_;
      r_449__47_ <= r_n_449__47_;
      r_449__46_ <= r_n_449__46_;
      r_449__45_ <= r_n_449__45_;
      r_449__44_ <= r_n_449__44_;
      r_449__43_ <= r_n_449__43_;
      r_449__42_ <= r_n_449__42_;
      r_449__41_ <= r_n_449__41_;
      r_449__40_ <= r_n_449__40_;
      r_449__39_ <= r_n_449__39_;
      r_449__38_ <= r_n_449__38_;
      r_449__37_ <= r_n_449__37_;
      r_449__36_ <= r_n_449__36_;
      r_449__35_ <= r_n_449__35_;
      r_449__34_ <= r_n_449__34_;
      r_449__33_ <= r_n_449__33_;
      r_449__32_ <= r_n_449__32_;
      r_449__31_ <= r_n_449__31_;
      r_449__30_ <= r_n_449__30_;
      r_449__29_ <= r_n_449__29_;
      r_449__28_ <= r_n_449__28_;
      r_449__27_ <= r_n_449__27_;
      r_449__26_ <= r_n_449__26_;
      r_449__25_ <= r_n_449__25_;
      r_449__24_ <= r_n_449__24_;
      r_449__23_ <= r_n_449__23_;
      r_449__22_ <= r_n_449__22_;
      r_449__21_ <= r_n_449__21_;
      r_449__20_ <= r_n_449__20_;
      r_449__19_ <= r_n_449__19_;
      r_449__18_ <= r_n_449__18_;
      r_449__17_ <= r_n_449__17_;
      r_449__16_ <= r_n_449__16_;
      r_449__15_ <= r_n_449__15_;
      r_449__14_ <= r_n_449__14_;
      r_449__13_ <= r_n_449__13_;
      r_449__12_ <= r_n_449__12_;
      r_449__11_ <= r_n_449__11_;
      r_449__10_ <= r_n_449__10_;
      r_449__9_ <= r_n_449__9_;
      r_449__8_ <= r_n_449__8_;
      r_449__7_ <= r_n_449__7_;
      r_449__6_ <= r_n_449__6_;
      r_449__5_ <= r_n_449__5_;
      r_449__4_ <= r_n_449__4_;
      r_449__3_ <= r_n_449__3_;
      r_449__2_ <= r_n_449__2_;
      r_449__1_ <= r_n_449__1_;
      r_449__0_ <= r_n_449__0_;
    end 
    if(N4034) begin
      r_450__63_ <= r_n_450__63_;
      r_450__62_ <= r_n_450__62_;
      r_450__61_ <= r_n_450__61_;
      r_450__60_ <= r_n_450__60_;
      r_450__59_ <= r_n_450__59_;
      r_450__58_ <= r_n_450__58_;
      r_450__57_ <= r_n_450__57_;
      r_450__56_ <= r_n_450__56_;
      r_450__55_ <= r_n_450__55_;
      r_450__54_ <= r_n_450__54_;
      r_450__53_ <= r_n_450__53_;
      r_450__52_ <= r_n_450__52_;
      r_450__51_ <= r_n_450__51_;
      r_450__50_ <= r_n_450__50_;
      r_450__49_ <= r_n_450__49_;
      r_450__48_ <= r_n_450__48_;
      r_450__47_ <= r_n_450__47_;
      r_450__46_ <= r_n_450__46_;
      r_450__45_ <= r_n_450__45_;
      r_450__44_ <= r_n_450__44_;
      r_450__43_ <= r_n_450__43_;
      r_450__42_ <= r_n_450__42_;
      r_450__41_ <= r_n_450__41_;
      r_450__40_ <= r_n_450__40_;
      r_450__39_ <= r_n_450__39_;
      r_450__38_ <= r_n_450__38_;
      r_450__37_ <= r_n_450__37_;
      r_450__36_ <= r_n_450__36_;
      r_450__35_ <= r_n_450__35_;
      r_450__34_ <= r_n_450__34_;
      r_450__33_ <= r_n_450__33_;
      r_450__32_ <= r_n_450__32_;
      r_450__31_ <= r_n_450__31_;
      r_450__30_ <= r_n_450__30_;
      r_450__29_ <= r_n_450__29_;
      r_450__28_ <= r_n_450__28_;
      r_450__27_ <= r_n_450__27_;
      r_450__26_ <= r_n_450__26_;
      r_450__25_ <= r_n_450__25_;
      r_450__24_ <= r_n_450__24_;
      r_450__23_ <= r_n_450__23_;
      r_450__22_ <= r_n_450__22_;
      r_450__21_ <= r_n_450__21_;
      r_450__20_ <= r_n_450__20_;
      r_450__19_ <= r_n_450__19_;
      r_450__18_ <= r_n_450__18_;
      r_450__17_ <= r_n_450__17_;
      r_450__16_ <= r_n_450__16_;
      r_450__15_ <= r_n_450__15_;
      r_450__14_ <= r_n_450__14_;
      r_450__13_ <= r_n_450__13_;
      r_450__12_ <= r_n_450__12_;
      r_450__11_ <= r_n_450__11_;
      r_450__10_ <= r_n_450__10_;
      r_450__9_ <= r_n_450__9_;
      r_450__8_ <= r_n_450__8_;
      r_450__7_ <= r_n_450__7_;
      r_450__6_ <= r_n_450__6_;
      r_450__5_ <= r_n_450__5_;
      r_450__4_ <= r_n_450__4_;
      r_450__3_ <= r_n_450__3_;
      r_450__2_ <= r_n_450__2_;
      r_450__1_ <= r_n_450__1_;
      r_450__0_ <= r_n_450__0_;
    end 
    if(N4035) begin
      r_451__63_ <= r_n_451__63_;
      r_451__62_ <= r_n_451__62_;
      r_451__61_ <= r_n_451__61_;
      r_451__60_ <= r_n_451__60_;
      r_451__59_ <= r_n_451__59_;
      r_451__58_ <= r_n_451__58_;
      r_451__57_ <= r_n_451__57_;
      r_451__56_ <= r_n_451__56_;
      r_451__55_ <= r_n_451__55_;
      r_451__54_ <= r_n_451__54_;
      r_451__53_ <= r_n_451__53_;
      r_451__52_ <= r_n_451__52_;
      r_451__51_ <= r_n_451__51_;
      r_451__50_ <= r_n_451__50_;
      r_451__49_ <= r_n_451__49_;
      r_451__48_ <= r_n_451__48_;
      r_451__47_ <= r_n_451__47_;
      r_451__46_ <= r_n_451__46_;
      r_451__45_ <= r_n_451__45_;
      r_451__44_ <= r_n_451__44_;
      r_451__43_ <= r_n_451__43_;
      r_451__42_ <= r_n_451__42_;
      r_451__41_ <= r_n_451__41_;
      r_451__40_ <= r_n_451__40_;
      r_451__39_ <= r_n_451__39_;
      r_451__38_ <= r_n_451__38_;
      r_451__37_ <= r_n_451__37_;
      r_451__36_ <= r_n_451__36_;
      r_451__35_ <= r_n_451__35_;
      r_451__34_ <= r_n_451__34_;
      r_451__33_ <= r_n_451__33_;
      r_451__32_ <= r_n_451__32_;
      r_451__31_ <= r_n_451__31_;
      r_451__30_ <= r_n_451__30_;
      r_451__29_ <= r_n_451__29_;
      r_451__28_ <= r_n_451__28_;
      r_451__27_ <= r_n_451__27_;
      r_451__26_ <= r_n_451__26_;
      r_451__25_ <= r_n_451__25_;
      r_451__24_ <= r_n_451__24_;
      r_451__23_ <= r_n_451__23_;
      r_451__22_ <= r_n_451__22_;
      r_451__21_ <= r_n_451__21_;
      r_451__20_ <= r_n_451__20_;
      r_451__19_ <= r_n_451__19_;
      r_451__18_ <= r_n_451__18_;
      r_451__17_ <= r_n_451__17_;
      r_451__16_ <= r_n_451__16_;
      r_451__15_ <= r_n_451__15_;
      r_451__14_ <= r_n_451__14_;
      r_451__13_ <= r_n_451__13_;
      r_451__12_ <= r_n_451__12_;
      r_451__11_ <= r_n_451__11_;
      r_451__10_ <= r_n_451__10_;
      r_451__9_ <= r_n_451__9_;
      r_451__8_ <= r_n_451__8_;
      r_451__7_ <= r_n_451__7_;
      r_451__6_ <= r_n_451__6_;
      r_451__5_ <= r_n_451__5_;
      r_451__4_ <= r_n_451__4_;
      r_451__3_ <= r_n_451__3_;
      r_451__2_ <= r_n_451__2_;
      r_451__1_ <= r_n_451__1_;
      r_451__0_ <= r_n_451__0_;
    end 
    if(N4036) begin
      r_452__63_ <= r_n_452__63_;
      r_452__62_ <= r_n_452__62_;
      r_452__61_ <= r_n_452__61_;
      r_452__60_ <= r_n_452__60_;
      r_452__59_ <= r_n_452__59_;
      r_452__58_ <= r_n_452__58_;
      r_452__57_ <= r_n_452__57_;
      r_452__56_ <= r_n_452__56_;
      r_452__55_ <= r_n_452__55_;
      r_452__54_ <= r_n_452__54_;
      r_452__53_ <= r_n_452__53_;
      r_452__52_ <= r_n_452__52_;
      r_452__51_ <= r_n_452__51_;
      r_452__50_ <= r_n_452__50_;
      r_452__49_ <= r_n_452__49_;
      r_452__48_ <= r_n_452__48_;
      r_452__47_ <= r_n_452__47_;
      r_452__46_ <= r_n_452__46_;
      r_452__45_ <= r_n_452__45_;
      r_452__44_ <= r_n_452__44_;
      r_452__43_ <= r_n_452__43_;
      r_452__42_ <= r_n_452__42_;
      r_452__41_ <= r_n_452__41_;
      r_452__40_ <= r_n_452__40_;
      r_452__39_ <= r_n_452__39_;
      r_452__38_ <= r_n_452__38_;
      r_452__37_ <= r_n_452__37_;
      r_452__36_ <= r_n_452__36_;
      r_452__35_ <= r_n_452__35_;
      r_452__34_ <= r_n_452__34_;
      r_452__33_ <= r_n_452__33_;
      r_452__32_ <= r_n_452__32_;
      r_452__31_ <= r_n_452__31_;
      r_452__30_ <= r_n_452__30_;
      r_452__29_ <= r_n_452__29_;
      r_452__28_ <= r_n_452__28_;
      r_452__27_ <= r_n_452__27_;
      r_452__26_ <= r_n_452__26_;
      r_452__25_ <= r_n_452__25_;
      r_452__24_ <= r_n_452__24_;
      r_452__23_ <= r_n_452__23_;
      r_452__22_ <= r_n_452__22_;
      r_452__21_ <= r_n_452__21_;
      r_452__20_ <= r_n_452__20_;
      r_452__19_ <= r_n_452__19_;
      r_452__18_ <= r_n_452__18_;
      r_452__17_ <= r_n_452__17_;
      r_452__16_ <= r_n_452__16_;
      r_452__15_ <= r_n_452__15_;
      r_452__14_ <= r_n_452__14_;
      r_452__13_ <= r_n_452__13_;
      r_452__12_ <= r_n_452__12_;
      r_452__11_ <= r_n_452__11_;
      r_452__10_ <= r_n_452__10_;
      r_452__9_ <= r_n_452__9_;
      r_452__8_ <= r_n_452__8_;
      r_452__7_ <= r_n_452__7_;
      r_452__6_ <= r_n_452__6_;
      r_452__5_ <= r_n_452__5_;
      r_452__4_ <= r_n_452__4_;
      r_452__3_ <= r_n_452__3_;
      r_452__2_ <= r_n_452__2_;
      r_452__1_ <= r_n_452__1_;
      r_452__0_ <= r_n_452__0_;
    end 
    if(N4037) begin
      r_453__63_ <= r_n_453__63_;
      r_453__62_ <= r_n_453__62_;
      r_453__61_ <= r_n_453__61_;
      r_453__60_ <= r_n_453__60_;
      r_453__59_ <= r_n_453__59_;
      r_453__58_ <= r_n_453__58_;
      r_453__57_ <= r_n_453__57_;
      r_453__56_ <= r_n_453__56_;
      r_453__55_ <= r_n_453__55_;
      r_453__54_ <= r_n_453__54_;
      r_453__53_ <= r_n_453__53_;
      r_453__52_ <= r_n_453__52_;
      r_453__51_ <= r_n_453__51_;
      r_453__50_ <= r_n_453__50_;
      r_453__49_ <= r_n_453__49_;
      r_453__48_ <= r_n_453__48_;
      r_453__47_ <= r_n_453__47_;
      r_453__46_ <= r_n_453__46_;
      r_453__45_ <= r_n_453__45_;
      r_453__44_ <= r_n_453__44_;
      r_453__43_ <= r_n_453__43_;
      r_453__42_ <= r_n_453__42_;
      r_453__41_ <= r_n_453__41_;
      r_453__40_ <= r_n_453__40_;
      r_453__39_ <= r_n_453__39_;
      r_453__38_ <= r_n_453__38_;
      r_453__37_ <= r_n_453__37_;
      r_453__36_ <= r_n_453__36_;
      r_453__35_ <= r_n_453__35_;
      r_453__34_ <= r_n_453__34_;
      r_453__33_ <= r_n_453__33_;
      r_453__32_ <= r_n_453__32_;
      r_453__31_ <= r_n_453__31_;
      r_453__30_ <= r_n_453__30_;
      r_453__29_ <= r_n_453__29_;
      r_453__28_ <= r_n_453__28_;
      r_453__27_ <= r_n_453__27_;
      r_453__26_ <= r_n_453__26_;
      r_453__25_ <= r_n_453__25_;
      r_453__24_ <= r_n_453__24_;
      r_453__23_ <= r_n_453__23_;
      r_453__22_ <= r_n_453__22_;
      r_453__21_ <= r_n_453__21_;
      r_453__20_ <= r_n_453__20_;
      r_453__19_ <= r_n_453__19_;
      r_453__18_ <= r_n_453__18_;
      r_453__17_ <= r_n_453__17_;
      r_453__16_ <= r_n_453__16_;
      r_453__15_ <= r_n_453__15_;
      r_453__14_ <= r_n_453__14_;
      r_453__13_ <= r_n_453__13_;
      r_453__12_ <= r_n_453__12_;
      r_453__11_ <= r_n_453__11_;
      r_453__10_ <= r_n_453__10_;
      r_453__9_ <= r_n_453__9_;
      r_453__8_ <= r_n_453__8_;
      r_453__7_ <= r_n_453__7_;
      r_453__6_ <= r_n_453__6_;
      r_453__5_ <= r_n_453__5_;
      r_453__4_ <= r_n_453__4_;
      r_453__3_ <= r_n_453__3_;
      r_453__2_ <= r_n_453__2_;
      r_453__1_ <= r_n_453__1_;
      r_453__0_ <= r_n_453__0_;
    end 
    if(N4038) begin
      r_454__63_ <= r_n_454__63_;
      r_454__62_ <= r_n_454__62_;
      r_454__61_ <= r_n_454__61_;
      r_454__60_ <= r_n_454__60_;
      r_454__59_ <= r_n_454__59_;
      r_454__58_ <= r_n_454__58_;
      r_454__57_ <= r_n_454__57_;
      r_454__56_ <= r_n_454__56_;
      r_454__55_ <= r_n_454__55_;
      r_454__54_ <= r_n_454__54_;
      r_454__53_ <= r_n_454__53_;
      r_454__52_ <= r_n_454__52_;
      r_454__51_ <= r_n_454__51_;
      r_454__50_ <= r_n_454__50_;
      r_454__49_ <= r_n_454__49_;
      r_454__48_ <= r_n_454__48_;
      r_454__47_ <= r_n_454__47_;
      r_454__46_ <= r_n_454__46_;
      r_454__45_ <= r_n_454__45_;
      r_454__44_ <= r_n_454__44_;
      r_454__43_ <= r_n_454__43_;
      r_454__42_ <= r_n_454__42_;
      r_454__41_ <= r_n_454__41_;
      r_454__40_ <= r_n_454__40_;
      r_454__39_ <= r_n_454__39_;
      r_454__38_ <= r_n_454__38_;
      r_454__37_ <= r_n_454__37_;
      r_454__36_ <= r_n_454__36_;
      r_454__35_ <= r_n_454__35_;
      r_454__34_ <= r_n_454__34_;
      r_454__33_ <= r_n_454__33_;
      r_454__32_ <= r_n_454__32_;
      r_454__31_ <= r_n_454__31_;
      r_454__30_ <= r_n_454__30_;
      r_454__29_ <= r_n_454__29_;
      r_454__28_ <= r_n_454__28_;
      r_454__27_ <= r_n_454__27_;
      r_454__26_ <= r_n_454__26_;
      r_454__25_ <= r_n_454__25_;
      r_454__24_ <= r_n_454__24_;
      r_454__23_ <= r_n_454__23_;
      r_454__22_ <= r_n_454__22_;
      r_454__21_ <= r_n_454__21_;
      r_454__20_ <= r_n_454__20_;
      r_454__19_ <= r_n_454__19_;
      r_454__18_ <= r_n_454__18_;
      r_454__17_ <= r_n_454__17_;
      r_454__16_ <= r_n_454__16_;
      r_454__15_ <= r_n_454__15_;
      r_454__14_ <= r_n_454__14_;
      r_454__13_ <= r_n_454__13_;
      r_454__12_ <= r_n_454__12_;
      r_454__11_ <= r_n_454__11_;
      r_454__10_ <= r_n_454__10_;
      r_454__9_ <= r_n_454__9_;
      r_454__8_ <= r_n_454__8_;
      r_454__7_ <= r_n_454__7_;
      r_454__6_ <= r_n_454__6_;
      r_454__5_ <= r_n_454__5_;
      r_454__4_ <= r_n_454__4_;
      r_454__3_ <= r_n_454__3_;
      r_454__2_ <= r_n_454__2_;
      r_454__1_ <= r_n_454__1_;
      r_454__0_ <= r_n_454__0_;
    end 
    if(N4039) begin
      r_455__63_ <= r_n_455__63_;
      r_455__62_ <= r_n_455__62_;
      r_455__61_ <= r_n_455__61_;
      r_455__60_ <= r_n_455__60_;
      r_455__59_ <= r_n_455__59_;
      r_455__58_ <= r_n_455__58_;
      r_455__57_ <= r_n_455__57_;
      r_455__56_ <= r_n_455__56_;
      r_455__55_ <= r_n_455__55_;
      r_455__54_ <= r_n_455__54_;
      r_455__53_ <= r_n_455__53_;
      r_455__52_ <= r_n_455__52_;
      r_455__51_ <= r_n_455__51_;
      r_455__50_ <= r_n_455__50_;
      r_455__49_ <= r_n_455__49_;
      r_455__48_ <= r_n_455__48_;
      r_455__47_ <= r_n_455__47_;
      r_455__46_ <= r_n_455__46_;
      r_455__45_ <= r_n_455__45_;
      r_455__44_ <= r_n_455__44_;
      r_455__43_ <= r_n_455__43_;
      r_455__42_ <= r_n_455__42_;
      r_455__41_ <= r_n_455__41_;
      r_455__40_ <= r_n_455__40_;
      r_455__39_ <= r_n_455__39_;
      r_455__38_ <= r_n_455__38_;
      r_455__37_ <= r_n_455__37_;
      r_455__36_ <= r_n_455__36_;
      r_455__35_ <= r_n_455__35_;
      r_455__34_ <= r_n_455__34_;
      r_455__33_ <= r_n_455__33_;
      r_455__32_ <= r_n_455__32_;
      r_455__31_ <= r_n_455__31_;
      r_455__30_ <= r_n_455__30_;
      r_455__29_ <= r_n_455__29_;
      r_455__28_ <= r_n_455__28_;
      r_455__27_ <= r_n_455__27_;
      r_455__26_ <= r_n_455__26_;
      r_455__25_ <= r_n_455__25_;
      r_455__24_ <= r_n_455__24_;
      r_455__23_ <= r_n_455__23_;
      r_455__22_ <= r_n_455__22_;
      r_455__21_ <= r_n_455__21_;
      r_455__20_ <= r_n_455__20_;
      r_455__19_ <= r_n_455__19_;
      r_455__18_ <= r_n_455__18_;
      r_455__17_ <= r_n_455__17_;
      r_455__16_ <= r_n_455__16_;
      r_455__15_ <= r_n_455__15_;
      r_455__14_ <= r_n_455__14_;
      r_455__13_ <= r_n_455__13_;
      r_455__12_ <= r_n_455__12_;
      r_455__11_ <= r_n_455__11_;
      r_455__10_ <= r_n_455__10_;
      r_455__9_ <= r_n_455__9_;
      r_455__8_ <= r_n_455__8_;
      r_455__7_ <= r_n_455__7_;
      r_455__6_ <= r_n_455__6_;
      r_455__5_ <= r_n_455__5_;
      r_455__4_ <= r_n_455__4_;
      r_455__3_ <= r_n_455__3_;
      r_455__2_ <= r_n_455__2_;
      r_455__1_ <= r_n_455__1_;
      r_455__0_ <= r_n_455__0_;
    end 
    if(N4040) begin
      r_456__63_ <= r_n_456__63_;
      r_456__62_ <= r_n_456__62_;
      r_456__61_ <= r_n_456__61_;
      r_456__60_ <= r_n_456__60_;
      r_456__59_ <= r_n_456__59_;
      r_456__58_ <= r_n_456__58_;
      r_456__57_ <= r_n_456__57_;
      r_456__56_ <= r_n_456__56_;
      r_456__55_ <= r_n_456__55_;
      r_456__54_ <= r_n_456__54_;
      r_456__53_ <= r_n_456__53_;
      r_456__52_ <= r_n_456__52_;
      r_456__51_ <= r_n_456__51_;
      r_456__50_ <= r_n_456__50_;
      r_456__49_ <= r_n_456__49_;
      r_456__48_ <= r_n_456__48_;
      r_456__47_ <= r_n_456__47_;
      r_456__46_ <= r_n_456__46_;
      r_456__45_ <= r_n_456__45_;
      r_456__44_ <= r_n_456__44_;
      r_456__43_ <= r_n_456__43_;
      r_456__42_ <= r_n_456__42_;
      r_456__41_ <= r_n_456__41_;
      r_456__40_ <= r_n_456__40_;
      r_456__39_ <= r_n_456__39_;
      r_456__38_ <= r_n_456__38_;
      r_456__37_ <= r_n_456__37_;
      r_456__36_ <= r_n_456__36_;
      r_456__35_ <= r_n_456__35_;
      r_456__34_ <= r_n_456__34_;
      r_456__33_ <= r_n_456__33_;
      r_456__32_ <= r_n_456__32_;
      r_456__31_ <= r_n_456__31_;
      r_456__30_ <= r_n_456__30_;
      r_456__29_ <= r_n_456__29_;
      r_456__28_ <= r_n_456__28_;
      r_456__27_ <= r_n_456__27_;
      r_456__26_ <= r_n_456__26_;
      r_456__25_ <= r_n_456__25_;
      r_456__24_ <= r_n_456__24_;
      r_456__23_ <= r_n_456__23_;
      r_456__22_ <= r_n_456__22_;
      r_456__21_ <= r_n_456__21_;
      r_456__20_ <= r_n_456__20_;
      r_456__19_ <= r_n_456__19_;
      r_456__18_ <= r_n_456__18_;
      r_456__17_ <= r_n_456__17_;
      r_456__16_ <= r_n_456__16_;
      r_456__15_ <= r_n_456__15_;
      r_456__14_ <= r_n_456__14_;
      r_456__13_ <= r_n_456__13_;
      r_456__12_ <= r_n_456__12_;
      r_456__11_ <= r_n_456__11_;
      r_456__10_ <= r_n_456__10_;
      r_456__9_ <= r_n_456__9_;
      r_456__8_ <= r_n_456__8_;
      r_456__7_ <= r_n_456__7_;
      r_456__6_ <= r_n_456__6_;
      r_456__5_ <= r_n_456__5_;
      r_456__4_ <= r_n_456__4_;
      r_456__3_ <= r_n_456__3_;
      r_456__2_ <= r_n_456__2_;
      r_456__1_ <= r_n_456__1_;
      r_456__0_ <= r_n_456__0_;
    end 
    if(N4041) begin
      r_457__63_ <= r_n_457__63_;
      r_457__62_ <= r_n_457__62_;
      r_457__61_ <= r_n_457__61_;
      r_457__60_ <= r_n_457__60_;
      r_457__59_ <= r_n_457__59_;
      r_457__58_ <= r_n_457__58_;
      r_457__57_ <= r_n_457__57_;
      r_457__56_ <= r_n_457__56_;
      r_457__55_ <= r_n_457__55_;
      r_457__54_ <= r_n_457__54_;
      r_457__53_ <= r_n_457__53_;
      r_457__52_ <= r_n_457__52_;
      r_457__51_ <= r_n_457__51_;
      r_457__50_ <= r_n_457__50_;
      r_457__49_ <= r_n_457__49_;
      r_457__48_ <= r_n_457__48_;
      r_457__47_ <= r_n_457__47_;
      r_457__46_ <= r_n_457__46_;
      r_457__45_ <= r_n_457__45_;
      r_457__44_ <= r_n_457__44_;
      r_457__43_ <= r_n_457__43_;
      r_457__42_ <= r_n_457__42_;
      r_457__41_ <= r_n_457__41_;
      r_457__40_ <= r_n_457__40_;
      r_457__39_ <= r_n_457__39_;
      r_457__38_ <= r_n_457__38_;
      r_457__37_ <= r_n_457__37_;
      r_457__36_ <= r_n_457__36_;
      r_457__35_ <= r_n_457__35_;
      r_457__34_ <= r_n_457__34_;
      r_457__33_ <= r_n_457__33_;
      r_457__32_ <= r_n_457__32_;
      r_457__31_ <= r_n_457__31_;
      r_457__30_ <= r_n_457__30_;
      r_457__29_ <= r_n_457__29_;
      r_457__28_ <= r_n_457__28_;
      r_457__27_ <= r_n_457__27_;
      r_457__26_ <= r_n_457__26_;
      r_457__25_ <= r_n_457__25_;
      r_457__24_ <= r_n_457__24_;
      r_457__23_ <= r_n_457__23_;
      r_457__22_ <= r_n_457__22_;
      r_457__21_ <= r_n_457__21_;
      r_457__20_ <= r_n_457__20_;
      r_457__19_ <= r_n_457__19_;
      r_457__18_ <= r_n_457__18_;
      r_457__17_ <= r_n_457__17_;
      r_457__16_ <= r_n_457__16_;
      r_457__15_ <= r_n_457__15_;
      r_457__14_ <= r_n_457__14_;
      r_457__13_ <= r_n_457__13_;
      r_457__12_ <= r_n_457__12_;
      r_457__11_ <= r_n_457__11_;
      r_457__10_ <= r_n_457__10_;
      r_457__9_ <= r_n_457__9_;
      r_457__8_ <= r_n_457__8_;
      r_457__7_ <= r_n_457__7_;
      r_457__6_ <= r_n_457__6_;
      r_457__5_ <= r_n_457__5_;
      r_457__4_ <= r_n_457__4_;
      r_457__3_ <= r_n_457__3_;
      r_457__2_ <= r_n_457__2_;
      r_457__1_ <= r_n_457__1_;
      r_457__0_ <= r_n_457__0_;
    end 
    if(N4042) begin
      r_458__63_ <= r_n_458__63_;
      r_458__62_ <= r_n_458__62_;
      r_458__61_ <= r_n_458__61_;
      r_458__60_ <= r_n_458__60_;
      r_458__59_ <= r_n_458__59_;
      r_458__58_ <= r_n_458__58_;
      r_458__57_ <= r_n_458__57_;
      r_458__56_ <= r_n_458__56_;
      r_458__55_ <= r_n_458__55_;
      r_458__54_ <= r_n_458__54_;
      r_458__53_ <= r_n_458__53_;
      r_458__52_ <= r_n_458__52_;
      r_458__51_ <= r_n_458__51_;
      r_458__50_ <= r_n_458__50_;
      r_458__49_ <= r_n_458__49_;
      r_458__48_ <= r_n_458__48_;
      r_458__47_ <= r_n_458__47_;
      r_458__46_ <= r_n_458__46_;
      r_458__45_ <= r_n_458__45_;
      r_458__44_ <= r_n_458__44_;
      r_458__43_ <= r_n_458__43_;
      r_458__42_ <= r_n_458__42_;
      r_458__41_ <= r_n_458__41_;
      r_458__40_ <= r_n_458__40_;
      r_458__39_ <= r_n_458__39_;
      r_458__38_ <= r_n_458__38_;
      r_458__37_ <= r_n_458__37_;
      r_458__36_ <= r_n_458__36_;
      r_458__35_ <= r_n_458__35_;
      r_458__34_ <= r_n_458__34_;
      r_458__33_ <= r_n_458__33_;
      r_458__32_ <= r_n_458__32_;
      r_458__31_ <= r_n_458__31_;
      r_458__30_ <= r_n_458__30_;
      r_458__29_ <= r_n_458__29_;
      r_458__28_ <= r_n_458__28_;
      r_458__27_ <= r_n_458__27_;
      r_458__26_ <= r_n_458__26_;
      r_458__25_ <= r_n_458__25_;
      r_458__24_ <= r_n_458__24_;
      r_458__23_ <= r_n_458__23_;
      r_458__22_ <= r_n_458__22_;
      r_458__21_ <= r_n_458__21_;
      r_458__20_ <= r_n_458__20_;
      r_458__19_ <= r_n_458__19_;
      r_458__18_ <= r_n_458__18_;
      r_458__17_ <= r_n_458__17_;
      r_458__16_ <= r_n_458__16_;
      r_458__15_ <= r_n_458__15_;
      r_458__14_ <= r_n_458__14_;
      r_458__13_ <= r_n_458__13_;
      r_458__12_ <= r_n_458__12_;
      r_458__11_ <= r_n_458__11_;
      r_458__10_ <= r_n_458__10_;
      r_458__9_ <= r_n_458__9_;
      r_458__8_ <= r_n_458__8_;
      r_458__7_ <= r_n_458__7_;
      r_458__6_ <= r_n_458__6_;
      r_458__5_ <= r_n_458__5_;
      r_458__4_ <= r_n_458__4_;
      r_458__3_ <= r_n_458__3_;
      r_458__2_ <= r_n_458__2_;
      r_458__1_ <= r_n_458__1_;
      r_458__0_ <= r_n_458__0_;
    end 
    if(N4043) begin
      r_459__63_ <= r_n_459__63_;
      r_459__62_ <= r_n_459__62_;
      r_459__61_ <= r_n_459__61_;
      r_459__60_ <= r_n_459__60_;
      r_459__59_ <= r_n_459__59_;
      r_459__58_ <= r_n_459__58_;
      r_459__57_ <= r_n_459__57_;
      r_459__56_ <= r_n_459__56_;
      r_459__55_ <= r_n_459__55_;
      r_459__54_ <= r_n_459__54_;
      r_459__53_ <= r_n_459__53_;
      r_459__52_ <= r_n_459__52_;
      r_459__51_ <= r_n_459__51_;
      r_459__50_ <= r_n_459__50_;
      r_459__49_ <= r_n_459__49_;
      r_459__48_ <= r_n_459__48_;
      r_459__47_ <= r_n_459__47_;
      r_459__46_ <= r_n_459__46_;
      r_459__45_ <= r_n_459__45_;
      r_459__44_ <= r_n_459__44_;
      r_459__43_ <= r_n_459__43_;
      r_459__42_ <= r_n_459__42_;
      r_459__41_ <= r_n_459__41_;
      r_459__40_ <= r_n_459__40_;
      r_459__39_ <= r_n_459__39_;
      r_459__38_ <= r_n_459__38_;
      r_459__37_ <= r_n_459__37_;
      r_459__36_ <= r_n_459__36_;
      r_459__35_ <= r_n_459__35_;
      r_459__34_ <= r_n_459__34_;
      r_459__33_ <= r_n_459__33_;
      r_459__32_ <= r_n_459__32_;
      r_459__31_ <= r_n_459__31_;
      r_459__30_ <= r_n_459__30_;
      r_459__29_ <= r_n_459__29_;
      r_459__28_ <= r_n_459__28_;
      r_459__27_ <= r_n_459__27_;
      r_459__26_ <= r_n_459__26_;
      r_459__25_ <= r_n_459__25_;
      r_459__24_ <= r_n_459__24_;
      r_459__23_ <= r_n_459__23_;
      r_459__22_ <= r_n_459__22_;
      r_459__21_ <= r_n_459__21_;
      r_459__20_ <= r_n_459__20_;
      r_459__19_ <= r_n_459__19_;
      r_459__18_ <= r_n_459__18_;
      r_459__17_ <= r_n_459__17_;
      r_459__16_ <= r_n_459__16_;
      r_459__15_ <= r_n_459__15_;
      r_459__14_ <= r_n_459__14_;
      r_459__13_ <= r_n_459__13_;
      r_459__12_ <= r_n_459__12_;
      r_459__11_ <= r_n_459__11_;
      r_459__10_ <= r_n_459__10_;
      r_459__9_ <= r_n_459__9_;
      r_459__8_ <= r_n_459__8_;
      r_459__7_ <= r_n_459__7_;
      r_459__6_ <= r_n_459__6_;
      r_459__5_ <= r_n_459__5_;
      r_459__4_ <= r_n_459__4_;
      r_459__3_ <= r_n_459__3_;
      r_459__2_ <= r_n_459__2_;
      r_459__1_ <= r_n_459__1_;
      r_459__0_ <= r_n_459__0_;
    end 
    if(N4044) begin
      r_460__63_ <= r_n_460__63_;
      r_460__62_ <= r_n_460__62_;
      r_460__61_ <= r_n_460__61_;
      r_460__60_ <= r_n_460__60_;
      r_460__59_ <= r_n_460__59_;
      r_460__58_ <= r_n_460__58_;
      r_460__57_ <= r_n_460__57_;
      r_460__56_ <= r_n_460__56_;
      r_460__55_ <= r_n_460__55_;
      r_460__54_ <= r_n_460__54_;
      r_460__53_ <= r_n_460__53_;
      r_460__52_ <= r_n_460__52_;
      r_460__51_ <= r_n_460__51_;
      r_460__50_ <= r_n_460__50_;
      r_460__49_ <= r_n_460__49_;
      r_460__48_ <= r_n_460__48_;
      r_460__47_ <= r_n_460__47_;
      r_460__46_ <= r_n_460__46_;
      r_460__45_ <= r_n_460__45_;
      r_460__44_ <= r_n_460__44_;
      r_460__43_ <= r_n_460__43_;
      r_460__42_ <= r_n_460__42_;
      r_460__41_ <= r_n_460__41_;
      r_460__40_ <= r_n_460__40_;
      r_460__39_ <= r_n_460__39_;
      r_460__38_ <= r_n_460__38_;
      r_460__37_ <= r_n_460__37_;
      r_460__36_ <= r_n_460__36_;
      r_460__35_ <= r_n_460__35_;
      r_460__34_ <= r_n_460__34_;
      r_460__33_ <= r_n_460__33_;
      r_460__32_ <= r_n_460__32_;
      r_460__31_ <= r_n_460__31_;
      r_460__30_ <= r_n_460__30_;
      r_460__29_ <= r_n_460__29_;
      r_460__28_ <= r_n_460__28_;
      r_460__27_ <= r_n_460__27_;
      r_460__26_ <= r_n_460__26_;
      r_460__25_ <= r_n_460__25_;
      r_460__24_ <= r_n_460__24_;
      r_460__23_ <= r_n_460__23_;
      r_460__22_ <= r_n_460__22_;
      r_460__21_ <= r_n_460__21_;
      r_460__20_ <= r_n_460__20_;
      r_460__19_ <= r_n_460__19_;
      r_460__18_ <= r_n_460__18_;
      r_460__17_ <= r_n_460__17_;
      r_460__16_ <= r_n_460__16_;
      r_460__15_ <= r_n_460__15_;
      r_460__14_ <= r_n_460__14_;
      r_460__13_ <= r_n_460__13_;
      r_460__12_ <= r_n_460__12_;
      r_460__11_ <= r_n_460__11_;
      r_460__10_ <= r_n_460__10_;
      r_460__9_ <= r_n_460__9_;
      r_460__8_ <= r_n_460__8_;
      r_460__7_ <= r_n_460__7_;
      r_460__6_ <= r_n_460__6_;
      r_460__5_ <= r_n_460__5_;
      r_460__4_ <= r_n_460__4_;
      r_460__3_ <= r_n_460__3_;
      r_460__2_ <= r_n_460__2_;
      r_460__1_ <= r_n_460__1_;
      r_460__0_ <= r_n_460__0_;
    end 
    if(N4045) begin
      r_461__63_ <= r_n_461__63_;
      r_461__62_ <= r_n_461__62_;
      r_461__61_ <= r_n_461__61_;
      r_461__60_ <= r_n_461__60_;
      r_461__59_ <= r_n_461__59_;
      r_461__58_ <= r_n_461__58_;
      r_461__57_ <= r_n_461__57_;
      r_461__56_ <= r_n_461__56_;
      r_461__55_ <= r_n_461__55_;
      r_461__54_ <= r_n_461__54_;
      r_461__53_ <= r_n_461__53_;
      r_461__52_ <= r_n_461__52_;
      r_461__51_ <= r_n_461__51_;
      r_461__50_ <= r_n_461__50_;
      r_461__49_ <= r_n_461__49_;
      r_461__48_ <= r_n_461__48_;
      r_461__47_ <= r_n_461__47_;
      r_461__46_ <= r_n_461__46_;
      r_461__45_ <= r_n_461__45_;
      r_461__44_ <= r_n_461__44_;
      r_461__43_ <= r_n_461__43_;
      r_461__42_ <= r_n_461__42_;
      r_461__41_ <= r_n_461__41_;
      r_461__40_ <= r_n_461__40_;
      r_461__39_ <= r_n_461__39_;
      r_461__38_ <= r_n_461__38_;
      r_461__37_ <= r_n_461__37_;
      r_461__36_ <= r_n_461__36_;
      r_461__35_ <= r_n_461__35_;
      r_461__34_ <= r_n_461__34_;
      r_461__33_ <= r_n_461__33_;
      r_461__32_ <= r_n_461__32_;
      r_461__31_ <= r_n_461__31_;
      r_461__30_ <= r_n_461__30_;
      r_461__29_ <= r_n_461__29_;
      r_461__28_ <= r_n_461__28_;
      r_461__27_ <= r_n_461__27_;
      r_461__26_ <= r_n_461__26_;
      r_461__25_ <= r_n_461__25_;
      r_461__24_ <= r_n_461__24_;
      r_461__23_ <= r_n_461__23_;
      r_461__22_ <= r_n_461__22_;
      r_461__21_ <= r_n_461__21_;
      r_461__20_ <= r_n_461__20_;
      r_461__19_ <= r_n_461__19_;
      r_461__18_ <= r_n_461__18_;
      r_461__17_ <= r_n_461__17_;
      r_461__16_ <= r_n_461__16_;
      r_461__15_ <= r_n_461__15_;
      r_461__14_ <= r_n_461__14_;
      r_461__13_ <= r_n_461__13_;
      r_461__12_ <= r_n_461__12_;
      r_461__11_ <= r_n_461__11_;
      r_461__10_ <= r_n_461__10_;
      r_461__9_ <= r_n_461__9_;
      r_461__8_ <= r_n_461__8_;
      r_461__7_ <= r_n_461__7_;
      r_461__6_ <= r_n_461__6_;
      r_461__5_ <= r_n_461__5_;
      r_461__4_ <= r_n_461__4_;
      r_461__3_ <= r_n_461__3_;
      r_461__2_ <= r_n_461__2_;
      r_461__1_ <= r_n_461__1_;
      r_461__0_ <= r_n_461__0_;
    end 
    if(N4046) begin
      r_462__63_ <= r_n_462__63_;
      r_462__62_ <= r_n_462__62_;
      r_462__61_ <= r_n_462__61_;
      r_462__60_ <= r_n_462__60_;
      r_462__59_ <= r_n_462__59_;
      r_462__58_ <= r_n_462__58_;
      r_462__57_ <= r_n_462__57_;
      r_462__56_ <= r_n_462__56_;
      r_462__55_ <= r_n_462__55_;
      r_462__54_ <= r_n_462__54_;
      r_462__53_ <= r_n_462__53_;
      r_462__52_ <= r_n_462__52_;
      r_462__51_ <= r_n_462__51_;
      r_462__50_ <= r_n_462__50_;
      r_462__49_ <= r_n_462__49_;
      r_462__48_ <= r_n_462__48_;
      r_462__47_ <= r_n_462__47_;
      r_462__46_ <= r_n_462__46_;
      r_462__45_ <= r_n_462__45_;
      r_462__44_ <= r_n_462__44_;
      r_462__43_ <= r_n_462__43_;
      r_462__42_ <= r_n_462__42_;
      r_462__41_ <= r_n_462__41_;
      r_462__40_ <= r_n_462__40_;
      r_462__39_ <= r_n_462__39_;
      r_462__38_ <= r_n_462__38_;
      r_462__37_ <= r_n_462__37_;
      r_462__36_ <= r_n_462__36_;
      r_462__35_ <= r_n_462__35_;
      r_462__34_ <= r_n_462__34_;
      r_462__33_ <= r_n_462__33_;
      r_462__32_ <= r_n_462__32_;
      r_462__31_ <= r_n_462__31_;
      r_462__30_ <= r_n_462__30_;
      r_462__29_ <= r_n_462__29_;
      r_462__28_ <= r_n_462__28_;
      r_462__27_ <= r_n_462__27_;
      r_462__26_ <= r_n_462__26_;
      r_462__25_ <= r_n_462__25_;
      r_462__24_ <= r_n_462__24_;
      r_462__23_ <= r_n_462__23_;
      r_462__22_ <= r_n_462__22_;
      r_462__21_ <= r_n_462__21_;
      r_462__20_ <= r_n_462__20_;
      r_462__19_ <= r_n_462__19_;
      r_462__18_ <= r_n_462__18_;
      r_462__17_ <= r_n_462__17_;
      r_462__16_ <= r_n_462__16_;
      r_462__15_ <= r_n_462__15_;
      r_462__14_ <= r_n_462__14_;
      r_462__13_ <= r_n_462__13_;
      r_462__12_ <= r_n_462__12_;
      r_462__11_ <= r_n_462__11_;
      r_462__10_ <= r_n_462__10_;
      r_462__9_ <= r_n_462__9_;
      r_462__8_ <= r_n_462__8_;
      r_462__7_ <= r_n_462__7_;
      r_462__6_ <= r_n_462__6_;
      r_462__5_ <= r_n_462__5_;
      r_462__4_ <= r_n_462__4_;
      r_462__3_ <= r_n_462__3_;
      r_462__2_ <= r_n_462__2_;
      r_462__1_ <= r_n_462__1_;
      r_462__0_ <= r_n_462__0_;
    end 
    if(N4047) begin
      r_463__63_ <= r_n_463__63_;
      r_463__62_ <= r_n_463__62_;
      r_463__61_ <= r_n_463__61_;
      r_463__60_ <= r_n_463__60_;
      r_463__59_ <= r_n_463__59_;
      r_463__58_ <= r_n_463__58_;
      r_463__57_ <= r_n_463__57_;
      r_463__56_ <= r_n_463__56_;
      r_463__55_ <= r_n_463__55_;
      r_463__54_ <= r_n_463__54_;
      r_463__53_ <= r_n_463__53_;
      r_463__52_ <= r_n_463__52_;
      r_463__51_ <= r_n_463__51_;
      r_463__50_ <= r_n_463__50_;
      r_463__49_ <= r_n_463__49_;
      r_463__48_ <= r_n_463__48_;
      r_463__47_ <= r_n_463__47_;
      r_463__46_ <= r_n_463__46_;
      r_463__45_ <= r_n_463__45_;
      r_463__44_ <= r_n_463__44_;
      r_463__43_ <= r_n_463__43_;
      r_463__42_ <= r_n_463__42_;
      r_463__41_ <= r_n_463__41_;
      r_463__40_ <= r_n_463__40_;
      r_463__39_ <= r_n_463__39_;
      r_463__38_ <= r_n_463__38_;
      r_463__37_ <= r_n_463__37_;
      r_463__36_ <= r_n_463__36_;
      r_463__35_ <= r_n_463__35_;
      r_463__34_ <= r_n_463__34_;
      r_463__33_ <= r_n_463__33_;
      r_463__32_ <= r_n_463__32_;
      r_463__31_ <= r_n_463__31_;
      r_463__30_ <= r_n_463__30_;
      r_463__29_ <= r_n_463__29_;
      r_463__28_ <= r_n_463__28_;
      r_463__27_ <= r_n_463__27_;
      r_463__26_ <= r_n_463__26_;
      r_463__25_ <= r_n_463__25_;
      r_463__24_ <= r_n_463__24_;
      r_463__23_ <= r_n_463__23_;
      r_463__22_ <= r_n_463__22_;
      r_463__21_ <= r_n_463__21_;
      r_463__20_ <= r_n_463__20_;
      r_463__19_ <= r_n_463__19_;
      r_463__18_ <= r_n_463__18_;
      r_463__17_ <= r_n_463__17_;
      r_463__16_ <= r_n_463__16_;
      r_463__15_ <= r_n_463__15_;
      r_463__14_ <= r_n_463__14_;
      r_463__13_ <= r_n_463__13_;
      r_463__12_ <= r_n_463__12_;
      r_463__11_ <= r_n_463__11_;
      r_463__10_ <= r_n_463__10_;
      r_463__9_ <= r_n_463__9_;
      r_463__8_ <= r_n_463__8_;
      r_463__7_ <= r_n_463__7_;
      r_463__6_ <= r_n_463__6_;
      r_463__5_ <= r_n_463__5_;
      r_463__4_ <= r_n_463__4_;
      r_463__3_ <= r_n_463__3_;
      r_463__2_ <= r_n_463__2_;
      r_463__1_ <= r_n_463__1_;
      r_463__0_ <= r_n_463__0_;
    end 
    if(N4048) begin
      r_464__63_ <= r_n_464__63_;
      r_464__62_ <= r_n_464__62_;
      r_464__61_ <= r_n_464__61_;
      r_464__60_ <= r_n_464__60_;
      r_464__59_ <= r_n_464__59_;
      r_464__58_ <= r_n_464__58_;
      r_464__57_ <= r_n_464__57_;
      r_464__56_ <= r_n_464__56_;
      r_464__55_ <= r_n_464__55_;
      r_464__54_ <= r_n_464__54_;
      r_464__53_ <= r_n_464__53_;
      r_464__52_ <= r_n_464__52_;
      r_464__51_ <= r_n_464__51_;
      r_464__50_ <= r_n_464__50_;
      r_464__49_ <= r_n_464__49_;
      r_464__48_ <= r_n_464__48_;
      r_464__47_ <= r_n_464__47_;
      r_464__46_ <= r_n_464__46_;
      r_464__45_ <= r_n_464__45_;
      r_464__44_ <= r_n_464__44_;
      r_464__43_ <= r_n_464__43_;
      r_464__42_ <= r_n_464__42_;
      r_464__41_ <= r_n_464__41_;
      r_464__40_ <= r_n_464__40_;
      r_464__39_ <= r_n_464__39_;
      r_464__38_ <= r_n_464__38_;
      r_464__37_ <= r_n_464__37_;
      r_464__36_ <= r_n_464__36_;
      r_464__35_ <= r_n_464__35_;
      r_464__34_ <= r_n_464__34_;
      r_464__33_ <= r_n_464__33_;
      r_464__32_ <= r_n_464__32_;
      r_464__31_ <= r_n_464__31_;
      r_464__30_ <= r_n_464__30_;
      r_464__29_ <= r_n_464__29_;
      r_464__28_ <= r_n_464__28_;
      r_464__27_ <= r_n_464__27_;
      r_464__26_ <= r_n_464__26_;
      r_464__25_ <= r_n_464__25_;
      r_464__24_ <= r_n_464__24_;
      r_464__23_ <= r_n_464__23_;
      r_464__22_ <= r_n_464__22_;
      r_464__21_ <= r_n_464__21_;
      r_464__20_ <= r_n_464__20_;
      r_464__19_ <= r_n_464__19_;
      r_464__18_ <= r_n_464__18_;
      r_464__17_ <= r_n_464__17_;
      r_464__16_ <= r_n_464__16_;
      r_464__15_ <= r_n_464__15_;
      r_464__14_ <= r_n_464__14_;
      r_464__13_ <= r_n_464__13_;
      r_464__12_ <= r_n_464__12_;
      r_464__11_ <= r_n_464__11_;
      r_464__10_ <= r_n_464__10_;
      r_464__9_ <= r_n_464__9_;
      r_464__8_ <= r_n_464__8_;
      r_464__7_ <= r_n_464__7_;
      r_464__6_ <= r_n_464__6_;
      r_464__5_ <= r_n_464__5_;
      r_464__4_ <= r_n_464__4_;
      r_464__3_ <= r_n_464__3_;
      r_464__2_ <= r_n_464__2_;
      r_464__1_ <= r_n_464__1_;
      r_464__0_ <= r_n_464__0_;
    end 
    if(N4049) begin
      r_465__63_ <= r_n_465__63_;
      r_465__62_ <= r_n_465__62_;
      r_465__61_ <= r_n_465__61_;
      r_465__60_ <= r_n_465__60_;
      r_465__59_ <= r_n_465__59_;
      r_465__58_ <= r_n_465__58_;
      r_465__57_ <= r_n_465__57_;
      r_465__56_ <= r_n_465__56_;
      r_465__55_ <= r_n_465__55_;
      r_465__54_ <= r_n_465__54_;
      r_465__53_ <= r_n_465__53_;
      r_465__52_ <= r_n_465__52_;
      r_465__51_ <= r_n_465__51_;
      r_465__50_ <= r_n_465__50_;
      r_465__49_ <= r_n_465__49_;
      r_465__48_ <= r_n_465__48_;
      r_465__47_ <= r_n_465__47_;
      r_465__46_ <= r_n_465__46_;
      r_465__45_ <= r_n_465__45_;
      r_465__44_ <= r_n_465__44_;
      r_465__43_ <= r_n_465__43_;
      r_465__42_ <= r_n_465__42_;
      r_465__41_ <= r_n_465__41_;
      r_465__40_ <= r_n_465__40_;
      r_465__39_ <= r_n_465__39_;
      r_465__38_ <= r_n_465__38_;
      r_465__37_ <= r_n_465__37_;
      r_465__36_ <= r_n_465__36_;
      r_465__35_ <= r_n_465__35_;
      r_465__34_ <= r_n_465__34_;
      r_465__33_ <= r_n_465__33_;
      r_465__32_ <= r_n_465__32_;
      r_465__31_ <= r_n_465__31_;
      r_465__30_ <= r_n_465__30_;
      r_465__29_ <= r_n_465__29_;
      r_465__28_ <= r_n_465__28_;
      r_465__27_ <= r_n_465__27_;
      r_465__26_ <= r_n_465__26_;
      r_465__25_ <= r_n_465__25_;
      r_465__24_ <= r_n_465__24_;
      r_465__23_ <= r_n_465__23_;
      r_465__22_ <= r_n_465__22_;
      r_465__21_ <= r_n_465__21_;
      r_465__20_ <= r_n_465__20_;
      r_465__19_ <= r_n_465__19_;
      r_465__18_ <= r_n_465__18_;
      r_465__17_ <= r_n_465__17_;
      r_465__16_ <= r_n_465__16_;
      r_465__15_ <= r_n_465__15_;
      r_465__14_ <= r_n_465__14_;
      r_465__13_ <= r_n_465__13_;
      r_465__12_ <= r_n_465__12_;
      r_465__11_ <= r_n_465__11_;
      r_465__10_ <= r_n_465__10_;
      r_465__9_ <= r_n_465__9_;
      r_465__8_ <= r_n_465__8_;
      r_465__7_ <= r_n_465__7_;
      r_465__6_ <= r_n_465__6_;
      r_465__5_ <= r_n_465__5_;
      r_465__4_ <= r_n_465__4_;
      r_465__3_ <= r_n_465__3_;
      r_465__2_ <= r_n_465__2_;
      r_465__1_ <= r_n_465__1_;
      r_465__0_ <= r_n_465__0_;
    end 
    if(N4050) begin
      r_466__63_ <= r_n_466__63_;
      r_466__62_ <= r_n_466__62_;
      r_466__61_ <= r_n_466__61_;
      r_466__60_ <= r_n_466__60_;
      r_466__59_ <= r_n_466__59_;
      r_466__58_ <= r_n_466__58_;
      r_466__57_ <= r_n_466__57_;
      r_466__56_ <= r_n_466__56_;
      r_466__55_ <= r_n_466__55_;
      r_466__54_ <= r_n_466__54_;
      r_466__53_ <= r_n_466__53_;
      r_466__52_ <= r_n_466__52_;
      r_466__51_ <= r_n_466__51_;
      r_466__50_ <= r_n_466__50_;
      r_466__49_ <= r_n_466__49_;
      r_466__48_ <= r_n_466__48_;
      r_466__47_ <= r_n_466__47_;
      r_466__46_ <= r_n_466__46_;
      r_466__45_ <= r_n_466__45_;
      r_466__44_ <= r_n_466__44_;
      r_466__43_ <= r_n_466__43_;
      r_466__42_ <= r_n_466__42_;
      r_466__41_ <= r_n_466__41_;
      r_466__40_ <= r_n_466__40_;
      r_466__39_ <= r_n_466__39_;
      r_466__38_ <= r_n_466__38_;
      r_466__37_ <= r_n_466__37_;
      r_466__36_ <= r_n_466__36_;
      r_466__35_ <= r_n_466__35_;
      r_466__34_ <= r_n_466__34_;
      r_466__33_ <= r_n_466__33_;
      r_466__32_ <= r_n_466__32_;
      r_466__31_ <= r_n_466__31_;
      r_466__30_ <= r_n_466__30_;
      r_466__29_ <= r_n_466__29_;
      r_466__28_ <= r_n_466__28_;
      r_466__27_ <= r_n_466__27_;
      r_466__26_ <= r_n_466__26_;
      r_466__25_ <= r_n_466__25_;
      r_466__24_ <= r_n_466__24_;
      r_466__23_ <= r_n_466__23_;
      r_466__22_ <= r_n_466__22_;
      r_466__21_ <= r_n_466__21_;
      r_466__20_ <= r_n_466__20_;
      r_466__19_ <= r_n_466__19_;
      r_466__18_ <= r_n_466__18_;
      r_466__17_ <= r_n_466__17_;
      r_466__16_ <= r_n_466__16_;
      r_466__15_ <= r_n_466__15_;
      r_466__14_ <= r_n_466__14_;
      r_466__13_ <= r_n_466__13_;
      r_466__12_ <= r_n_466__12_;
      r_466__11_ <= r_n_466__11_;
      r_466__10_ <= r_n_466__10_;
      r_466__9_ <= r_n_466__9_;
      r_466__8_ <= r_n_466__8_;
      r_466__7_ <= r_n_466__7_;
      r_466__6_ <= r_n_466__6_;
      r_466__5_ <= r_n_466__5_;
      r_466__4_ <= r_n_466__4_;
      r_466__3_ <= r_n_466__3_;
      r_466__2_ <= r_n_466__2_;
      r_466__1_ <= r_n_466__1_;
      r_466__0_ <= r_n_466__0_;
    end 
    if(N4051) begin
      r_467__63_ <= r_n_467__63_;
      r_467__62_ <= r_n_467__62_;
      r_467__61_ <= r_n_467__61_;
      r_467__60_ <= r_n_467__60_;
      r_467__59_ <= r_n_467__59_;
      r_467__58_ <= r_n_467__58_;
      r_467__57_ <= r_n_467__57_;
      r_467__56_ <= r_n_467__56_;
      r_467__55_ <= r_n_467__55_;
      r_467__54_ <= r_n_467__54_;
      r_467__53_ <= r_n_467__53_;
      r_467__52_ <= r_n_467__52_;
      r_467__51_ <= r_n_467__51_;
      r_467__50_ <= r_n_467__50_;
      r_467__49_ <= r_n_467__49_;
      r_467__48_ <= r_n_467__48_;
      r_467__47_ <= r_n_467__47_;
      r_467__46_ <= r_n_467__46_;
      r_467__45_ <= r_n_467__45_;
      r_467__44_ <= r_n_467__44_;
      r_467__43_ <= r_n_467__43_;
      r_467__42_ <= r_n_467__42_;
      r_467__41_ <= r_n_467__41_;
      r_467__40_ <= r_n_467__40_;
      r_467__39_ <= r_n_467__39_;
      r_467__38_ <= r_n_467__38_;
      r_467__37_ <= r_n_467__37_;
      r_467__36_ <= r_n_467__36_;
      r_467__35_ <= r_n_467__35_;
      r_467__34_ <= r_n_467__34_;
      r_467__33_ <= r_n_467__33_;
      r_467__32_ <= r_n_467__32_;
      r_467__31_ <= r_n_467__31_;
      r_467__30_ <= r_n_467__30_;
      r_467__29_ <= r_n_467__29_;
      r_467__28_ <= r_n_467__28_;
      r_467__27_ <= r_n_467__27_;
      r_467__26_ <= r_n_467__26_;
      r_467__25_ <= r_n_467__25_;
      r_467__24_ <= r_n_467__24_;
      r_467__23_ <= r_n_467__23_;
      r_467__22_ <= r_n_467__22_;
      r_467__21_ <= r_n_467__21_;
      r_467__20_ <= r_n_467__20_;
      r_467__19_ <= r_n_467__19_;
      r_467__18_ <= r_n_467__18_;
      r_467__17_ <= r_n_467__17_;
      r_467__16_ <= r_n_467__16_;
      r_467__15_ <= r_n_467__15_;
      r_467__14_ <= r_n_467__14_;
      r_467__13_ <= r_n_467__13_;
      r_467__12_ <= r_n_467__12_;
      r_467__11_ <= r_n_467__11_;
      r_467__10_ <= r_n_467__10_;
      r_467__9_ <= r_n_467__9_;
      r_467__8_ <= r_n_467__8_;
      r_467__7_ <= r_n_467__7_;
      r_467__6_ <= r_n_467__6_;
      r_467__5_ <= r_n_467__5_;
      r_467__4_ <= r_n_467__4_;
      r_467__3_ <= r_n_467__3_;
      r_467__2_ <= r_n_467__2_;
      r_467__1_ <= r_n_467__1_;
      r_467__0_ <= r_n_467__0_;
    end 
    if(N4052) begin
      r_468__63_ <= r_n_468__63_;
      r_468__62_ <= r_n_468__62_;
      r_468__61_ <= r_n_468__61_;
      r_468__60_ <= r_n_468__60_;
      r_468__59_ <= r_n_468__59_;
      r_468__58_ <= r_n_468__58_;
      r_468__57_ <= r_n_468__57_;
      r_468__56_ <= r_n_468__56_;
      r_468__55_ <= r_n_468__55_;
      r_468__54_ <= r_n_468__54_;
      r_468__53_ <= r_n_468__53_;
      r_468__52_ <= r_n_468__52_;
      r_468__51_ <= r_n_468__51_;
      r_468__50_ <= r_n_468__50_;
      r_468__49_ <= r_n_468__49_;
      r_468__48_ <= r_n_468__48_;
      r_468__47_ <= r_n_468__47_;
      r_468__46_ <= r_n_468__46_;
      r_468__45_ <= r_n_468__45_;
      r_468__44_ <= r_n_468__44_;
      r_468__43_ <= r_n_468__43_;
      r_468__42_ <= r_n_468__42_;
      r_468__41_ <= r_n_468__41_;
      r_468__40_ <= r_n_468__40_;
      r_468__39_ <= r_n_468__39_;
      r_468__38_ <= r_n_468__38_;
      r_468__37_ <= r_n_468__37_;
      r_468__36_ <= r_n_468__36_;
      r_468__35_ <= r_n_468__35_;
      r_468__34_ <= r_n_468__34_;
      r_468__33_ <= r_n_468__33_;
      r_468__32_ <= r_n_468__32_;
      r_468__31_ <= r_n_468__31_;
      r_468__30_ <= r_n_468__30_;
      r_468__29_ <= r_n_468__29_;
      r_468__28_ <= r_n_468__28_;
      r_468__27_ <= r_n_468__27_;
      r_468__26_ <= r_n_468__26_;
      r_468__25_ <= r_n_468__25_;
      r_468__24_ <= r_n_468__24_;
      r_468__23_ <= r_n_468__23_;
      r_468__22_ <= r_n_468__22_;
      r_468__21_ <= r_n_468__21_;
      r_468__20_ <= r_n_468__20_;
      r_468__19_ <= r_n_468__19_;
      r_468__18_ <= r_n_468__18_;
      r_468__17_ <= r_n_468__17_;
      r_468__16_ <= r_n_468__16_;
      r_468__15_ <= r_n_468__15_;
      r_468__14_ <= r_n_468__14_;
      r_468__13_ <= r_n_468__13_;
      r_468__12_ <= r_n_468__12_;
      r_468__11_ <= r_n_468__11_;
      r_468__10_ <= r_n_468__10_;
      r_468__9_ <= r_n_468__9_;
      r_468__8_ <= r_n_468__8_;
      r_468__7_ <= r_n_468__7_;
      r_468__6_ <= r_n_468__6_;
      r_468__5_ <= r_n_468__5_;
      r_468__4_ <= r_n_468__4_;
      r_468__3_ <= r_n_468__3_;
      r_468__2_ <= r_n_468__2_;
      r_468__1_ <= r_n_468__1_;
      r_468__0_ <= r_n_468__0_;
    end 
    if(N4053) begin
      r_469__63_ <= r_n_469__63_;
      r_469__62_ <= r_n_469__62_;
      r_469__61_ <= r_n_469__61_;
      r_469__60_ <= r_n_469__60_;
      r_469__59_ <= r_n_469__59_;
      r_469__58_ <= r_n_469__58_;
      r_469__57_ <= r_n_469__57_;
      r_469__56_ <= r_n_469__56_;
      r_469__55_ <= r_n_469__55_;
      r_469__54_ <= r_n_469__54_;
      r_469__53_ <= r_n_469__53_;
      r_469__52_ <= r_n_469__52_;
      r_469__51_ <= r_n_469__51_;
      r_469__50_ <= r_n_469__50_;
      r_469__49_ <= r_n_469__49_;
      r_469__48_ <= r_n_469__48_;
      r_469__47_ <= r_n_469__47_;
      r_469__46_ <= r_n_469__46_;
      r_469__45_ <= r_n_469__45_;
      r_469__44_ <= r_n_469__44_;
      r_469__43_ <= r_n_469__43_;
      r_469__42_ <= r_n_469__42_;
      r_469__41_ <= r_n_469__41_;
      r_469__40_ <= r_n_469__40_;
      r_469__39_ <= r_n_469__39_;
      r_469__38_ <= r_n_469__38_;
      r_469__37_ <= r_n_469__37_;
      r_469__36_ <= r_n_469__36_;
      r_469__35_ <= r_n_469__35_;
      r_469__34_ <= r_n_469__34_;
      r_469__33_ <= r_n_469__33_;
      r_469__32_ <= r_n_469__32_;
      r_469__31_ <= r_n_469__31_;
      r_469__30_ <= r_n_469__30_;
      r_469__29_ <= r_n_469__29_;
      r_469__28_ <= r_n_469__28_;
      r_469__27_ <= r_n_469__27_;
      r_469__26_ <= r_n_469__26_;
      r_469__25_ <= r_n_469__25_;
      r_469__24_ <= r_n_469__24_;
      r_469__23_ <= r_n_469__23_;
      r_469__22_ <= r_n_469__22_;
      r_469__21_ <= r_n_469__21_;
      r_469__20_ <= r_n_469__20_;
      r_469__19_ <= r_n_469__19_;
      r_469__18_ <= r_n_469__18_;
      r_469__17_ <= r_n_469__17_;
      r_469__16_ <= r_n_469__16_;
      r_469__15_ <= r_n_469__15_;
      r_469__14_ <= r_n_469__14_;
      r_469__13_ <= r_n_469__13_;
      r_469__12_ <= r_n_469__12_;
      r_469__11_ <= r_n_469__11_;
      r_469__10_ <= r_n_469__10_;
      r_469__9_ <= r_n_469__9_;
      r_469__8_ <= r_n_469__8_;
      r_469__7_ <= r_n_469__7_;
      r_469__6_ <= r_n_469__6_;
      r_469__5_ <= r_n_469__5_;
      r_469__4_ <= r_n_469__4_;
      r_469__3_ <= r_n_469__3_;
      r_469__2_ <= r_n_469__2_;
      r_469__1_ <= r_n_469__1_;
      r_469__0_ <= r_n_469__0_;
    end 
    if(N4054) begin
      r_470__63_ <= r_n_470__63_;
      r_470__62_ <= r_n_470__62_;
      r_470__61_ <= r_n_470__61_;
      r_470__60_ <= r_n_470__60_;
      r_470__59_ <= r_n_470__59_;
      r_470__58_ <= r_n_470__58_;
      r_470__57_ <= r_n_470__57_;
      r_470__56_ <= r_n_470__56_;
      r_470__55_ <= r_n_470__55_;
      r_470__54_ <= r_n_470__54_;
      r_470__53_ <= r_n_470__53_;
      r_470__52_ <= r_n_470__52_;
      r_470__51_ <= r_n_470__51_;
      r_470__50_ <= r_n_470__50_;
      r_470__49_ <= r_n_470__49_;
      r_470__48_ <= r_n_470__48_;
      r_470__47_ <= r_n_470__47_;
      r_470__46_ <= r_n_470__46_;
      r_470__45_ <= r_n_470__45_;
      r_470__44_ <= r_n_470__44_;
      r_470__43_ <= r_n_470__43_;
      r_470__42_ <= r_n_470__42_;
      r_470__41_ <= r_n_470__41_;
      r_470__40_ <= r_n_470__40_;
      r_470__39_ <= r_n_470__39_;
      r_470__38_ <= r_n_470__38_;
      r_470__37_ <= r_n_470__37_;
      r_470__36_ <= r_n_470__36_;
      r_470__35_ <= r_n_470__35_;
      r_470__34_ <= r_n_470__34_;
      r_470__33_ <= r_n_470__33_;
      r_470__32_ <= r_n_470__32_;
      r_470__31_ <= r_n_470__31_;
      r_470__30_ <= r_n_470__30_;
      r_470__29_ <= r_n_470__29_;
      r_470__28_ <= r_n_470__28_;
      r_470__27_ <= r_n_470__27_;
      r_470__26_ <= r_n_470__26_;
      r_470__25_ <= r_n_470__25_;
      r_470__24_ <= r_n_470__24_;
      r_470__23_ <= r_n_470__23_;
      r_470__22_ <= r_n_470__22_;
      r_470__21_ <= r_n_470__21_;
      r_470__20_ <= r_n_470__20_;
      r_470__19_ <= r_n_470__19_;
      r_470__18_ <= r_n_470__18_;
      r_470__17_ <= r_n_470__17_;
      r_470__16_ <= r_n_470__16_;
      r_470__15_ <= r_n_470__15_;
      r_470__14_ <= r_n_470__14_;
      r_470__13_ <= r_n_470__13_;
      r_470__12_ <= r_n_470__12_;
      r_470__11_ <= r_n_470__11_;
      r_470__10_ <= r_n_470__10_;
      r_470__9_ <= r_n_470__9_;
      r_470__8_ <= r_n_470__8_;
      r_470__7_ <= r_n_470__7_;
      r_470__6_ <= r_n_470__6_;
      r_470__5_ <= r_n_470__5_;
      r_470__4_ <= r_n_470__4_;
      r_470__3_ <= r_n_470__3_;
      r_470__2_ <= r_n_470__2_;
      r_470__1_ <= r_n_470__1_;
      r_470__0_ <= r_n_470__0_;
    end 
    if(N4055) begin
      r_471__63_ <= r_n_471__63_;
      r_471__62_ <= r_n_471__62_;
      r_471__61_ <= r_n_471__61_;
      r_471__60_ <= r_n_471__60_;
      r_471__59_ <= r_n_471__59_;
      r_471__58_ <= r_n_471__58_;
      r_471__57_ <= r_n_471__57_;
      r_471__56_ <= r_n_471__56_;
      r_471__55_ <= r_n_471__55_;
      r_471__54_ <= r_n_471__54_;
      r_471__53_ <= r_n_471__53_;
      r_471__52_ <= r_n_471__52_;
      r_471__51_ <= r_n_471__51_;
      r_471__50_ <= r_n_471__50_;
      r_471__49_ <= r_n_471__49_;
      r_471__48_ <= r_n_471__48_;
      r_471__47_ <= r_n_471__47_;
      r_471__46_ <= r_n_471__46_;
      r_471__45_ <= r_n_471__45_;
      r_471__44_ <= r_n_471__44_;
      r_471__43_ <= r_n_471__43_;
      r_471__42_ <= r_n_471__42_;
      r_471__41_ <= r_n_471__41_;
      r_471__40_ <= r_n_471__40_;
      r_471__39_ <= r_n_471__39_;
      r_471__38_ <= r_n_471__38_;
      r_471__37_ <= r_n_471__37_;
      r_471__36_ <= r_n_471__36_;
      r_471__35_ <= r_n_471__35_;
      r_471__34_ <= r_n_471__34_;
      r_471__33_ <= r_n_471__33_;
      r_471__32_ <= r_n_471__32_;
      r_471__31_ <= r_n_471__31_;
      r_471__30_ <= r_n_471__30_;
      r_471__29_ <= r_n_471__29_;
      r_471__28_ <= r_n_471__28_;
      r_471__27_ <= r_n_471__27_;
      r_471__26_ <= r_n_471__26_;
      r_471__25_ <= r_n_471__25_;
      r_471__24_ <= r_n_471__24_;
      r_471__23_ <= r_n_471__23_;
      r_471__22_ <= r_n_471__22_;
      r_471__21_ <= r_n_471__21_;
      r_471__20_ <= r_n_471__20_;
      r_471__19_ <= r_n_471__19_;
      r_471__18_ <= r_n_471__18_;
      r_471__17_ <= r_n_471__17_;
      r_471__16_ <= r_n_471__16_;
      r_471__15_ <= r_n_471__15_;
      r_471__14_ <= r_n_471__14_;
      r_471__13_ <= r_n_471__13_;
      r_471__12_ <= r_n_471__12_;
      r_471__11_ <= r_n_471__11_;
      r_471__10_ <= r_n_471__10_;
      r_471__9_ <= r_n_471__9_;
      r_471__8_ <= r_n_471__8_;
      r_471__7_ <= r_n_471__7_;
      r_471__6_ <= r_n_471__6_;
      r_471__5_ <= r_n_471__5_;
      r_471__4_ <= r_n_471__4_;
      r_471__3_ <= r_n_471__3_;
      r_471__2_ <= r_n_471__2_;
      r_471__1_ <= r_n_471__1_;
      r_471__0_ <= r_n_471__0_;
    end 
    if(N4056) begin
      r_472__63_ <= r_n_472__63_;
      r_472__62_ <= r_n_472__62_;
      r_472__61_ <= r_n_472__61_;
      r_472__60_ <= r_n_472__60_;
      r_472__59_ <= r_n_472__59_;
      r_472__58_ <= r_n_472__58_;
      r_472__57_ <= r_n_472__57_;
      r_472__56_ <= r_n_472__56_;
      r_472__55_ <= r_n_472__55_;
      r_472__54_ <= r_n_472__54_;
      r_472__53_ <= r_n_472__53_;
      r_472__52_ <= r_n_472__52_;
      r_472__51_ <= r_n_472__51_;
      r_472__50_ <= r_n_472__50_;
      r_472__49_ <= r_n_472__49_;
      r_472__48_ <= r_n_472__48_;
      r_472__47_ <= r_n_472__47_;
      r_472__46_ <= r_n_472__46_;
      r_472__45_ <= r_n_472__45_;
      r_472__44_ <= r_n_472__44_;
      r_472__43_ <= r_n_472__43_;
      r_472__42_ <= r_n_472__42_;
      r_472__41_ <= r_n_472__41_;
      r_472__40_ <= r_n_472__40_;
      r_472__39_ <= r_n_472__39_;
      r_472__38_ <= r_n_472__38_;
      r_472__37_ <= r_n_472__37_;
      r_472__36_ <= r_n_472__36_;
      r_472__35_ <= r_n_472__35_;
      r_472__34_ <= r_n_472__34_;
      r_472__33_ <= r_n_472__33_;
      r_472__32_ <= r_n_472__32_;
      r_472__31_ <= r_n_472__31_;
      r_472__30_ <= r_n_472__30_;
      r_472__29_ <= r_n_472__29_;
      r_472__28_ <= r_n_472__28_;
      r_472__27_ <= r_n_472__27_;
      r_472__26_ <= r_n_472__26_;
      r_472__25_ <= r_n_472__25_;
      r_472__24_ <= r_n_472__24_;
      r_472__23_ <= r_n_472__23_;
      r_472__22_ <= r_n_472__22_;
      r_472__21_ <= r_n_472__21_;
      r_472__20_ <= r_n_472__20_;
      r_472__19_ <= r_n_472__19_;
      r_472__18_ <= r_n_472__18_;
      r_472__17_ <= r_n_472__17_;
      r_472__16_ <= r_n_472__16_;
      r_472__15_ <= r_n_472__15_;
      r_472__14_ <= r_n_472__14_;
      r_472__13_ <= r_n_472__13_;
      r_472__12_ <= r_n_472__12_;
      r_472__11_ <= r_n_472__11_;
      r_472__10_ <= r_n_472__10_;
      r_472__9_ <= r_n_472__9_;
      r_472__8_ <= r_n_472__8_;
      r_472__7_ <= r_n_472__7_;
      r_472__6_ <= r_n_472__6_;
      r_472__5_ <= r_n_472__5_;
      r_472__4_ <= r_n_472__4_;
      r_472__3_ <= r_n_472__3_;
      r_472__2_ <= r_n_472__2_;
      r_472__1_ <= r_n_472__1_;
      r_472__0_ <= r_n_472__0_;
    end 
    if(N4057) begin
      r_473__63_ <= r_n_473__63_;
      r_473__62_ <= r_n_473__62_;
      r_473__61_ <= r_n_473__61_;
      r_473__60_ <= r_n_473__60_;
      r_473__59_ <= r_n_473__59_;
      r_473__58_ <= r_n_473__58_;
      r_473__57_ <= r_n_473__57_;
      r_473__56_ <= r_n_473__56_;
      r_473__55_ <= r_n_473__55_;
      r_473__54_ <= r_n_473__54_;
      r_473__53_ <= r_n_473__53_;
      r_473__52_ <= r_n_473__52_;
      r_473__51_ <= r_n_473__51_;
      r_473__50_ <= r_n_473__50_;
      r_473__49_ <= r_n_473__49_;
      r_473__48_ <= r_n_473__48_;
      r_473__47_ <= r_n_473__47_;
      r_473__46_ <= r_n_473__46_;
      r_473__45_ <= r_n_473__45_;
      r_473__44_ <= r_n_473__44_;
      r_473__43_ <= r_n_473__43_;
      r_473__42_ <= r_n_473__42_;
      r_473__41_ <= r_n_473__41_;
      r_473__40_ <= r_n_473__40_;
      r_473__39_ <= r_n_473__39_;
      r_473__38_ <= r_n_473__38_;
      r_473__37_ <= r_n_473__37_;
      r_473__36_ <= r_n_473__36_;
      r_473__35_ <= r_n_473__35_;
      r_473__34_ <= r_n_473__34_;
      r_473__33_ <= r_n_473__33_;
      r_473__32_ <= r_n_473__32_;
      r_473__31_ <= r_n_473__31_;
      r_473__30_ <= r_n_473__30_;
      r_473__29_ <= r_n_473__29_;
      r_473__28_ <= r_n_473__28_;
      r_473__27_ <= r_n_473__27_;
      r_473__26_ <= r_n_473__26_;
      r_473__25_ <= r_n_473__25_;
      r_473__24_ <= r_n_473__24_;
      r_473__23_ <= r_n_473__23_;
      r_473__22_ <= r_n_473__22_;
      r_473__21_ <= r_n_473__21_;
      r_473__20_ <= r_n_473__20_;
      r_473__19_ <= r_n_473__19_;
      r_473__18_ <= r_n_473__18_;
      r_473__17_ <= r_n_473__17_;
      r_473__16_ <= r_n_473__16_;
      r_473__15_ <= r_n_473__15_;
      r_473__14_ <= r_n_473__14_;
      r_473__13_ <= r_n_473__13_;
      r_473__12_ <= r_n_473__12_;
      r_473__11_ <= r_n_473__11_;
      r_473__10_ <= r_n_473__10_;
      r_473__9_ <= r_n_473__9_;
      r_473__8_ <= r_n_473__8_;
      r_473__7_ <= r_n_473__7_;
      r_473__6_ <= r_n_473__6_;
      r_473__5_ <= r_n_473__5_;
      r_473__4_ <= r_n_473__4_;
      r_473__3_ <= r_n_473__3_;
      r_473__2_ <= r_n_473__2_;
      r_473__1_ <= r_n_473__1_;
      r_473__0_ <= r_n_473__0_;
    end 
    if(N4058) begin
      r_474__63_ <= r_n_474__63_;
      r_474__62_ <= r_n_474__62_;
      r_474__61_ <= r_n_474__61_;
      r_474__60_ <= r_n_474__60_;
      r_474__59_ <= r_n_474__59_;
      r_474__58_ <= r_n_474__58_;
      r_474__57_ <= r_n_474__57_;
      r_474__56_ <= r_n_474__56_;
      r_474__55_ <= r_n_474__55_;
      r_474__54_ <= r_n_474__54_;
      r_474__53_ <= r_n_474__53_;
      r_474__52_ <= r_n_474__52_;
      r_474__51_ <= r_n_474__51_;
      r_474__50_ <= r_n_474__50_;
      r_474__49_ <= r_n_474__49_;
      r_474__48_ <= r_n_474__48_;
      r_474__47_ <= r_n_474__47_;
      r_474__46_ <= r_n_474__46_;
      r_474__45_ <= r_n_474__45_;
      r_474__44_ <= r_n_474__44_;
      r_474__43_ <= r_n_474__43_;
      r_474__42_ <= r_n_474__42_;
      r_474__41_ <= r_n_474__41_;
      r_474__40_ <= r_n_474__40_;
      r_474__39_ <= r_n_474__39_;
      r_474__38_ <= r_n_474__38_;
      r_474__37_ <= r_n_474__37_;
      r_474__36_ <= r_n_474__36_;
      r_474__35_ <= r_n_474__35_;
      r_474__34_ <= r_n_474__34_;
      r_474__33_ <= r_n_474__33_;
      r_474__32_ <= r_n_474__32_;
      r_474__31_ <= r_n_474__31_;
      r_474__30_ <= r_n_474__30_;
      r_474__29_ <= r_n_474__29_;
      r_474__28_ <= r_n_474__28_;
      r_474__27_ <= r_n_474__27_;
      r_474__26_ <= r_n_474__26_;
      r_474__25_ <= r_n_474__25_;
      r_474__24_ <= r_n_474__24_;
      r_474__23_ <= r_n_474__23_;
      r_474__22_ <= r_n_474__22_;
      r_474__21_ <= r_n_474__21_;
      r_474__20_ <= r_n_474__20_;
      r_474__19_ <= r_n_474__19_;
      r_474__18_ <= r_n_474__18_;
      r_474__17_ <= r_n_474__17_;
      r_474__16_ <= r_n_474__16_;
      r_474__15_ <= r_n_474__15_;
      r_474__14_ <= r_n_474__14_;
      r_474__13_ <= r_n_474__13_;
      r_474__12_ <= r_n_474__12_;
      r_474__11_ <= r_n_474__11_;
      r_474__10_ <= r_n_474__10_;
      r_474__9_ <= r_n_474__9_;
      r_474__8_ <= r_n_474__8_;
      r_474__7_ <= r_n_474__7_;
      r_474__6_ <= r_n_474__6_;
      r_474__5_ <= r_n_474__5_;
      r_474__4_ <= r_n_474__4_;
      r_474__3_ <= r_n_474__3_;
      r_474__2_ <= r_n_474__2_;
      r_474__1_ <= r_n_474__1_;
      r_474__0_ <= r_n_474__0_;
    end 
    if(N4059) begin
      r_475__63_ <= r_n_475__63_;
      r_475__62_ <= r_n_475__62_;
      r_475__61_ <= r_n_475__61_;
      r_475__60_ <= r_n_475__60_;
      r_475__59_ <= r_n_475__59_;
      r_475__58_ <= r_n_475__58_;
      r_475__57_ <= r_n_475__57_;
      r_475__56_ <= r_n_475__56_;
      r_475__55_ <= r_n_475__55_;
      r_475__54_ <= r_n_475__54_;
      r_475__53_ <= r_n_475__53_;
      r_475__52_ <= r_n_475__52_;
      r_475__51_ <= r_n_475__51_;
      r_475__50_ <= r_n_475__50_;
      r_475__49_ <= r_n_475__49_;
      r_475__48_ <= r_n_475__48_;
      r_475__47_ <= r_n_475__47_;
      r_475__46_ <= r_n_475__46_;
      r_475__45_ <= r_n_475__45_;
      r_475__44_ <= r_n_475__44_;
      r_475__43_ <= r_n_475__43_;
      r_475__42_ <= r_n_475__42_;
      r_475__41_ <= r_n_475__41_;
      r_475__40_ <= r_n_475__40_;
      r_475__39_ <= r_n_475__39_;
      r_475__38_ <= r_n_475__38_;
      r_475__37_ <= r_n_475__37_;
      r_475__36_ <= r_n_475__36_;
      r_475__35_ <= r_n_475__35_;
      r_475__34_ <= r_n_475__34_;
      r_475__33_ <= r_n_475__33_;
      r_475__32_ <= r_n_475__32_;
      r_475__31_ <= r_n_475__31_;
      r_475__30_ <= r_n_475__30_;
      r_475__29_ <= r_n_475__29_;
      r_475__28_ <= r_n_475__28_;
      r_475__27_ <= r_n_475__27_;
      r_475__26_ <= r_n_475__26_;
      r_475__25_ <= r_n_475__25_;
      r_475__24_ <= r_n_475__24_;
      r_475__23_ <= r_n_475__23_;
      r_475__22_ <= r_n_475__22_;
      r_475__21_ <= r_n_475__21_;
      r_475__20_ <= r_n_475__20_;
      r_475__19_ <= r_n_475__19_;
      r_475__18_ <= r_n_475__18_;
      r_475__17_ <= r_n_475__17_;
      r_475__16_ <= r_n_475__16_;
      r_475__15_ <= r_n_475__15_;
      r_475__14_ <= r_n_475__14_;
      r_475__13_ <= r_n_475__13_;
      r_475__12_ <= r_n_475__12_;
      r_475__11_ <= r_n_475__11_;
      r_475__10_ <= r_n_475__10_;
      r_475__9_ <= r_n_475__9_;
      r_475__8_ <= r_n_475__8_;
      r_475__7_ <= r_n_475__7_;
      r_475__6_ <= r_n_475__6_;
      r_475__5_ <= r_n_475__5_;
      r_475__4_ <= r_n_475__4_;
      r_475__3_ <= r_n_475__3_;
      r_475__2_ <= r_n_475__2_;
      r_475__1_ <= r_n_475__1_;
      r_475__0_ <= r_n_475__0_;
    end 
    if(N4060) begin
      r_476__63_ <= r_n_476__63_;
      r_476__62_ <= r_n_476__62_;
      r_476__61_ <= r_n_476__61_;
      r_476__60_ <= r_n_476__60_;
      r_476__59_ <= r_n_476__59_;
      r_476__58_ <= r_n_476__58_;
      r_476__57_ <= r_n_476__57_;
      r_476__56_ <= r_n_476__56_;
      r_476__55_ <= r_n_476__55_;
      r_476__54_ <= r_n_476__54_;
      r_476__53_ <= r_n_476__53_;
      r_476__52_ <= r_n_476__52_;
      r_476__51_ <= r_n_476__51_;
      r_476__50_ <= r_n_476__50_;
      r_476__49_ <= r_n_476__49_;
      r_476__48_ <= r_n_476__48_;
      r_476__47_ <= r_n_476__47_;
      r_476__46_ <= r_n_476__46_;
      r_476__45_ <= r_n_476__45_;
      r_476__44_ <= r_n_476__44_;
      r_476__43_ <= r_n_476__43_;
      r_476__42_ <= r_n_476__42_;
      r_476__41_ <= r_n_476__41_;
      r_476__40_ <= r_n_476__40_;
      r_476__39_ <= r_n_476__39_;
      r_476__38_ <= r_n_476__38_;
      r_476__37_ <= r_n_476__37_;
      r_476__36_ <= r_n_476__36_;
      r_476__35_ <= r_n_476__35_;
      r_476__34_ <= r_n_476__34_;
      r_476__33_ <= r_n_476__33_;
      r_476__32_ <= r_n_476__32_;
      r_476__31_ <= r_n_476__31_;
      r_476__30_ <= r_n_476__30_;
      r_476__29_ <= r_n_476__29_;
      r_476__28_ <= r_n_476__28_;
      r_476__27_ <= r_n_476__27_;
      r_476__26_ <= r_n_476__26_;
      r_476__25_ <= r_n_476__25_;
      r_476__24_ <= r_n_476__24_;
      r_476__23_ <= r_n_476__23_;
      r_476__22_ <= r_n_476__22_;
      r_476__21_ <= r_n_476__21_;
      r_476__20_ <= r_n_476__20_;
      r_476__19_ <= r_n_476__19_;
      r_476__18_ <= r_n_476__18_;
      r_476__17_ <= r_n_476__17_;
      r_476__16_ <= r_n_476__16_;
      r_476__15_ <= r_n_476__15_;
      r_476__14_ <= r_n_476__14_;
      r_476__13_ <= r_n_476__13_;
      r_476__12_ <= r_n_476__12_;
      r_476__11_ <= r_n_476__11_;
      r_476__10_ <= r_n_476__10_;
      r_476__9_ <= r_n_476__9_;
      r_476__8_ <= r_n_476__8_;
      r_476__7_ <= r_n_476__7_;
      r_476__6_ <= r_n_476__6_;
      r_476__5_ <= r_n_476__5_;
      r_476__4_ <= r_n_476__4_;
      r_476__3_ <= r_n_476__3_;
      r_476__2_ <= r_n_476__2_;
      r_476__1_ <= r_n_476__1_;
      r_476__0_ <= r_n_476__0_;
    end 
    if(N4061) begin
      r_477__63_ <= r_n_477__63_;
      r_477__62_ <= r_n_477__62_;
      r_477__61_ <= r_n_477__61_;
      r_477__60_ <= r_n_477__60_;
      r_477__59_ <= r_n_477__59_;
      r_477__58_ <= r_n_477__58_;
      r_477__57_ <= r_n_477__57_;
      r_477__56_ <= r_n_477__56_;
      r_477__55_ <= r_n_477__55_;
      r_477__54_ <= r_n_477__54_;
      r_477__53_ <= r_n_477__53_;
      r_477__52_ <= r_n_477__52_;
      r_477__51_ <= r_n_477__51_;
      r_477__50_ <= r_n_477__50_;
      r_477__49_ <= r_n_477__49_;
      r_477__48_ <= r_n_477__48_;
      r_477__47_ <= r_n_477__47_;
      r_477__46_ <= r_n_477__46_;
      r_477__45_ <= r_n_477__45_;
      r_477__44_ <= r_n_477__44_;
      r_477__43_ <= r_n_477__43_;
      r_477__42_ <= r_n_477__42_;
      r_477__41_ <= r_n_477__41_;
      r_477__40_ <= r_n_477__40_;
      r_477__39_ <= r_n_477__39_;
      r_477__38_ <= r_n_477__38_;
      r_477__37_ <= r_n_477__37_;
      r_477__36_ <= r_n_477__36_;
      r_477__35_ <= r_n_477__35_;
      r_477__34_ <= r_n_477__34_;
      r_477__33_ <= r_n_477__33_;
      r_477__32_ <= r_n_477__32_;
      r_477__31_ <= r_n_477__31_;
      r_477__30_ <= r_n_477__30_;
      r_477__29_ <= r_n_477__29_;
      r_477__28_ <= r_n_477__28_;
      r_477__27_ <= r_n_477__27_;
      r_477__26_ <= r_n_477__26_;
      r_477__25_ <= r_n_477__25_;
      r_477__24_ <= r_n_477__24_;
      r_477__23_ <= r_n_477__23_;
      r_477__22_ <= r_n_477__22_;
      r_477__21_ <= r_n_477__21_;
      r_477__20_ <= r_n_477__20_;
      r_477__19_ <= r_n_477__19_;
      r_477__18_ <= r_n_477__18_;
      r_477__17_ <= r_n_477__17_;
      r_477__16_ <= r_n_477__16_;
      r_477__15_ <= r_n_477__15_;
      r_477__14_ <= r_n_477__14_;
      r_477__13_ <= r_n_477__13_;
      r_477__12_ <= r_n_477__12_;
      r_477__11_ <= r_n_477__11_;
      r_477__10_ <= r_n_477__10_;
      r_477__9_ <= r_n_477__9_;
      r_477__8_ <= r_n_477__8_;
      r_477__7_ <= r_n_477__7_;
      r_477__6_ <= r_n_477__6_;
      r_477__5_ <= r_n_477__5_;
      r_477__4_ <= r_n_477__4_;
      r_477__3_ <= r_n_477__3_;
      r_477__2_ <= r_n_477__2_;
      r_477__1_ <= r_n_477__1_;
      r_477__0_ <= r_n_477__0_;
    end 
    if(N4062) begin
      r_478__63_ <= r_n_478__63_;
      r_478__62_ <= r_n_478__62_;
      r_478__61_ <= r_n_478__61_;
      r_478__60_ <= r_n_478__60_;
      r_478__59_ <= r_n_478__59_;
      r_478__58_ <= r_n_478__58_;
      r_478__57_ <= r_n_478__57_;
      r_478__56_ <= r_n_478__56_;
      r_478__55_ <= r_n_478__55_;
      r_478__54_ <= r_n_478__54_;
      r_478__53_ <= r_n_478__53_;
      r_478__52_ <= r_n_478__52_;
      r_478__51_ <= r_n_478__51_;
      r_478__50_ <= r_n_478__50_;
      r_478__49_ <= r_n_478__49_;
      r_478__48_ <= r_n_478__48_;
      r_478__47_ <= r_n_478__47_;
      r_478__46_ <= r_n_478__46_;
      r_478__45_ <= r_n_478__45_;
      r_478__44_ <= r_n_478__44_;
      r_478__43_ <= r_n_478__43_;
      r_478__42_ <= r_n_478__42_;
      r_478__41_ <= r_n_478__41_;
      r_478__40_ <= r_n_478__40_;
      r_478__39_ <= r_n_478__39_;
      r_478__38_ <= r_n_478__38_;
      r_478__37_ <= r_n_478__37_;
      r_478__36_ <= r_n_478__36_;
      r_478__35_ <= r_n_478__35_;
      r_478__34_ <= r_n_478__34_;
      r_478__33_ <= r_n_478__33_;
      r_478__32_ <= r_n_478__32_;
      r_478__31_ <= r_n_478__31_;
      r_478__30_ <= r_n_478__30_;
      r_478__29_ <= r_n_478__29_;
      r_478__28_ <= r_n_478__28_;
      r_478__27_ <= r_n_478__27_;
      r_478__26_ <= r_n_478__26_;
      r_478__25_ <= r_n_478__25_;
      r_478__24_ <= r_n_478__24_;
      r_478__23_ <= r_n_478__23_;
      r_478__22_ <= r_n_478__22_;
      r_478__21_ <= r_n_478__21_;
      r_478__20_ <= r_n_478__20_;
      r_478__19_ <= r_n_478__19_;
      r_478__18_ <= r_n_478__18_;
      r_478__17_ <= r_n_478__17_;
      r_478__16_ <= r_n_478__16_;
      r_478__15_ <= r_n_478__15_;
      r_478__14_ <= r_n_478__14_;
      r_478__13_ <= r_n_478__13_;
      r_478__12_ <= r_n_478__12_;
      r_478__11_ <= r_n_478__11_;
      r_478__10_ <= r_n_478__10_;
      r_478__9_ <= r_n_478__9_;
      r_478__8_ <= r_n_478__8_;
      r_478__7_ <= r_n_478__7_;
      r_478__6_ <= r_n_478__6_;
      r_478__5_ <= r_n_478__5_;
      r_478__4_ <= r_n_478__4_;
      r_478__3_ <= r_n_478__3_;
      r_478__2_ <= r_n_478__2_;
      r_478__1_ <= r_n_478__1_;
      r_478__0_ <= r_n_478__0_;
    end 
    if(N4063) begin
      r_479__63_ <= r_n_479__63_;
      r_479__62_ <= r_n_479__62_;
      r_479__61_ <= r_n_479__61_;
      r_479__60_ <= r_n_479__60_;
      r_479__59_ <= r_n_479__59_;
      r_479__58_ <= r_n_479__58_;
      r_479__57_ <= r_n_479__57_;
      r_479__56_ <= r_n_479__56_;
      r_479__55_ <= r_n_479__55_;
      r_479__54_ <= r_n_479__54_;
      r_479__53_ <= r_n_479__53_;
      r_479__52_ <= r_n_479__52_;
      r_479__51_ <= r_n_479__51_;
      r_479__50_ <= r_n_479__50_;
      r_479__49_ <= r_n_479__49_;
      r_479__48_ <= r_n_479__48_;
      r_479__47_ <= r_n_479__47_;
      r_479__46_ <= r_n_479__46_;
      r_479__45_ <= r_n_479__45_;
      r_479__44_ <= r_n_479__44_;
      r_479__43_ <= r_n_479__43_;
      r_479__42_ <= r_n_479__42_;
      r_479__41_ <= r_n_479__41_;
      r_479__40_ <= r_n_479__40_;
      r_479__39_ <= r_n_479__39_;
      r_479__38_ <= r_n_479__38_;
      r_479__37_ <= r_n_479__37_;
      r_479__36_ <= r_n_479__36_;
      r_479__35_ <= r_n_479__35_;
      r_479__34_ <= r_n_479__34_;
      r_479__33_ <= r_n_479__33_;
      r_479__32_ <= r_n_479__32_;
      r_479__31_ <= r_n_479__31_;
      r_479__30_ <= r_n_479__30_;
      r_479__29_ <= r_n_479__29_;
      r_479__28_ <= r_n_479__28_;
      r_479__27_ <= r_n_479__27_;
      r_479__26_ <= r_n_479__26_;
      r_479__25_ <= r_n_479__25_;
      r_479__24_ <= r_n_479__24_;
      r_479__23_ <= r_n_479__23_;
      r_479__22_ <= r_n_479__22_;
      r_479__21_ <= r_n_479__21_;
      r_479__20_ <= r_n_479__20_;
      r_479__19_ <= r_n_479__19_;
      r_479__18_ <= r_n_479__18_;
      r_479__17_ <= r_n_479__17_;
      r_479__16_ <= r_n_479__16_;
      r_479__15_ <= r_n_479__15_;
      r_479__14_ <= r_n_479__14_;
      r_479__13_ <= r_n_479__13_;
      r_479__12_ <= r_n_479__12_;
      r_479__11_ <= r_n_479__11_;
      r_479__10_ <= r_n_479__10_;
      r_479__9_ <= r_n_479__9_;
      r_479__8_ <= r_n_479__8_;
      r_479__7_ <= r_n_479__7_;
      r_479__6_ <= r_n_479__6_;
      r_479__5_ <= r_n_479__5_;
      r_479__4_ <= r_n_479__4_;
      r_479__3_ <= r_n_479__3_;
      r_479__2_ <= r_n_479__2_;
      r_479__1_ <= r_n_479__1_;
      r_479__0_ <= r_n_479__0_;
    end 
    if(N4064) begin
      r_480__63_ <= r_n_480__63_;
      r_480__62_ <= r_n_480__62_;
      r_480__61_ <= r_n_480__61_;
      r_480__60_ <= r_n_480__60_;
      r_480__59_ <= r_n_480__59_;
      r_480__58_ <= r_n_480__58_;
      r_480__57_ <= r_n_480__57_;
      r_480__56_ <= r_n_480__56_;
      r_480__55_ <= r_n_480__55_;
      r_480__54_ <= r_n_480__54_;
      r_480__53_ <= r_n_480__53_;
      r_480__52_ <= r_n_480__52_;
      r_480__51_ <= r_n_480__51_;
      r_480__50_ <= r_n_480__50_;
      r_480__49_ <= r_n_480__49_;
      r_480__48_ <= r_n_480__48_;
      r_480__47_ <= r_n_480__47_;
      r_480__46_ <= r_n_480__46_;
      r_480__45_ <= r_n_480__45_;
      r_480__44_ <= r_n_480__44_;
      r_480__43_ <= r_n_480__43_;
      r_480__42_ <= r_n_480__42_;
      r_480__41_ <= r_n_480__41_;
      r_480__40_ <= r_n_480__40_;
      r_480__39_ <= r_n_480__39_;
      r_480__38_ <= r_n_480__38_;
      r_480__37_ <= r_n_480__37_;
      r_480__36_ <= r_n_480__36_;
      r_480__35_ <= r_n_480__35_;
      r_480__34_ <= r_n_480__34_;
      r_480__33_ <= r_n_480__33_;
      r_480__32_ <= r_n_480__32_;
      r_480__31_ <= r_n_480__31_;
      r_480__30_ <= r_n_480__30_;
      r_480__29_ <= r_n_480__29_;
      r_480__28_ <= r_n_480__28_;
      r_480__27_ <= r_n_480__27_;
      r_480__26_ <= r_n_480__26_;
      r_480__25_ <= r_n_480__25_;
      r_480__24_ <= r_n_480__24_;
      r_480__23_ <= r_n_480__23_;
      r_480__22_ <= r_n_480__22_;
      r_480__21_ <= r_n_480__21_;
      r_480__20_ <= r_n_480__20_;
      r_480__19_ <= r_n_480__19_;
      r_480__18_ <= r_n_480__18_;
      r_480__17_ <= r_n_480__17_;
      r_480__16_ <= r_n_480__16_;
      r_480__15_ <= r_n_480__15_;
      r_480__14_ <= r_n_480__14_;
      r_480__13_ <= r_n_480__13_;
      r_480__12_ <= r_n_480__12_;
      r_480__11_ <= r_n_480__11_;
      r_480__10_ <= r_n_480__10_;
      r_480__9_ <= r_n_480__9_;
      r_480__8_ <= r_n_480__8_;
      r_480__7_ <= r_n_480__7_;
      r_480__6_ <= r_n_480__6_;
      r_480__5_ <= r_n_480__5_;
      r_480__4_ <= r_n_480__4_;
      r_480__3_ <= r_n_480__3_;
      r_480__2_ <= r_n_480__2_;
      r_480__1_ <= r_n_480__1_;
      r_480__0_ <= r_n_480__0_;
    end 
    if(N4065) begin
      r_481__63_ <= r_n_481__63_;
      r_481__62_ <= r_n_481__62_;
      r_481__61_ <= r_n_481__61_;
      r_481__60_ <= r_n_481__60_;
      r_481__59_ <= r_n_481__59_;
      r_481__58_ <= r_n_481__58_;
      r_481__57_ <= r_n_481__57_;
      r_481__56_ <= r_n_481__56_;
      r_481__55_ <= r_n_481__55_;
      r_481__54_ <= r_n_481__54_;
      r_481__53_ <= r_n_481__53_;
      r_481__52_ <= r_n_481__52_;
      r_481__51_ <= r_n_481__51_;
      r_481__50_ <= r_n_481__50_;
      r_481__49_ <= r_n_481__49_;
      r_481__48_ <= r_n_481__48_;
      r_481__47_ <= r_n_481__47_;
      r_481__46_ <= r_n_481__46_;
      r_481__45_ <= r_n_481__45_;
      r_481__44_ <= r_n_481__44_;
      r_481__43_ <= r_n_481__43_;
      r_481__42_ <= r_n_481__42_;
      r_481__41_ <= r_n_481__41_;
      r_481__40_ <= r_n_481__40_;
      r_481__39_ <= r_n_481__39_;
      r_481__38_ <= r_n_481__38_;
      r_481__37_ <= r_n_481__37_;
      r_481__36_ <= r_n_481__36_;
      r_481__35_ <= r_n_481__35_;
      r_481__34_ <= r_n_481__34_;
      r_481__33_ <= r_n_481__33_;
      r_481__32_ <= r_n_481__32_;
      r_481__31_ <= r_n_481__31_;
      r_481__30_ <= r_n_481__30_;
      r_481__29_ <= r_n_481__29_;
      r_481__28_ <= r_n_481__28_;
      r_481__27_ <= r_n_481__27_;
      r_481__26_ <= r_n_481__26_;
      r_481__25_ <= r_n_481__25_;
      r_481__24_ <= r_n_481__24_;
      r_481__23_ <= r_n_481__23_;
      r_481__22_ <= r_n_481__22_;
      r_481__21_ <= r_n_481__21_;
      r_481__20_ <= r_n_481__20_;
      r_481__19_ <= r_n_481__19_;
      r_481__18_ <= r_n_481__18_;
      r_481__17_ <= r_n_481__17_;
      r_481__16_ <= r_n_481__16_;
      r_481__15_ <= r_n_481__15_;
      r_481__14_ <= r_n_481__14_;
      r_481__13_ <= r_n_481__13_;
      r_481__12_ <= r_n_481__12_;
      r_481__11_ <= r_n_481__11_;
      r_481__10_ <= r_n_481__10_;
      r_481__9_ <= r_n_481__9_;
      r_481__8_ <= r_n_481__8_;
      r_481__7_ <= r_n_481__7_;
      r_481__6_ <= r_n_481__6_;
      r_481__5_ <= r_n_481__5_;
      r_481__4_ <= r_n_481__4_;
      r_481__3_ <= r_n_481__3_;
      r_481__2_ <= r_n_481__2_;
      r_481__1_ <= r_n_481__1_;
      r_481__0_ <= r_n_481__0_;
    end 
    if(N4066) begin
      r_482__63_ <= r_n_482__63_;
      r_482__62_ <= r_n_482__62_;
      r_482__61_ <= r_n_482__61_;
      r_482__60_ <= r_n_482__60_;
      r_482__59_ <= r_n_482__59_;
      r_482__58_ <= r_n_482__58_;
      r_482__57_ <= r_n_482__57_;
      r_482__56_ <= r_n_482__56_;
      r_482__55_ <= r_n_482__55_;
      r_482__54_ <= r_n_482__54_;
      r_482__53_ <= r_n_482__53_;
      r_482__52_ <= r_n_482__52_;
      r_482__51_ <= r_n_482__51_;
      r_482__50_ <= r_n_482__50_;
      r_482__49_ <= r_n_482__49_;
      r_482__48_ <= r_n_482__48_;
      r_482__47_ <= r_n_482__47_;
      r_482__46_ <= r_n_482__46_;
      r_482__45_ <= r_n_482__45_;
      r_482__44_ <= r_n_482__44_;
      r_482__43_ <= r_n_482__43_;
      r_482__42_ <= r_n_482__42_;
      r_482__41_ <= r_n_482__41_;
      r_482__40_ <= r_n_482__40_;
      r_482__39_ <= r_n_482__39_;
      r_482__38_ <= r_n_482__38_;
      r_482__37_ <= r_n_482__37_;
      r_482__36_ <= r_n_482__36_;
      r_482__35_ <= r_n_482__35_;
      r_482__34_ <= r_n_482__34_;
      r_482__33_ <= r_n_482__33_;
      r_482__32_ <= r_n_482__32_;
      r_482__31_ <= r_n_482__31_;
      r_482__30_ <= r_n_482__30_;
      r_482__29_ <= r_n_482__29_;
      r_482__28_ <= r_n_482__28_;
      r_482__27_ <= r_n_482__27_;
      r_482__26_ <= r_n_482__26_;
      r_482__25_ <= r_n_482__25_;
      r_482__24_ <= r_n_482__24_;
      r_482__23_ <= r_n_482__23_;
      r_482__22_ <= r_n_482__22_;
      r_482__21_ <= r_n_482__21_;
      r_482__20_ <= r_n_482__20_;
      r_482__19_ <= r_n_482__19_;
      r_482__18_ <= r_n_482__18_;
      r_482__17_ <= r_n_482__17_;
      r_482__16_ <= r_n_482__16_;
      r_482__15_ <= r_n_482__15_;
      r_482__14_ <= r_n_482__14_;
      r_482__13_ <= r_n_482__13_;
      r_482__12_ <= r_n_482__12_;
      r_482__11_ <= r_n_482__11_;
      r_482__10_ <= r_n_482__10_;
      r_482__9_ <= r_n_482__9_;
      r_482__8_ <= r_n_482__8_;
      r_482__7_ <= r_n_482__7_;
      r_482__6_ <= r_n_482__6_;
      r_482__5_ <= r_n_482__5_;
      r_482__4_ <= r_n_482__4_;
      r_482__3_ <= r_n_482__3_;
      r_482__2_ <= r_n_482__2_;
      r_482__1_ <= r_n_482__1_;
      r_482__0_ <= r_n_482__0_;
    end 
    if(N4067) begin
      r_483__63_ <= r_n_483__63_;
      r_483__62_ <= r_n_483__62_;
      r_483__61_ <= r_n_483__61_;
      r_483__60_ <= r_n_483__60_;
      r_483__59_ <= r_n_483__59_;
      r_483__58_ <= r_n_483__58_;
      r_483__57_ <= r_n_483__57_;
      r_483__56_ <= r_n_483__56_;
      r_483__55_ <= r_n_483__55_;
      r_483__54_ <= r_n_483__54_;
      r_483__53_ <= r_n_483__53_;
      r_483__52_ <= r_n_483__52_;
      r_483__51_ <= r_n_483__51_;
      r_483__50_ <= r_n_483__50_;
      r_483__49_ <= r_n_483__49_;
      r_483__48_ <= r_n_483__48_;
      r_483__47_ <= r_n_483__47_;
      r_483__46_ <= r_n_483__46_;
      r_483__45_ <= r_n_483__45_;
      r_483__44_ <= r_n_483__44_;
      r_483__43_ <= r_n_483__43_;
      r_483__42_ <= r_n_483__42_;
      r_483__41_ <= r_n_483__41_;
      r_483__40_ <= r_n_483__40_;
      r_483__39_ <= r_n_483__39_;
      r_483__38_ <= r_n_483__38_;
      r_483__37_ <= r_n_483__37_;
      r_483__36_ <= r_n_483__36_;
      r_483__35_ <= r_n_483__35_;
      r_483__34_ <= r_n_483__34_;
      r_483__33_ <= r_n_483__33_;
      r_483__32_ <= r_n_483__32_;
      r_483__31_ <= r_n_483__31_;
      r_483__30_ <= r_n_483__30_;
      r_483__29_ <= r_n_483__29_;
      r_483__28_ <= r_n_483__28_;
      r_483__27_ <= r_n_483__27_;
      r_483__26_ <= r_n_483__26_;
      r_483__25_ <= r_n_483__25_;
      r_483__24_ <= r_n_483__24_;
      r_483__23_ <= r_n_483__23_;
      r_483__22_ <= r_n_483__22_;
      r_483__21_ <= r_n_483__21_;
      r_483__20_ <= r_n_483__20_;
      r_483__19_ <= r_n_483__19_;
      r_483__18_ <= r_n_483__18_;
      r_483__17_ <= r_n_483__17_;
      r_483__16_ <= r_n_483__16_;
      r_483__15_ <= r_n_483__15_;
      r_483__14_ <= r_n_483__14_;
      r_483__13_ <= r_n_483__13_;
      r_483__12_ <= r_n_483__12_;
      r_483__11_ <= r_n_483__11_;
      r_483__10_ <= r_n_483__10_;
      r_483__9_ <= r_n_483__9_;
      r_483__8_ <= r_n_483__8_;
      r_483__7_ <= r_n_483__7_;
      r_483__6_ <= r_n_483__6_;
      r_483__5_ <= r_n_483__5_;
      r_483__4_ <= r_n_483__4_;
      r_483__3_ <= r_n_483__3_;
      r_483__2_ <= r_n_483__2_;
      r_483__1_ <= r_n_483__1_;
      r_483__0_ <= r_n_483__0_;
    end 
    if(N4068) begin
      r_484__63_ <= r_n_484__63_;
      r_484__62_ <= r_n_484__62_;
      r_484__61_ <= r_n_484__61_;
      r_484__60_ <= r_n_484__60_;
      r_484__59_ <= r_n_484__59_;
      r_484__58_ <= r_n_484__58_;
      r_484__57_ <= r_n_484__57_;
      r_484__56_ <= r_n_484__56_;
      r_484__55_ <= r_n_484__55_;
      r_484__54_ <= r_n_484__54_;
      r_484__53_ <= r_n_484__53_;
      r_484__52_ <= r_n_484__52_;
      r_484__51_ <= r_n_484__51_;
      r_484__50_ <= r_n_484__50_;
      r_484__49_ <= r_n_484__49_;
      r_484__48_ <= r_n_484__48_;
      r_484__47_ <= r_n_484__47_;
      r_484__46_ <= r_n_484__46_;
      r_484__45_ <= r_n_484__45_;
      r_484__44_ <= r_n_484__44_;
      r_484__43_ <= r_n_484__43_;
      r_484__42_ <= r_n_484__42_;
      r_484__41_ <= r_n_484__41_;
      r_484__40_ <= r_n_484__40_;
      r_484__39_ <= r_n_484__39_;
      r_484__38_ <= r_n_484__38_;
      r_484__37_ <= r_n_484__37_;
      r_484__36_ <= r_n_484__36_;
      r_484__35_ <= r_n_484__35_;
      r_484__34_ <= r_n_484__34_;
      r_484__33_ <= r_n_484__33_;
      r_484__32_ <= r_n_484__32_;
      r_484__31_ <= r_n_484__31_;
      r_484__30_ <= r_n_484__30_;
      r_484__29_ <= r_n_484__29_;
      r_484__28_ <= r_n_484__28_;
      r_484__27_ <= r_n_484__27_;
      r_484__26_ <= r_n_484__26_;
      r_484__25_ <= r_n_484__25_;
      r_484__24_ <= r_n_484__24_;
      r_484__23_ <= r_n_484__23_;
      r_484__22_ <= r_n_484__22_;
      r_484__21_ <= r_n_484__21_;
      r_484__20_ <= r_n_484__20_;
      r_484__19_ <= r_n_484__19_;
      r_484__18_ <= r_n_484__18_;
      r_484__17_ <= r_n_484__17_;
      r_484__16_ <= r_n_484__16_;
      r_484__15_ <= r_n_484__15_;
      r_484__14_ <= r_n_484__14_;
      r_484__13_ <= r_n_484__13_;
      r_484__12_ <= r_n_484__12_;
      r_484__11_ <= r_n_484__11_;
      r_484__10_ <= r_n_484__10_;
      r_484__9_ <= r_n_484__9_;
      r_484__8_ <= r_n_484__8_;
      r_484__7_ <= r_n_484__7_;
      r_484__6_ <= r_n_484__6_;
      r_484__5_ <= r_n_484__5_;
      r_484__4_ <= r_n_484__4_;
      r_484__3_ <= r_n_484__3_;
      r_484__2_ <= r_n_484__2_;
      r_484__1_ <= r_n_484__1_;
      r_484__0_ <= r_n_484__0_;
    end 
    if(N4069) begin
      r_485__63_ <= r_n_485__63_;
      r_485__62_ <= r_n_485__62_;
      r_485__61_ <= r_n_485__61_;
      r_485__60_ <= r_n_485__60_;
      r_485__59_ <= r_n_485__59_;
      r_485__58_ <= r_n_485__58_;
      r_485__57_ <= r_n_485__57_;
      r_485__56_ <= r_n_485__56_;
      r_485__55_ <= r_n_485__55_;
      r_485__54_ <= r_n_485__54_;
      r_485__53_ <= r_n_485__53_;
      r_485__52_ <= r_n_485__52_;
      r_485__51_ <= r_n_485__51_;
      r_485__50_ <= r_n_485__50_;
      r_485__49_ <= r_n_485__49_;
      r_485__48_ <= r_n_485__48_;
      r_485__47_ <= r_n_485__47_;
      r_485__46_ <= r_n_485__46_;
      r_485__45_ <= r_n_485__45_;
      r_485__44_ <= r_n_485__44_;
      r_485__43_ <= r_n_485__43_;
      r_485__42_ <= r_n_485__42_;
      r_485__41_ <= r_n_485__41_;
      r_485__40_ <= r_n_485__40_;
      r_485__39_ <= r_n_485__39_;
      r_485__38_ <= r_n_485__38_;
      r_485__37_ <= r_n_485__37_;
      r_485__36_ <= r_n_485__36_;
      r_485__35_ <= r_n_485__35_;
      r_485__34_ <= r_n_485__34_;
      r_485__33_ <= r_n_485__33_;
      r_485__32_ <= r_n_485__32_;
      r_485__31_ <= r_n_485__31_;
      r_485__30_ <= r_n_485__30_;
      r_485__29_ <= r_n_485__29_;
      r_485__28_ <= r_n_485__28_;
      r_485__27_ <= r_n_485__27_;
      r_485__26_ <= r_n_485__26_;
      r_485__25_ <= r_n_485__25_;
      r_485__24_ <= r_n_485__24_;
      r_485__23_ <= r_n_485__23_;
      r_485__22_ <= r_n_485__22_;
      r_485__21_ <= r_n_485__21_;
      r_485__20_ <= r_n_485__20_;
      r_485__19_ <= r_n_485__19_;
      r_485__18_ <= r_n_485__18_;
      r_485__17_ <= r_n_485__17_;
      r_485__16_ <= r_n_485__16_;
      r_485__15_ <= r_n_485__15_;
      r_485__14_ <= r_n_485__14_;
      r_485__13_ <= r_n_485__13_;
      r_485__12_ <= r_n_485__12_;
      r_485__11_ <= r_n_485__11_;
      r_485__10_ <= r_n_485__10_;
      r_485__9_ <= r_n_485__9_;
      r_485__8_ <= r_n_485__8_;
      r_485__7_ <= r_n_485__7_;
      r_485__6_ <= r_n_485__6_;
      r_485__5_ <= r_n_485__5_;
      r_485__4_ <= r_n_485__4_;
      r_485__3_ <= r_n_485__3_;
      r_485__2_ <= r_n_485__2_;
      r_485__1_ <= r_n_485__1_;
      r_485__0_ <= r_n_485__0_;
    end 
    if(N4070) begin
      r_486__63_ <= r_n_486__63_;
      r_486__62_ <= r_n_486__62_;
      r_486__61_ <= r_n_486__61_;
      r_486__60_ <= r_n_486__60_;
      r_486__59_ <= r_n_486__59_;
      r_486__58_ <= r_n_486__58_;
      r_486__57_ <= r_n_486__57_;
      r_486__56_ <= r_n_486__56_;
      r_486__55_ <= r_n_486__55_;
      r_486__54_ <= r_n_486__54_;
      r_486__53_ <= r_n_486__53_;
      r_486__52_ <= r_n_486__52_;
      r_486__51_ <= r_n_486__51_;
      r_486__50_ <= r_n_486__50_;
      r_486__49_ <= r_n_486__49_;
      r_486__48_ <= r_n_486__48_;
      r_486__47_ <= r_n_486__47_;
      r_486__46_ <= r_n_486__46_;
      r_486__45_ <= r_n_486__45_;
      r_486__44_ <= r_n_486__44_;
      r_486__43_ <= r_n_486__43_;
      r_486__42_ <= r_n_486__42_;
      r_486__41_ <= r_n_486__41_;
      r_486__40_ <= r_n_486__40_;
      r_486__39_ <= r_n_486__39_;
      r_486__38_ <= r_n_486__38_;
      r_486__37_ <= r_n_486__37_;
      r_486__36_ <= r_n_486__36_;
      r_486__35_ <= r_n_486__35_;
      r_486__34_ <= r_n_486__34_;
      r_486__33_ <= r_n_486__33_;
      r_486__32_ <= r_n_486__32_;
      r_486__31_ <= r_n_486__31_;
      r_486__30_ <= r_n_486__30_;
      r_486__29_ <= r_n_486__29_;
      r_486__28_ <= r_n_486__28_;
      r_486__27_ <= r_n_486__27_;
      r_486__26_ <= r_n_486__26_;
      r_486__25_ <= r_n_486__25_;
      r_486__24_ <= r_n_486__24_;
      r_486__23_ <= r_n_486__23_;
      r_486__22_ <= r_n_486__22_;
      r_486__21_ <= r_n_486__21_;
      r_486__20_ <= r_n_486__20_;
      r_486__19_ <= r_n_486__19_;
      r_486__18_ <= r_n_486__18_;
      r_486__17_ <= r_n_486__17_;
      r_486__16_ <= r_n_486__16_;
      r_486__15_ <= r_n_486__15_;
      r_486__14_ <= r_n_486__14_;
      r_486__13_ <= r_n_486__13_;
      r_486__12_ <= r_n_486__12_;
      r_486__11_ <= r_n_486__11_;
      r_486__10_ <= r_n_486__10_;
      r_486__9_ <= r_n_486__9_;
      r_486__8_ <= r_n_486__8_;
      r_486__7_ <= r_n_486__7_;
      r_486__6_ <= r_n_486__6_;
      r_486__5_ <= r_n_486__5_;
      r_486__4_ <= r_n_486__4_;
      r_486__3_ <= r_n_486__3_;
      r_486__2_ <= r_n_486__2_;
      r_486__1_ <= r_n_486__1_;
      r_486__0_ <= r_n_486__0_;
    end 
    if(N4071) begin
      r_487__63_ <= r_n_487__63_;
      r_487__62_ <= r_n_487__62_;
      r_487__61_ <= r_n_487__61_;
      r_487__60_ <= r_n_487__60_;
      r_487__59_ <= r_n_487__59_;
      r_487__58_ <= r_n_487__58_;
      r_487__57_ <= r_n_487__57_;
      r_487__56_ <= r_n_487__56_;
      r_487__55_ <= r_n_487__55_;
      r_487__54_ <= r_n_487__54_;
      r_487__53_ <= r_n_487__53_;
      r_487__52_ <= r_n_487__52_;
      r_487__51_ <= r_n_487__51_;
      r_487__50_ <= r_n_487__50_;
      r_487__49_ <= r_n_487__49_;
      r_487__48_ <= r_n_487__48_;
      r_487__47_ <= r_n_487__47_;
      r_487__46_ <= r_n_487__46_;
      r_487__45_ <= r_n_487__45_;
      r_487__44_ <= r_n_487__44_;
      r_487__43_ <= r_n_487__43_;
      r_487__42_ <= r_n_487__42_;
      r_487__41_ <= r_n_487__41_;
      r_487__40_ <= r_n_487__40_;
      r_487__39_ <= r_n_487__39_;
      r_487__38_ <= r_n_487__38_;
      r_487__37_ <= r_n_487__37_;
      r_487__36_ <= r_n_487__36_;
      r_487__35_ <= r_n_487__35_;
      r_487__34_ <= r_n_487__34_;
      r_487__33_ <= r_n_487__33_;
      r_487__32_ <= r_n_487__32_;
      r_487__31_ <= r_n_487__31_;
      r_487__30_ <= r_n_487__30_;
      r_487__29_ <= r_n_487__29_;
      r_487__28_ <= r_n_487__28_;
      r_487__27_ <= r_n_487__27_;
      r_487__26_ <= r_n_487__26_;
      r_487__25_ <= r_n_487__25_;
      r_487__24_ <= r_n_487__24_;
      r_487__23_ <= r_n_487__23_;
      r_487__22_ <= r_n_487__22_;
      r_487__21_ <= r_n_487__21_;
      r_487__20_ <= r_n_487__20_;
      r_487__19_ <= r_n_487__19_;
      r_487__18_ <= r_n_487__18_;
      r_487__17_ <= r_n_487__17_;
      r_487__16_ <= r_n_487__16_;
      r_487__15_ <= r_n_487__15_;
      r_487__14_ <= r_n_487__14_;
      r_487__13_ <= r_n_487__13_;
      r_487__12_ <= r_n_487__12_;
      r_487__11_ <= r_n_487__11_;
      r_487__10_ <= r_n_487__10_;
      r_487__9_ <= r_n_487__9_;
      r_487__8_ <= r_n_487__8_;
      r_487__7_ <= r_n_487__7_;
      r_487__6_ <= r_n_487__6_;
      r_487__5_ <= r_n_487__5_;
      r_487__4_ <= r_n_487__4_;
      r_487__3_ <= r_n_487__3_;
      r_487__2_ <= r_n_487__2_;
      r_487__1_ <= r_n_487__1_;
      r_487__0_ <= r_n_487__0_;
    end 
    if(N4072) begin
      r_488__63_ <= r_n_488__63_;
      r_488__62_ <= r_n_488__62_;
      r_488__61_ <= r_n_488__61_;
      r_488__60_ <= r_n_488__60_;
      r_488__59_ <= r_n_488__59_;
      r_488__58_ <= r_n_488__58_;
      r_488__57_ <= r_n_488__57_;
      r_488__56_ <= r_n_488__56_;
      r_488__55_ <= r_n_488__55_;
      r_488__54_ <= r_n_488__54_;
      r_488__53_ <= r_n_488__53_;
      r_488__52_ <= r_n_488__52_;
      r_488__51_ <= r_n_488__51_;
      r_488__50_ <= r_n_488__50_;
      r_488__49_ <= r_n_488__49_;
      r_488__48_ <= r_n_488__48_;
      r_488__47_ <= r_n_488__47_;
      r_488__46_ <= r_n_488__46_;
      r_488__45_ <= r_n_488__45_;
      r_488__44_ <= r_n_488__44_;
      r_488__43_ <= r_n_488__43_;
      r_488__42_ <= r_n_488__42_;
      r_488__41_ <= r_n_488__41_;
      r_488__40_ <= r_n_488__40_;
      r_488__39_ <= r_n_488__39_;
      r_488__38_ <= r_n_488__38_;
      r_488__37_ <= r_n_488__37_;
      r_488__36_ <= r_n_488__36_;
      r_488__35_ <= r_n_488__35_;
      r_488__34_ <= r_n_488__34_;
      r_488__33_ <= r_n_488__33_;
      r_488__32_ <= r_n_488__32_;
      r_488__31_ <= r_n_488__31_;
      r_488__30_ <= r_n_488__30_;
      r_488__29_ <= r_n_488__29_;
      r_488__28_ <= r_n_488__28_;
      r_488__27_ <= r_n_488__27_;
      r_488__26_ <= r_n_488__26_;
      r_488__25_ <= r_n_488__25_;
      r_488__24_ <= r_n_488__24_;
      r_488__23_ <= r_n_488__23_;
      r_488__22_ <= r_n_488__22_;
      r_488__21_ <= r_n_488__21_;
      r_488__20_ <= r_n_488__20_;
      r_488__19_ <= r_n_488__19_;
      r_488__18_ <= r_n_488__18_;
      r_488__17_ <= r_n_488__17_;
      r_488__16_ <= r_n_488__16_;
      r_488__15_ <= r_n_488__15_;
      r_488__14_ <= r_n_488__14_;
      r_488__13_ <= r_n_488__13_;
      r_488__12_ <= r_n_488__12_;
      r_488__11_ <= r_n_488__11_;
      r_488__10_ <= r_n_488__10_;
      r_488__9_ <= r_n_488__9_;
      r_488__8_ <= r_n_488__8_;
      r_488__7_ <= r_n_488__7_;
      r_488__6_ <= r_n_488__6_;
      r_488__5_ <= r_n_488__5_;
      r_488__4_ <= r_n_488__4_;
      r_488__3_ <= r_n_488__3_;
      r_488__2_ <= r_n_488__2_;
      r_488__1_ <= r_n_488__1_;
      r_488__0_ <= r_n_488__0_;
    end 
    if(N4073) begin
      r_489__63_ <= r_n_489__63_;
      r_489__62_ <= r_n_489__62_;
      r_489__61_ <= r_n_489__61_;
      r_489__60_ <= r_n_489__60_;
      r_489__59_ <= r_n_489__59_;
      r_489__58_ <= r_n_489__58_;
      r_489__57_ <= r_n_489__57_;
      r_489__56_ <= r_n_489__56_;
      r_489__55_ <= r_n_489__55_;
      r_489__54_ <= r_n_489__54_;
      r_489__53_ <= r_n_489__53_;
      r_489__52_ <= r_n_489__52_;
      r_489__51_ <= r_n_489__51_;
      r_489__50_ <= r_n_489__50_;
      r_489__49_ <= r_n_489__49_;
      r_489__48_ <= r_n_489__48_;
      r_489__47_ <= r_n_489__47_;
      r_489__46_ <= r_n_489__46_;
      r_489__45_ <= r_n_489__45_;
      r_489__44_ <= r_n_489__44_;
      r_489__43_ <= r_n_489__43_;
      r_489__42_ <= r_n_489__42_;
      r_489__41_ <= r_n_489__41_;
      r_489__40_ <= r_n_489__40_;
      r_489__39_ <= r_n_489__39_;
      r_489__38_ <= r_n_489__38_;
      r_489__37_ <= r_n_489__37_;
      r_489__36_ <= r_n_489__36_;
      r_489__35_ <= r_n_489__35_;
      r_489__34_ <= r_n_489__34_;
      r_489__33_ <= r_n_489__33_;
      r_489__32_ <= r_n_489__32_;
      r_489__31_ <= r_n_489__31_;
      r_489__30_ <= r_n_489__30_;
      r_489__29_ <= r_n_489__29_;
      r_489__28_ <= r_n_489__28_;
      r_489__27_ <= r_n_489__27_;
      r_489__26_ <= r_n_489__26_;
      r_489__25_ <= r_n_489__25_;
      r_489__24_ <= r_n_489__24_;
      r_489__23_ <= r_n_489__23_;
      r_489__22_ <= r_n_489__22_;
      r_489__21_ <= r_n_489__21_;
      r_489__20_ <= r_n_489__20_;
      r_489__19_ <= r_n_489__19_;
      r_489__18_ <= r_n_489__18_;
      r_489__17_ <= r_n_489__17_;
      r_489__16_ <= r_n_489__16_;
      r_489__15_ <= r_n_489__15_;
      r_489__14_ <= r_n_489__14_;
      r_489__13_ <= r_n_489__13_;
      r_489__12_ <= r_n_489__12_;
      r_489__11_ <= r_n_489__11_;
      r_489__10_ <= r_n_489__10_;
      r_489__9_ <= r_n_489__9_;
      r_489__8_ <= r_n_489__8_;
      r_489__7_ <= r_n_489__7_;
      r_489__6_ <= r_n_489__6_;
      r_489__5_ <= r_n_489__5_;
      r_489__4_ <= r_n_489__4_;
      r_489__3_ <= r_n_489__3_;
      r_489__2_ <= r_n_489__2_;
      r_489__1_ <= r_n_489__1_;
      r_489__0_ <= r_n_489__0_;
    end 
    if(N4074) begin
      r_490__63_ <= r_n_490__63_;
      r_490__62_ <= r_n_490__62_;
      r_490__61_ <= r_n_490__61_;
      r_490__60_ <= r_n_490__60_;
      r_490__59_ <= r_n_490__59_;
      r_490__58_ <= r_n_490__58_;
      r_490__57_ <= r_n_490__57_;
      r_490__56_ <= r_n_490__56_;
      r_490__55_ <= r_n_490__55_;
      r_490__54_ <= r_n_490__54_;
      r_490__53_ <= r_n_490__53_;
      r_490__52_ <= r_n_490__52_;
      r_490__51_ <= r_n_490__51_;
      r_490__50_ <= r_n_490__50_;
      r_490__49_ <= r_n_490__49_;
      r_490__48_ <= r_n_490__48_;
      r_490__47_ <= r_n_490__47_;
      r_490__46_ <= r_n_490__46_;
      r_490__45_ <= r_n_490__45_;
      r_490__44_ <= r_n_490__44_;
      r_490__43_ <= r_n_490__43_;
      r_490__42_ <= r_n_490__42_;
      r_490__41_ <= r_n_490__41_;
      r_490__40_ <= r_n_490__40_;
      r_490__39_ <= r_n_490__39_;
      r_490__38_ <= r_n_490__38_;
      r_490__37_ <= r_n_490__37_;
      r_490__36_ <= r_n_490__36_;
      r_490__35_ <= r_n_490__35_;
      r_490__34_ <= r_n_490__34_;
      r_490__33_ <= r_n_490__33_;
      r_490__32_ <= r_n_490__32_;
      r_490__31_ <= r_n_490__31_;
      r_490__30_ <= r_n_490__30_;
      r_490__29_ <= r_n_490__29_;
      r_490__28_ <= r_n_490__28_;
      r_490__27_ <= r_n_490__27_;
      r_490__26_ <= r_n_490__26_;
      r_490__25_ <= r_n_490__25_;
      r_490__24_ <= r_n_490__24_;
      r_490__23_ <= r_n_490__23_;
      r_490__22_ <= r_n_490__22_;
      r_490__21_ <= r_n_490__21_;
      r_490__20_ <= r_n_490__20_;
      r_490__19_ <= r_n_490__19_;
      r_490__18_ <= r_n_490__18_;
      r_490__17_ <= r_n_490__17_;
      r_490__16_ <= r_n_490__16_;
      r_490__15_ <= r_n_490__15_;
      r_490__14_ <= r_n_490__14_;
      r_490__13_ <= r_n_490__13_;
      r_490__12_ <= r_n_490__12_;
      r_490__11_ <= r_n_490__11_;
      r_490__10_ <= r_n_490__10_;
      r_490__9_ <= r_n_490__9_;
      r_490__8_ <= r_n_490__8_;
      r_490__7_ <= r_n_490__7_;
      r_490__6_ <= r_n_490__6_;
      r_490__5_ <= r_n_490__5_;
      r_490__4_ <= r_n_490__4_;
      r_490__3_ <= r_n_490__3_;
      r_490__2_ <= r_n_490__2_;
      r_490__1_ <= r_n_490__1_;
      r_490__0_ <= r_n_490__0_;
    end 
    if(N4075) begin
      r_491__63_ <= r_n_491__63_;
      r_491__62_ <= r_n_491__62_;
      r_491__61_ <= r_n_491__61_;
      r_491__60_ <= r_n_491__60_;
      r_491__59_ <= r_n_491__59_;
      r_491__58_ <= r_n_491__58_;
      r_491__57_ <= r_n_491__57_;
      r_491__56_ <= r_n_491__56_;
      r_491__55_ <= r_n_491__55_;
      r_491__54_ <= r_n_491__54_;
      r_491__53_ <= r_n_491__53_;
      r_491__52_ <= r_n_491__52_;
      r_491__51_ <= r_n_491__51_;
      r_491__50_ <= r_n_491__50_;
      r_491__49_ <= r_n_491__49_;
      r_491__48_ <= r_n_491__48_;
      r_491__47_ <= r_n_491__47_;
      r_491__46_ <= r_n_491__46_;
      r_491__45_ <= r_n_491__45_;
      r_491__44_ <= r_n_491__44_;
      r_491__43_ <= r_n_491__43_;
      r_491__42_ <= r_n_491__42_;
      r_491__41_ <= r_n_491__41_;
      r_491__40_ <= r_n_491__40_;
      r_491__39_ <= r_n_491__39_;
      r_491__38_ <= r_n_491__38_;
      r_491__37_ <= r_n_491__37_;
      r_491__36_ <= r_n_491__36_;
      r_491__35_ <= r_n_491__35_;
      r_491__34_ <= r_n_491__34_;
      r_491__33_ <= r_n_491__33_;
      r_491__32_ <= r_n_491__32_;
      r_491__31_ <= r_n_491__31_;
      r_491__30_ <= r_n_491__30_;
      r_491__29_ <= r_n_491__29_;
      r_491__28_ <= r_n_491__28_;
      r_491__27_ <= r_n_491__27_;
      r_491__26_ <= r_n_491__26_;
      r_491__25_ <= r_n_491__25_;
      r_491__24_ <= r_n_491__24_;
      r_491__23_ <= r_n_491__23_;
      r_491__22_ <= r_n_491__22_;
      r_491__21_ <= r_n_491__21_;
      r_491__20_ <= r_n_491__20_;
      r_491__19_ <= r_n_491__19_;
      r_491__18_ <= r_n_491__18_;
      r_491__17_ <= r_n_491__17_;
      r_491__16_ <= r_n_491__16_;
      r_491__15_ <= r_n_491__15_;
      r_491__14_ <= r_n_491__14_;
      r_491__13_ <= r_n_491__13_;
      r_491__12_ <= r_n_491__12_;
      r_491__11_ <= r_n_491__11_;
      r_491__10_ <= r_n_491__10_;
      r_491__9_ <= r_n_491__9_;
      r_491__8_ <= r_n_491__8_;
      r_491__7_ <= r_n_491__7_;
      r_491__6_ <= r_n_491__6_;
      r_491__5_ <= r_n_491__5_;
      r_491__4_ <= r_n_491__4_;
      r_491__3_ <= r_n_491__3_;
      r_491__2_ <= r_n_491__2_;
      r_491__1_ <= r_n_491__1_;
      r_491__0_ <= r_n_491__0_;
    end 
    if(N4076) begin
      r_492__63_ <= r_n_492__63_;
      r_492__62_ <= r_n_492__62_;
      r_492__61_ <= r_n_492__61_;
      r_492__60_ <= r_n_492__60_;
      r_492__59_ <= r_n_492__59_;
      r_492__58_ <= r_n_492__58_;
      r_492__57_ <= r_n_492__57_;
      r_492__56_ <= r_n_492__56_;
      r_492__55_ <= r_n_492__55_;
      r_492__54_ <= r_n_492__54_;
      r_492__53_ <= r_n_492__53_;
      r_492__52_ <= r_n_492__52_;
      r_492__51_ <= r_n_492__51_;
      r_492__50_ <= r_n_492__50_;
      r_492__49_ <= r_n_492__49_;
      r_492__48_ <= r_n_492__48_;
      r_492__47_ <= r_n_492__47_;
      r_492__46_ <= r_n_492__46_;
      r_492__45_ <= r_n_492__45_;
      r_492__44_ <= r_n_492__44_;
      r_492__43_ <= r_n_492__43_;
      r_492__42_ <= r_n_492__42_;
      r_492__41_ <= r_n_492__41_;
      r_492__40_ <= r_n_492__40_;
      r_492__39_ <= r_n_492__39_;
      r_492__38_ <= r_n_492__38_;
      r_492__37_ <= r_n_492__37_;
      r_492__36_ <= r_n_492__36_;
      r_492__35_ <= r_n_492__35_;
      r_492__34_ <= r_n_492__34_;
      r_492__33_ <= r_n_492__33_;
      r_492__32_ <= r_n_492__32_;
      r_492__31_ <= r_n_492__31_;
      r_492__30_ <= r_n_492__30_;
      r_492__29_ <= r_n_492__29_;
      r_492__28_ <= r_n_492__28_;
      r_492__27_ <= r_n_492__27_;
      r_492__26_ <= r_n_492__26_;
      r_492__25_ <= r_n_492__25_;
      r_492__24_ <= r_n_492__24_;
      r_492__23_ <= r_n_492__23_;
      r_492__22_ <= r_n_492__22_;
      r_492__21_ <= r_n_492__21_;
      r_492__20_ <= r_n_492__20_;
      r_492__19_ <= r_n_492__19_;
      r_492__18_ <= r_n_492__18_;
      r_492__17_ <= r_n_492__17_;
      r_492__16_ <= r_n_492__16_;
      r_492__15_ <= r_n_492__15_;
      r_492__14_ <= r_n_492__14_;
      r_492__13_ <= r_n_492__13_;
      r_492__12_ <= r_n_492__12_;
      r_492__11_ <= r_n_492__11_;
      r_492__10_ <= r_n_492__10_;
      r_492__9_ <= r_n_492__9_;
      r_492__8_ <= r_n_492__8_;
      r_492__7_ <= r_n_492__7_;
      r_492__6_ <= r_n_492__6_;
      r_492__5_ <= r_n_492__5_;
      r_492__4_ <= r_n_492__4_;
      r_492__3_ <= r_n_492__3_;
      r_492__2_ <= r_n_492__2_;
      r_492__1_ <= r_n_492__1_;
      r_492__0_ <= r_n_492__0_;
    end 
    if(N4077) begin
      r_493__63_ <= r_n_493__63_;
      r_493__62_ <= r_n_493__62_;
      r_493__61_ <= r_n_493__61_;
      r_493__60_ <= r_n_493__60_;
      r_493__59_ <= r_n_493__59_;
      r_493__58_ <= r_n_493__58_;
      r_493__57_ <= r_n_493__57_;
      r_493__56_ <= r_n_493__56_;
      r_493__55_ <= r_n_493__55_;
      r_493__54_ <= r_n_493__54_;
      r_493__53_ <= r_n_493__53_;
      r_493__52_ <= r_n_493__52_;
      r_493__51_ <= r_n_493__51_;
      r_493__50_ <= r_n_493__50_;
      r_493__49_ <= r_n_493__49_;
      r_493__48_ <= r_n_493__48_;
      r_493__47_ <= r_n_493__47_;
      r_493__46_ <= r_n_493__46_;
      r_493__45_ <= r_n_493__45_;
      r_493__44_ <= r_n_493__44_;
      r_493__43_ <= r_n_493__43_;
      r_493__42_ <= r_n_493__42_;
      r_493__41_ <= r_n_493__41_;
      r_493__40_ <= r_n_493__40_;
      r_493__39_ <= r_n_493__39_;
      r_493__38_ <= r_n_493__38_;
      r_493__37_ <= r_n_493__37_;
      r_493__36_ <= r_n_493__36_;
      r_493__35_ <= r_n_493__35_;
      r_493__34_ <= r_n_493__34_;
      r_493__33_ <= r_n_493__33_;
      r_493__32_ <= r_n_493__32_;
      r_493__31_ <= r_n_493__31_;
      r_493__30_ <= r_n_493__30_;
      r_493__29_ <= r_n_493__29_;
      r_493__28_ <= r_n_493__28_;
      r_493__27_ <= r_n_493__27_;
      r_493__26_ <= r_n_493__26_;
      r_493__25_ <= r_n_493__25_;
      r_493__24_ <= r_n_493__24_;
      r_493__23_ <= r_n_493__23_;
      r_493__22_ <= r_n_493__22_;
      r_493__21_ <= r_n_493__21_;
      r_493__20_ <= r_n_493__20_;
      r_493__19_ <= r_n_493__19_;
      r_493__18_ <= r_n_493__18_;
      r_493__17_ <= r_n_493__17_;
      r_493__16_ <= r_n_493__16_;
      r_493__15_ <= r_n_493__15_;
      r_493__14_ <= r_n_493__14_;
      r_493__13_ <= r_n_493__13_;
      r_493__12_ <= r_n_493__12_;
      r_493__11_ <= r_n_493__11_;
      r_493__10_ <= r_n_493__10_;
      r_493__9_ <= r_n_493__9_;
      r_493__8_ <= r_n_493__8_;
      r_493__7_ <= r_n_493__7_;
      r_493__6_ <= r_n_493__6_;
      r_493__5_ <= r_n_493__5_;
      r_493__4_ <= r_n_493__4_;
      r_493__3_ <= r_n_493__3_;
      r_493__2_ <= r_n_493__2_;
      r_493__1_ <= r_n_493__1_;
      r_493__0_ <= r_n_493__0_;
    end 
    if(N4078) begin
      r_494__63_ <= r_n_494__63_;
      r_494__62_ <= r_n_494__62_;
      r_494__61_ <= r_n_494__61_;
      r_494__60_ <= r_n_494__60_;
      r_494__59_ <= r_n_494__59_;
      r_494__58_ <= r_n_494__58_;
      r_494__57_ <= r_n_494__57_;
      r_494__56_ <= r_n_494__56_;
      r_494__55_ <= r_n_494__55_;
      r_494__54_ <= r_n_494__54_;
      r_494__53_ <= r_n_494__53_;
      r_494__52_ <= r_n_494__52_;
      r_494__51_ <= r_n_494__51_;
      r_494__50_ <= r_n_494__50_;
      r_494__49_ <= r_n_494__49_;
      r_494__48_ <= r_n_494__48_;
      r_494__47_ <= r_n_494__47_;
      r_494__46_ <= r_n_494__46_;
      r_494__45_ <= r_n_494__45_;
      r_494__44_ <= r_n_494__44_;
      r_494__43_ <= r_n_494__43_;
      r_494__42_ <= r_n_494__42_;
      r_494__41_ <= r_n_494__41_;
      r_494__40_ <= r_n_494__40_;
      r_494__39_ <= r_n_494__39_;
      r_494__38_ <= r_n_494__38_;
      r_494__37_ <= r_n_494__37_;
      r_494__36_ <= r_n_494__36_;
      r_494__35_ <= r_n_494__35_;
      r_494__34_ <= r_n_494__34_;
      r_494__33_ <= r_n_494__33_;
      r_494__32_ <= r_n_494__32_;
      r_494__31_ <= r_n_494__31_;
      r_494__30_ <= r_n_494__30_;
      r_494__29_ <= r_n_494__29_;
      r_494__28_ <= r_n_494__28_;
      r_494__27_ <= r_n_494__27_;
      r_494__26_ <= r_n_494__26_;
      r_494__25_ <= r_n_494__25_;
      r_494__24_ <= r_n_494__24_;
      r_494__23_ <= r_n_494__23_;
      r_494__22_ <= r_n_494__22_;
      r_494__21_ <= r_n_494__21_;
      r_494__20_ <= r_n_494__20_;
      r_494__19_ <= r_n_494__19_;
      r_494__18_ <= r_n_494__18_;
      r_494__17_ <= r_n_494__17_;
      r_494__16_ <= r_n_494__16_;
      r_494__15_ <= r_n_494__15_;
      r_494__14_ <= r_n_494__14_;
      r_494__13_ <= r_n_494__13_;
      r_494__12_ <= r_n_494__12_;
      r_494__11_ <= r_n_494__11_;
      r_494__10_ <= r_n_494__10_;
      r_494__9_ <= r_n_494__9_;
      r_494__8_ <= r_n_494__8_;
      r_494__7_ <= r_n_494__7_;
      r_494__6_ <= r_n_494__6_;
      r_494__5_ <= r_n_494__5_;
      r_494__4_ <= r_n_494__4_;
      r_494__3_ <= r_n_494__3_;
      r_494__2_ <= r_n_494__2_;
      r_494__1_ <= r_n_494__1_;
      r_494__0_ <= r_n_494__0_;
    end 
    if(N4079) begin
      r_495__63_ <= r_n_495__63_;
      r_495__62_ <= r_n_495__62_;
      r_495__61_ <= r_n_495__61_;
      r_495__60_ <= r_n_495__60_;
      r_495__59_ <= r_n_495__59_;
      r_495__58_ <= r_n_495__58_;
      r_495__57_ <= r_n_495__57_;
      r_495__56_ <= r_n_495__56_;
      r_495__55_ <= r_n_495__55_;
      r_495__54_ <= r_n_495__54_;
      r_495__53_ <= r_n_495__53_;
      r_495__52_ <= r_n_495__52_;
      r_495__51_ <= r_n_495__51_;
      r_495__50_ <= r_n_495__50_;
      r_495__49_ <= r_n_495__49_;
      r_495__48_ <= r_n_495__48_;
      r_495__47_ <= r_n_495__47_;
      r_495__46_ <= r_n_495__46_;
      r_495__45_ <= r_n_495__45_;
      r_495__44_ <= r_n_495__44_;
      r_495__43_ <= r_n_495__43_;
      r_495__42_ <= r_n_495__42_;
      r_495__41_ <= r_n_495__41_;
      r_495__40_ <= r_n_495__40_;
      r_495__39_ <= r_n_495__39_;
      r_495__38_ <= r_n_495__38_;
      r_495__37_ <= r_n_495__37_;
      r_495__36_ <= r_n_495__36_;
      r_495__35_ <= r_n_495__35_;
      r_495__34_ <= r_n_495__34_;
      r_495__33_ <= r_n_495__33_;
      r_495__32_ <= r_n_495__32_;
      r_495__31_ <= r_n_495__31_;
      r_495__30_ <= r_n_495__30_;
      r_495__29_ <= r_n_495__29_;
      r_495__28_ <= r_n_495__28_;
      r_495__27_ <= r_n_495__27_;
      r_495__26_ <= r_n_495__26_;
      r_495__25_ <= r_n_495__25_;
      r_495__24_ <= r_n_495__24_;
      r_495__23_ <= r_n_495__23_;
      r_495__22_ <= r_n_495__22_;
      r_495__21_ <= r_n_495__21_;
      r_495__20_ <= r_n_495__20_;
      r_495__19_ <= r_n_495__19_;
      r_495__18_ <= r_n_495__18_;
      r_495__17_ <= r_n_495__17_;
      r_495__16_ <= r_n_495__16_;
      r_495__15_ <= r_n_495__15_;
      r_495__14_ <= r_n_495__14_;
      r_495__13_ <= r_n_495__13_;
      r_495__12_ <= r_n_495__12_;
      r_495__11_ <= r_n_495__11_;
      r_495__10_ <= r_n_495__10_;
      r_495__9_ <= r_n_495__9_;
      r_495__8_ <= r_n_495__8_;
      r_495__7_ <= r_n_495__7_;
      r_495__6_ <= r_n_495__6_;
      r_495__5_ <= r_n_495__5_;
      r_495__4_ <= r_n_495__4_;
      r_495__3_ <= r_n_495__3_;
      r_495__2_ <= r_n_495__2_;
      r_495__1_ <= r_n_495__1_;
      r_495__0_ <= r_n_495__0_;
    end 
    if(N4080) begin
      r_496__63_ <= r_n_496__63_;
      r_496__62_ <= r_n_496__62_;
      r_496__61_ <= r_n_496__61_;
      r_496__60_ <= r_n_496__60_;
      r_496__59_ <= r_n_496__59_;
      r_496__58_ <= r_n_496__58_;
      r_496__57_ <= r_n_496__57_;
      r_496__56_ <= r_n_496__56_;
      r_496__55_ <= r_n_496__55_;
      r_496__54_ <= r_n_496__54_;
      r_496__53_ <= r_n_496__53_;
      r_496__52_ <= r_n_496__52_;
      r_496__51_ <= r_n_496__51_;
      r_496__50_ <= r_n_496__50_;
      r_496__49_ <= r_n_496__49_;
      r_496__48_ <= r_n_496__48_;
      r_496__47_ <= r_n_496__47_;
      r_496__46_ <= r_n_496__46_;
      r_496__45_ <= r_n_496__45_;
      r_496__44_ <= r_n_496__44_;
      r_496__43_ <= r_n_496__43_;
      r_496__42_ <= r_n_496__42_;
      r_496__41_ <= r_n_496__41_;
      r_496__40_ <= r_n_496__40_;
      r_496__39_ <= r_n_496__39_;
      r_496__38_ <= r_n_496__38_;
      r_496__37_ <= r_n_496__37_;
      r_496__36_ <= r_n_496__36_;
      r_496__35_ <= r_n_496__35_;
      r_496__34_ <= r_n_496__34_;
      r_496__33_ <= r_n_496__33_;
      r_496__32_ <= r_n_496__32_;
      r_496__31_ <= r_n_496__31_;
      r_496__30_ <= r_n_496__30_;
      r_496__29_ <= r_n_496__29_;
      r_496__28_ <= r_n_496__28_;
      r_496__27_ <= r_n_496__27_;
      r_496__26_ <= r_n_496__26_;
      r_496__25_ <= r_n_496__25_;
      r_496__24_ <= r_n_496__24_;
      r_496__23_ <= r_n_496__23_;
      r_496__22_ <= r_n_496__22_;
      r_496__21_ <= r_n_496__21_;
      r_496__20_ <= r_n_496__20_;
      r_496__19_ <= r_n_496__19_;
      r_496__18_ <= r_n_496__18_;
      r_496__17_ <= r_n_496__17_;
      r_496__16_ <= r_n_496__16_;
      r_496__15_ <= r_n_496__15_;
      r_496__14_ <= r_n_496__14_;
      r_496__13_ <= r_n_496__13_;
      r_496__12_ <= r_n_496__12_;
      r_496__11_ <= r_n_496__11_;
      r_496__10_ <= r_n_496__10_;
      r_496__9_ <= r_n_496__9_;
      r_496__8_ <= r_n_496__8_;
      r_496__7_ <= r_n_496__7_;
      r_496__6_ <= r_n_496__6_;
      r_496__5_ <= r_n_496__5_;
      r_496__4_ <= r_n_496__4_;
      r_496__3_ <= r_n_496__3_;
      r_496__2_ <= r_n_496__2_;
      r_496__1_ <= r_n_496__1_;
      r_496__0_ <= r_n_496__0_;
    end 
    if(N4081) begin
      r_497__63_ <= r_n_497__63_;
      r_497__62_ <= r_n_497__62_;
      r_497__61_ <= r_n_497__61_;
      r_497__60_ <= r_n_497__60_;
      r_497__59_ <= r_n_497__59_;
      r_497__58_ <= r_n_497__58_;
      r_497__57_ <= r_n_497__57_;
      r_497__56_ <= r_n_497__56_;
      r_497__55_ <= r_n_497__55_;
      r_497__54_ <= r_n_497__54_;
      r_497__53_ <= r_n_497__53_;
      r_497__52_ <= r_n_497__52_;
      r_497__51_ <= r_n_497__51_;
      r_497__50_ <= r_n_497__50_;
      r_497__49_ <= r_n_497__49_;
      r_497__48_ <= r_n_497__48_;
      r_497__47_ <= r_n_497__47_;
      r_497__46_ <= r_n_497__46_;
      r_497__45_ <= r_n_497__45_;
      r_497__44_ <= r_n_497__44_;
      r_497__43_ <= r_n_497__43_;
      r_497__42_ <= r_n_497__42_;
      r_497__41_ <= r_n_497__41_;
      r_497__40_ <= r_n_497__40_;
      r_497__39_ <= r_n_497__39_;
      r_497__38_ <= r_n_497__38_;
      r_497__37_ <= r_n_497__37_;
      r_497__36_ <= r_n_497__36_;
      r_497__35_ <= r_n_497__35_;
      r_497__34_ <= r_n_497__34_;
      r_497__33_ <= r_n_497__33_;
      r_497__32_ <= r_n_497__32_;
      r_497__31_ <= r_n_497__31_;
      r_497__30_ <= r_n_497__30_;
      r_497__29_ <= r_n_497__29_;
      r_497__28_ <= r_n_497__28_;
      r_497__27_ <= r_n_497__27_;
      r_497__26_ <= r_n_497__26_;
      r_497__25_ <= r_n_497__25_;
      r_497__24_ <= r_n_497__24_;
      r_497__23_ <= r_n_497__23_;
      r_497__22_ <= r_n_497__22_;
      r_497__21_ <= r_n_497__21_;
      r_497__20_ <= r_n_497__20_;
      r_497__19_ <= r_n_497__19_;
      r_497__18_ <= r_n_497__18_;
      r_497__17_ <= r_n_497__17_;
      r_497__16_ <= r_n_497__16_;
      r_497__15_ <= r_n_497__15_;
      r_497__14_ <= r_n_497__14_;
      r_497__13_ <= r_n_497__13_;
      r_497__12_ <= r_n_497__12_;
      r_497__11_ <= r_n_497__11_;
      r_497__10_ <= r_n_497__10_;
      r_497__9_ <= r_n_497__9_;
      r_497__8_ <= r_n_497__8_;
      r_497__7_ <= r_n_497__7_;
      r_497__6_ <= r_n_497__6_;
      r_497__5_ <= r_n_497__5_;
      r_497__4_ <= r_n_497__4_;
      r_497__3_ <= r_n_497__3_;
      r_497__2_ <= r_n_497__2_;
      r_497__1_ <= r_n_497__1_;
      r_497__0_ <= r_n_497__0_;
    end 
    if(N4082) begin
      r_498__63_ <= r_n_498__63_;
      r_498__62_ <= r_n_498__62_;
      r_498__61_ <= r_n_498__61_;
      r_498__60_ <= r_n_498__60_;
      r_498__59_ <= r_n_498__59_;
      r_498__58_ <= r_n_498__58_;
      r_498__57_ <= r_n_498__57_;
      r_498__56_ <= r_n_498__56_;
      r_498__55_ <= r_n_498__55_;
      r_498__54_ <= r_n_498__54_;
      r_498__53_ <= r_n_498__53_;
      r_498__52_ <= r_n_498__52_;
      r_498__51_ <= r_n_498__51_;
      r_498__50_ <= r_n_498__50_;
      r_498__49_ <= r_n_498__49_;
      r_498__48_ <= r_n_498__48_;
      r_498__47_ <= r_n_498__47_;
      r_498__46_ <= r_n_498__46_;
      r_498__45_ <= r_n_498__45_;
      r_498__44_ <= r_n_498__44_;
      r_498__43_ <= r_n_498__43_;
      r_498__42_ <= r_n_498__42_;
      r_498__41_ <= r_n_498__41_;
      r_498__40_ <= r_n_498__40_;
      r_498__39_ <= r_n_498__39_;
      r_498__38_ <= r_n_498__38_;
      r_498__37_ <= r_n_498__37_;
      r_498__36_ <= r_n_498__36_;
      r_498__35_ <= r_n_498__35_;
      r_498__34_ <= r_n_498__34_;
      r_498__33_ <= r_n_498__33_;
      r_498__32_ <= r_n_498__32_;
      r_498__31_ <= r_n_498__31_;
      r_498__30_ <= r_n_498__30_;
      r_498__29_ <= r_n_498__29_;
      r_498__28_ <= r_n_498__28_;
      r_498__27_ <= r_n_498__27_;
      r_498__26_ <= r_n_498__26_;
      r_498__25_ <= r_n_498__25_;
      r_498__24_ <= r_n_498__24_;
      r_498__23_ <= r_n_498__23_;
      r_498__22_ <= r_n_498__22_;
      r_498__21_ <= r_n_498__21_;
      r_498__20_ <= r_n_498__20_;
      r_498__19_ <= r_n_498__19_;
      r_498__18_ <= r_n_498__18_;
      r_498__17_ <= r_n_498__17_;
      r_498__16_ <= r_n_498__16_;
      r_498__15_ <= r_n_498__15_;
      r_498__14_ <= r_n_498__14_;
      r_498__13_ <= r_n_498__13_;
      r_498__12_ <= r_n_498__12_;
      r_498__11_ <= r_n_498__11_;
      r_498__10_ <= r_n_498__10_;
      r_498__9_ <= r_n_498__9_;
      r_498__8_ <= r_n_498__8_;
      r_498__7_ <= r_n_498__7_;
      r_498__6_ <= r_n_498__6_;
      r_498__5_ <= r_n_498__5_;
      r_498__4_ <= r_n_498__4_;
      r_498__3_ <= r_n_498__3_;
      r_498__2_ <= r_n_498__2_;
      r_498__1_ <= r_n_498__1_;
      r_498__0_ <= r_n_498__0_;
    end 
    if(N4083) begin
      r_499__63_ <= r_n_499__63_;
      r_499__62_ <= r_n_499__62_;
      r_499__61_ <= r_n_499__61_;
      r_499__60_ <= r_n_499__60_;
      r_499__59_ <= r_n_499__59_;
      r_499__58_ <= r_n_499__58_;
      r_499__57_ <= r_n_499__57_;
      r_499__56_ <= r_n_499__56_;
      r_499__55_ <= r_n_499__55_;
      r_499__54_ <= r_n_499__54_;
      r_499__53_ <= r_n_499__53_;
      r_499__52_ <= r_n_499__52_;
      r_499__51_ <= r_n_499__51_;
      r_499__50_ <= r_n_499__50_;
      r_499__49_ <= r_n_499__49_;
      r_499__48_ <= r_n_499__48_;
      r_499__47_ <= r_n_499__47_;
      r_499__46_ <= r_n_499__46_;
      r_499__45_ <= r_n_499__45_;
      r_499__44_ <= r_n_499__44_;
      r_499__43_ <= r_n_499__43_;
      r_499__42_ <= r_n_499__42_;
      r_499__41_ <= r_n_499__41_;
      r_499__40_ <= r_n_499__40_;
      r_499__39_ <= r_n_499__39_;
      r_499__38_ <= r_n_499__38_;
      r_499__37_ <= r_n_499__37_;
      r_499__36_ <= r_n_499__36_;
      r_499__35_ <= r_n_499__35_;
      r_499__34_ <= r_n_499__34_;
      r_499__33_ <= r_n_499__33_;
      r_499__32_ <= r_n_499__32_;
      r_499__31_ <= r_n_499__31_;
      r_499__30_ <= r_n_499__30_;
      r_499__29_ <= r_n_499__29_;
      r_499__28_ <= r_n_499__28_;
      r_499__27_ <= r_n_499__27_;
      r_499__26_ <= r_n_499__26_;
      r_499__25_ <= r_n_499__25_;
      r_499__24_ <= r_n_499__24_;
      r_499__23_ <= r_n_499__23_;
      r_499__22_ <= r_n_499__22_;
      r_499__21_ <= r_n_499__21_;
      r_499__20_ <= r_n_499__20_;
      r_499__19_ <= r_n_499__19_;
      r_499__18_ <= r_n_499__18_;
      r_499__17_ <= r_n_499__17_;
      r_499__16_ <= r_n_499__16_;
      r_499__15_ <= r_n_499__15_;
      r_499__14_ <= r_n_499__14_;
      r_499__13_ <= r_n_499__13_;
      r_499__12_ <= r_n_499__12_;
      r_499__11_ <= r_n_499__11_;
      r_499__10_ <= r_n_499__10_;
      r_499__9_ <= r_n_499__9_;
      r_499__8_ <= r_n_499__8_;
      r_499__7_ <= r_n_499__7_;
      r_499__6_ <= r_n_499__6_;
      r_499__5_ <= r_n_499__5_;
      r_499__4_ <= r_n_499__4_;
      r_499__3_ <= r_n_499__3_;
      r_499__2_ <= r_n_499__2_;
      r_499__1_ <= r_n_499__1_;
      r_499__0_ <= r_n_499__0_;
    end 
    if(N4084) begin
      r_500__63_ <= r_n_500__63_;
      r_500__62_ <= r_n_500__62_;
      r_500__61_ <= r_n_500__61_;
      r_500__60_ <= r_n_500__60_;
      r_500__59_ <= r_n_500__59_;
      r_500__58_ <= r_n_500__58_;
      r_500__57_ <= r_n_500__57_;
      r_500__56_ <= r_n_500__56_;
      r_500__55_ <= r_n_500__55_;
      r_500__54_ <= r_n_500__54_;
      r_500__53_ <= r_n_500__53_;
      r_500__52_ <= r_n_500__52_;
      r_500__51_ <= r_n_500__51_;
      r_500__50_ <= r_n_500__50_;
      r_500__49_ <= r_n_500__49_;
      r_500__48_ <= r_n_500__48_;
      r_500__47_ <= r_n_500__47_;
      r_500__46_ <= r_n_500__46_;
      r_500__45_ <= r_n_500__45_;
      r_500__44_ <= r_n_500__44_;
      r_500__43_ <= r_n_500__43_;
      r_500__42_ <= r_n_500__42_;
      r_500__41_ <= r_n_500__41_;
      r_500__40_ <= r_n_500__40_;
      r_500__39_ <= r_n_500__39_;
      r_500__38_ <= r_n_500__38_;
      r_500__37_ <= r_n_500__37_;
      r_500__36_ <= r_n_500__36_;
      r_500__35_ <= r_n_500__35_;
      r_500__34_ <= r_n_500__34_;
      r_500__33_ <= r_n_500__33_;
      r_500__32_ <= r_n_500__32_;
      r_500__31_ <= r_n_500__31_;
      r_500__30_ <= r_n_500__30_;
      r_500__29_ <= r_n_500__29_;
      r_500__28_ <= r_n_500__28_;
      r_500__27_ <= r_n_500__27_;
      r_500__26_ <= r_n_500__26_;
      r_500__25_ <= r_n_500__25_;
      r_500__24_ <= r_n_500__24_;
      r_500__23_ <= r_n_500__23_;
      r_500__22_ <= r_n_500__22_;
      r_500__21_ <= r_n_500__21_;
      r_500__20_ <= r_n_500__20_;
      r_500__19_ <= r_n_500__19_;
      r_500__18_ <= r_n_500__18_;
      r_500__17_ <= r_n_500__17_;
      r_500__16_ <= r_n_500__16_;
      r_500__15_ <= r_n_500__15_;
      r_500__14_ <= r_n_500__14_;
      r_500__13_ <= r_n_500__13_;
      r_500__12_ <= r_n_500__12_;
      r_500__11_ <= r_n_500__11_;
      r_500__10_ <= r_n_500__10_;
      r_500__9_ <= r_n_500__9_;
      r_500__8_ <= r_n_500__8_;
      r_500__7_ <= r_n_500__7_;
      r_500__6_ <= r_n_500__6_;
      r_500__5_ <= r_n_500__5_;
      r_500__4_ <= r_n_500__4_;
      r_500__3_ <= r_n_500__3_;
      r_500__2_ <= r_n_500__2_;
      r_500__1_ <= r_n_500__1_;
      r_500__0_ <= r_n_500__0_;
    end 
    if(N4085) begin
      r_501__63_ <= r_n_501__63_;
      r_501__62_ <= r_n_501__62_;
      r_501__61_ <= r_n_501__61_;
      r_501__60_ <= r_n_501__60_;
      r_501__59_ <= r_n_501__59_;
      r_501__58_ <= r_n_501__58_;
      r_501__57_ <= r_n_501__57_;
      r_501__56_ <= r_n_501__56_;
      r_501__55_ <= r_n_501__55_;
      r_501__54_ <= r_n_501__54_;
      r_501__53_ <= r_n_501__53_;
      r_501__52_ <= r_n_501__52_;
      r_501__51_ <= r_n_501__51_;
      r_501__50_ <= r_n_501__50_;
      r_501__49_ <= r_n_501__49_;
      r_501__48_ <= r_n_501__48_;
      r_501__47_ <= r_n_501__47_;
      r_501__46_ <= r_n_501__46_;
      r_501__45_ <= r_n_501__45_;
      r_501__44_ <= r_n_501__44_;
      r_501__43_ <= r_n_501__43_;
      r_501__42_ <= r_n_501__42_;
      r_501__41_ <= r_n_501__41_;
      r_501__40_ <= r_n_501__40_;
      r_501__39_ <= r_n_501__39_;
      r_501__38_ <= r_n_501__38_;
      r_501__37_ <= r_n_501__37_;
      r_501__36_ <= r_n_501__36_;
      r_501__35_ <= r_n_501__35_;
      r_501__34_ <= r_n_501__34_;
      r_501__33_ <= r_n_501__33_;
      r_501__32_ <= r_n_501__32_;
      r_501__31_ <= r_n_501__31_;
      r_501__30_ <= r_n_501__30_;
      r_501__29_ <= r_n_501__29_;
      r_501__28_ <= r_n_501__28_;
      r_501__27_ <= r_n_501__27_;
      r_501__26_ <= r_n_501__26_;
      r_501__25_ <= r_n_501__25_;
      r_501__24_ <= r_n_501__24_;
      r_501__23_ <= r_n_501__23_;
      r_501__22_ <= r_n_501__22_;
      r_501__21_ <= r_n_501__21_;
      r_501__20_ <= r_n_501__20_;
      r_501__19_ <= r_n_501__19_;
      r_501__18_ <= r_n_501__18_;
      r_501__17_ <= r_n_501__17_;
      r_501__16_ <= r_n_501__16_;
      r_501__15_ <= r_n_501__15_;
      r_501__14_ <= r_n_501__14_;
      r_501__13_ <= r_n_501__13_;
      r_501__12_ <= r_n_501__12_;
      r_501__11_ <= r_n_501__11_;
      r_501__10_ <= r_n_501__10_;
      r_501__9_ <= r_n_501__9_;
      r_501__8_ <= r_n_501__8_;
      r_501__7_ <= r_n_501__7_;
      r_501__6_ <= r_n_501__6_;
      r_501__5_ <= r_n_501__5_;
      r_501__4_ <= r_n_501__4_;
      r_501__3_ <= r_n_501__3_;
      r_501__2_ <= r_n_501__2_;
      r_501__1_ <= r_n_501__1_;
      r_501__0_ <= r_n_501__0_;
    end 
    if(N4086) begin
      r_502__63_ <= r_n_502__63_;
      r_502__62_ <= r_n_502__62_;
      r_502__61_ <= r_n_502__61_;
      r_502__60_ <= r_n_502__60_;
      r_502__59_ <= r_n_502__59_;
      r_502__58_ <= r_n_502__58_;
      r_502__57_ <= r_n_502__57_;
      r_502__56_ <= r_n_502__56_;
      r_502__55_ <= r_n_502__55_;
      r_502__54_ <= r_n_502__54_;
      r_502__53_ <= r_n_502__53_;
      r_502__52_ <= r_n_502__52_;
      r_502__51_ <= r_n_502__51_;
      r_502__50_ <= r_n_502__50_;
      r_502__49_ <= r_n_502__49_;
      r_502__48_ <= r_n_502__48_;
      r_502__47_ <= r_n_502__47_;
      r_502__46_ <= r_n_502__46_;
      r_502__45_ <= r_n_502__45_;
      r_502__44_ <= r_n_502__44_;
      r_502__43_ <= r_n_502__43_;
      r_502__42_ <= r_n_502__42_;
      r_502__41_ <= r_n_502__41_;
      r_502__40_ <= r_n_502__40_;
      r_502__39_ <= r_n_502__39_;
      r_502__38_ <= r_n_502__38_;
      r_502__37_ <= r_n_502__37_;
      r_502__36_ <= r_n_502__36_;
      r_502__35_ <= r_n_502__35_;
      r_502__34_ <= r_n_502__34_;
      r_502__33_ <= r_n_502__33_;
      r_502__32_ <= r_n_502__32_;
      r_502__31_ <= r_n_502__31_;
      r_502__30_ <= r_n_502__30_;
      r_502__29_ <= r_n_502__29_;
      r_502__28_ <= r_n_502__28_;
      r_502__27_ <= r_n_502__27_;
      r_502__26_ <= r_n_502__26_;
      r_502__25_ <= r_n_502__25_;
      r_502__24_ <= r_n_502__24_;
      r_502__23_ <= r_n_502__23_;
      r_502__22_ <= r_n_502__22_;
      r_502__21_ <= r_n_502__21_;
      r_502__20_ <= r_n_502__20_;
      r_502__19_ <= r_n_502__19_;
      r_502__18_ <= r_n_502__18_;
      r_502__17_ <= r_n_502__17_;
      r_502__16_ <= r_n_502__16_;
      r_502__15_ <= r_n_502__15_;
      r_502__14_ <= r_n_502__14_;
      r_502__13_ <= r_n_502__13_;
      r_502__12_ <= r_n_502__12_;
      r_502__11_ <= r_n_502__11_;
      r_502__10_ <= r_n_502__10_;
      r_502__9_ <= r_n_502__9_;
      r_502__8_ <= r_n_502__8_;
      r_502__7_ <= r_n_502__7_;
      r_502__6_ <= r_n_502__6_;
      r_502__5_ <= r_n_502__5_;
      r_502__4_ <= r_n_502__4_;
      r_502__3_ <= r_n_502__3_;
      r_502__2_ <= r_n_502__2_;
      r_502__1_ <= r_n_502__1_;
      r_502__0_ <= r_n_502__0_;
    end 
    if(N4087) begin
      r_503__63_ <= r_n_503__63_;
      r_503__62_ <= r_n_503__62_;
      r_503__61_ <= r_n_503__61_;
      r_503__60_ <= r_n_503__60_;
      r_503__59_ <= r_n_503__59_;
      r_503__58_ <= r_n_503__58_;
      r_503__57_ <= r_n_503__57_;
      r_503__56_ <= r_n_503__56_;
      r_503__55_ <= r_n_503__55_;
      r_503__54_ <= r_n_503__54_;
      r_503__53_ <= r_n_503__53_;
      r_503__52_ <= r_n_503__52_;
      r_503__51_ <= r_n_503__51_;
      r_503__50_ <= r_n_503__50_;
      r_503__49_ <= r_n_503__49_;
      r_503__48_ <= r_n_503__48_;
      r_503__47_ <= r_n_503__47_;
      r_503__46_ <= r_n_503__46_;
      r_503__45_ <= r_n_503__45_;
      r_503__44_ <= r_n_503__44_;
      r_503__43_ <= r_n_503__43_;
      r_503__42_ <= r_n_503__42_;
      r_503__41_ <= r_n_503__41_;
      r_503__40_ <= r_n_503__40_;
      r_503__39_ <= r_n_503__39_;
      r_503__38_ <= r_n_503__38_;
      r_503__37_ <= r_n_503__37_;
      r_503__36_ <= r_n_503__36_;
      r_503__35_ <= r_n_503__35_;
      r_503__34_ <= r_n_503__34_;
      r_503__33_ <= r_n_503__33_;
      r_503__32_ <= r_n_503__32_;
      r_503__31_ <= r_n_503__31_;
      r_503__30_ <= r_n_503__30_;
      r_503__29_ <= r_n_503__29_;
      r_503__28_ <= r_n_503__28_;
      r_503__27_ <= r_n_503__27_;
      r_503__26_ <= r_n_503__26_;
      r_503__25_ <= r_n_503__25_;
      r_503__24_ <= r_n_503__24_;
      r_503__23_ <= r_n_503__23_;
      r_503__22_ <= r_n_503__22_;
      r_503__21_ <= r_n_503__21_;
      r_503__20_ <= r_n_503__20_;
      r_503__19_ <= r_n_503__19_;
      r_503__18_ <= r_n_503__18_;
      r_503__17_ <= r_n_503__17_;
      r_503__16_ <= r_n_503__16_;
      r_503__15_ <= r_n_503__15_;
      r_503__14_ <= r_n_503__14_;
      r_503__13_ <= r_n_503__13_;
      r_503__12_ <= r_n_503__12_;
      r_503__11_ <= r_n_503__11_;
      r_503__10_ <= r_n_503__10_;
      r_503__9_ <= r_n_503__9_;
      r_503__8_ <= r_n_503__8_;
      r_503__7_ <= r_n_503__7_;
      r_503__6_ <= r_n_503__6_;
      r_503__5_ <= r_n_503__5_;
      r_503__4_ <= r_n_503__4_;
      r_503__3_ <= r_n_503__3_;
      r_503__2_ <= r_n_503__2_;
      r_503__1_ <= r_n_503__1_;
      r_503__0_ <= r_n_503__0_;
    end 
    if(N4088) begin
      r_504__63_ <= r_n_504__63_;
      r_504__62_ <= r_n_504__62_;
      r_504__61_ <= r_n_504__61_;
      r_504__60_ <= r_n_504__60_;
      r_504__59_ <= r_n_504__59_;
      r_504__58_ <= r_n_504__58_;
      r_504__57_ <= r_n_504__57_;
      r_504__56_ <= r_n_504__56_;
      r_504__55_ <= r_n_504__55_;
      r_504__54_ <= r_n_504__54_;
      r_504__53_ <= r_n_504__53_;
      r_504__52_ <= r_n_504__52_;
      r_504__51_ <= r_n_504__51_;
      r_504__50_ <= r_n_504__50_;
      r_504__49_ <= r_n_504__49_;
      r_504__48_ <= r_n_504__48_;
      r_504__47_ <= r_n_504__47_;
      r_504__46_ <= r_n_504__46_;
      r_504__45_ <= r_n_504__45_;
      r_504__44_ <= r_n_504__44_;
      r_504__43_ <= r_n_504__43_;
      r_504__42_ <= r_n_504__42_;
      r_504__41_ <= r_n_504__41_;
      r_504__40_ <= r_n_504__40_;
      r_504__39_ <= r_n_504__39_;
      r_504__38_ <= r_n_504__38_;
      r_504__37_ <= r_n_504__37_;
      r_504__36_ <= r_n_504__36_;
      r_504__35_ <= r_n_504__35_;
      r_504__34_ <= r_n_504__34_;
      r_504__33_ <= r_n_504__33_;
      r_504__32_ <= r_n_504__32_;
      r_504__31_ <= r_n_504__31_;
      r_504__30_ <= r_n_504__30_;
      r_504__29_ <= r_n_504__29_;
      r_504__28_ <= r_n_504__28_;
      r_504__27_ <= r_n_504__27_;
      r_504__26_ <= r_n_504__26_;
      r_504__25_ <= r_n_504__25_;
      r_504__24_ <= r_n_504__24_;
      r_504__23_ <= r_n_504__23_;
      r_504__22_ <= r_n_504__22_;
      r_504__21_ <= r_n_504__21_;
      r_504__20_ <= r_n_504__20_;
      r_504__19_ <= r_n_504__19_;
      r_504__18_ <= r_n_504__18_;
      r_504__17_ <= r_n_504__17_;
      r_504__16_ <= r_n_504__16_;
      r_504__15_ <= r_n_504__15_;
      r_504__14_ <= r_n_504__14_;
      r_504__13_ <= r_n_504__13_;
      r_504__12_ <= r_n_504__12_;
      r_504__11_ <= r_n_504__11_;
      r_504__10_ <= r_n_504__10_;
      r_504__9_ <= r_n_504__9_;
      r_504__8_ <= r_n_504__8_;
      r_504__7_ <= r_n_504__7_;
      r_504__6_ <= r_n_504__6_;
      r_504__5_ <= r_n_504__5_;
      r_504__4_ <= r_n_504__4_;
      r_504__3_ <= r_n_504__3_;
      r_504__2_ <= r_n_504__2_;
      r_504__1_ <= r_n_504__1_;
      r_504__0_ <= r_n_504__0_;
    end 
    if(N4089) begin
      r_505__63_ <= r_n_505__63_;
      r_505__62_ <= r_n_505__62_;
      r_505__61_ <= r_n_505__61_;
      r_505__60_ <= r_n_505__60_;
      r_505__59_ <= r_n_505__59_;
      r_505__58_ <= r_n_505__58_;
      r_505__57_ <= r_n_505__57_;
      r_505__56_ <= r_n_505__56_;
      r_505__55_ <= r_n_505__55_;
      r_505__54_ <= r_n_505__54_;
      r_505__53_ <= r_n_505__53_;
      r_505__52_ <= r_n_505__52_;
      r_505__51_ <= r_n_505__51_;
      r_505__50_ <= r_n_505__50_;
      r_505__49_ <= r_n_505__49_;
      r_505__48_ <= r_n_505__48_;
      r_505__47_ <= r_n_505__47_;
      r_505__46_ <= r_n_505__46_;
      r_505__45_ <= r_n_505__45_;
      r_505__44_ <= r_n_505__44_;
      r_505__43_ <= r_n_505__43_;
      r_505__42_ <= r_n_505__42_;
      r_505__41_ <= r_n_505__41_;
      r_505__40_ <= r_n_505__40_;
      r_505__39_ <= r_n_505__39_;
      r_505__38_ <= r_n_505__38_;
      r_505__37_ <= r_n_505__37_;
      r_505__36_ <= r_n_505__36_;
      r_505__35_ <= r_n_505__35_;
      r_505__34_ <= r_n_505__34_;
      r_505__33_ <= r_n_505__33_;
      r_505__32_ <= r_n_505__32_;
      r_505__31_ <= r_n_505__31_;
      r_505__30_ <= r_n_505__30_;
      r_505__29_ <= r_n_505__29_;
      r_505__28_ <= r_n_505__28_;
      r_505__27_ <= r_n_505__27_;
      r_505__26_ <= r_n_505__26_;
      r_505__25_ <= r_n_505__25_;
      r_505__24_ <= r_n_505__24_;
      r_505__23_ <= r_n_505__23_;
      r_505__22_ <= r_n_505__22_;
      r_505__21_ <= r_n_505__21_;
      r_505__20_ <= r_n_505__20_;
      r_505__19_ <= r_n_505__19_;
      r_505__18_ <= r_n_505__18_;
      r_505__17_ <= r_n_505__17_;
      r_505__16_ <= r_n_505__16_;
      r_505__15_ <= r_n_505__15_;
      r_505__14_ <= r_n_505__14_;
      r_505__13_ <= r_n_505__13_;
      r_505__12_ <= r_n_505__12_;
      r_505__11_ <= r_n_505__11_;
      r_505__10_ <= r_n_505__10_;
      r_505__9_ <= r_n_505__9_;
      r_505__8_ <= r_n_505__8_;
      r_505__7_ <= r_n_505__7_;
      r_505__6_ <= r_n_505__6_;
      r_505__5_ <= r_n_505__5_;
      r_505__4_ <= r_n_505__4_;
      r_505__3_ <= r_n_505__3_;
      r_505__2_ <= r_n_505__2_;
      r_505__1_ <= r_n_505__1_;
      r_505__0_ <= r_n_505__0_;
    end 
    if(N4090) begin
      r_506__63_ <= r_n_506__63_;
      r_506__62_ <= r_n_506__62_;
      r_506__61_ <= r_n_506__61_;
      r_506__60_ <= r_n_506__60_;
      r_506__59_ <= r_n_506__59_;
      r_506__58_ <= r_n_506__58_;
      r_506__57_ <= r_n_506__57_;
      r_506__56_ <= r_n_506__56_;
      r_506__55_ <= r_n_506__55_;
      r_506__54_ <= r_n_506__54_;
      r_506__53_ <= r_n_506__53_;
      r_506__52_ <= r_n_506__52_;
      r_506__51_ <= r_n_506__51_;
      r_506__50_ <= r_n_506__50_;
      r_506__49_ <= r_n_506__49_;
      r_506__48_ <= r_n_506__48_;
      r_506__47_ <= r_n_506__47_;
      r_506__46_ <= r_n_506__46_;
      r_506__45_ <= r_n_506__45_;
      r_506__44_ <= r_n_506__44_;
      r_506__43_ <= r_n_506__43_;
      r_506__42_ <= r_n_506__42_;
      r_506__41_ <= r_n_506__41_;
      r_506__40_ <= r_n_506__40_;
      r_506__39_ <= r_n_506__39_;
      r_506__38_ <= r_n_506__38_;
      r_506__37_ <= r_n_506__37_;
      r_506__36_ <= r_n_506__36_;
      r_506__35_ <= r_n_506__35_;
      r_506__34_ <= r_n_506__34_;
      r_506__33_ <= r_n_506__33_;
      r_506__32_ <= r_n_506__32_;
      r_506__31_ <= r_n_506__31_;
      r_506__30_ <= r_n_506__30_;
      r_506__29_ <= r_n_506__29_;
      r_506__28_ <= r_n_506__28_;
      r_506__27_ <= r_n_506__27_;
      r_506__26_ <= r_n_506__26_;
      r_506__25_ <= r_n_506__25_;
      r_506__24_ <= r_n_506__24_;
      r_506__23_ <= r_n_506__23_;
      r_506__22_ <= r_n_506__22_;
      r_506__21_ <= r_n_506__21_;
      r_506__20_ <= r_n_506__20_;
      r_506__19_ <= r_n_506__19_;
      r_506__18_ <= r_n_506__18_;
      r_506__17_ <= r_n_506__17_;
      r_506__16_ <= r_n_506__16_;
      r_506__15_ <= r_n_506__15_;
      r_506__14_ <= r_n_506__14_;
      r_506__13_ <= r_n_506__13_;
      r_506__12_ <= r_n_506__12_;
      r_506__11_ <= r_n_506__11_;
      r_506__10_ <= r_n_506__10_;
      r_506__9_ <= r_n_506__9_;
      r_506__8_ <= r_n_506__8_;
      r_506__7_ <= r_n_506__7_;
      r_506__6_ <= r_n_506__6_;
      r_506__5_ <= r_n_506__5_;
      r_506__4_ <= r_n_506__4_;
      r_506__3_ <= r_n_506__3_;
      r_506__2_ <= r_n_506__2_;
      r_506__1_ <= r_n_506__1_;
      r_506__0_ <= r_n_506__0_;
    end 
    if(N4091) begin
      r_507__63_ <= r_n_507__63_;
      r_507__62_ <= r_n_507__62_;
      r_507__61_ <= r_n_507__61_;
      r_507__60_ <= r_n_507__60_;
      r_507__59_ <= r_n_507__59_;
      r_507__58_ <= r_n_507__58_;
      r_507__57_ <= r_n_507__57_;
      r_507__56_ <= r_n_507__56_;
      r_507__55_ <= r_n_507__55_;
      r_507__54_ <= r_n_507__54_;
      r_507__53_ <= r_n_507__53_;
      r_507__52_ <= r_n_507__52_;
      r_507__51_ <= r_n_507__51_;
      r_507__50_ <= r_n_507__50_;
      r_507__49_ <= r_n_507__49_;
      r_507__48_ <= r_n_507__48_;
      r_507__47_ <= r_n_507__47_;
      r_507__46_ <= r_n_507__46_;
      r_507__45_ <= r_n_507__45_;
      r_507__44_ <= r_n_507__44_;
      r_507__43_ <= r_n_507__43_;
      r_507__42_ <= r_n_507__42_;
      r_507__41_ <= r_n_507__41_;
      r_507__40_ <= r_n_507__40_;
      r_507__39_ <= r_n_507__39_;
      r_507__38_ <= r_n_507__38_;
      r_507__37_ <= r_n_507__37_;
      r_507__36_ <= r_n_507__36_;
      r_507__35_ <= r_n_507__35_;
      r_507__34_ <= r_n_507__34_;
      r_507__33_ <= r_n_507__33_;
      r_507__32_ <= r_n_507__32_;
      r_507__31_ <= r_n_507__31_;
      r_507__30_ <= r_n_507__30_;
      r_507__29_ <= r_n_507__29_;
      r_507__28_ <= r_n_507__28_;
      r_507__27_ <= r_n_507__27_;
      r_507__26_ <= r_n_507__26_;
      r_507__25_ <= r_n_507__25_;
      r_507__24_ <= r_n_507__24_;
      r_507__23_ <= r_n_507__23_;
      r_507__22_ <= r_n_507__22_;
      r_507__21_ <= r_n_507__21_;
      r_507__20_ <= r_n_507__20_;
      r_507__19_ <= r_n_507__19_;
      r_507__18_ <= r_n_507__18_;
      r_507__17_ <= r_n_507__17_;
      r_507__16_ <= r_n_507__16_;
      r_507__15_ <= r_n_507__15_;
      r_507__14_ <= r_n_507__14_;
      r_507__13_ <= r_n_507__13_;
      r_507__12_ <= r_n_507__12_;
      r_507__11_ <= r_n_507__11_;
      r_507__10_ <= r_n_507__10_;
      r_507__9_ <= r_n_507__9_;
      r_507__8_ <= r_n_507__8_;
      r_507__7_ <= r_n_507__7_;
      r_507__6_ <= r_n_507__6_;
      r_507__5_ <= r_n_507__5_;
      r_507__4_ <= r_n_507__4_;
      r_507__3_ <= r_n_507__3_;
      r_507__2_ <= r_n_507__2_;
      r_507__1_ <= r_n_507__1_;
      r_507__0_ <= r_n_507__0_;
    end 
    if(N4092) begin
      r_508__63_ <= r_n_508__63_;
      r_508__62_ <= r_n_508__62_;
      r_508__61_ <= r_n_508__61_;
      r_508__60_ <= r_n_508__60_;
      r_508__59_ <= r_n_508__59_;
      r_508__58_ <= r_n_508__58_;
      r_508__57_ <= r_n_508__57_;
      r_508__56_ <= r_n_508__56_;
      r_508__55_ <= r_n_508__55_;
      r_508__54_ <= r_n_508__54_;
      r_508__53_ <= r_n_508__53_;
      r_508__52_ <= r_n_508__52_;
      r_508__51_ <= r_n_508__51_;
      r_508__50_ <= r_n_508__50_;
      r_508__49_ <= r_n_508__49_;
      r_508__48_ <= r_n_508__48_;
      r_508__47_ <= r_n_508__47_;
      r_508__46_ <= r_n_508__46_;
      r_508__45_ <= r_n_508__45_;
      r_508__44_ <= r_n_508__44_;
      r_508__43_ <= r_n_508__43_;
      r_508__42_ <= r_n_508__42_;
      r_508__41_ <= r_n_508__41_;
      r_508__40_ <= r_n_508__40_;
      r_508__39_ <= r_n_508__39_;
      r_508__38_ <= r_n_508__38_;
      r_508__37_ <= r_n_508__37_;
      r_508__36_ <= r_n_508__36_;
      r_508__35_ <= r_n_508__35_;
      r_508__34_ <= r_n_508__34_;
      r_508__33_ <= r_n_508__33_;
      r_508__32_ <= r_n_508__32_;
      r_508__31_ <= r_n_508__31_;
      r_508__30_ <= r_n_508__30_;
      r_508__29_ <= r_n_508__29_;
      r_508__28_ <= r_n_508__28_;
      r_508__27_ <= r_n_508__27_;
      r_508__26_ <= r_n_508__26_;
      r_508__25_ <= r_n_508__25_;
      r_508__24_ <= r_n_508__24_;
      r_508__23_ <= r_n_508__23_;
      r_508__22_ <= r_n_508__22_;
      r_508__21_ <= r_n_508__21_;
      r_508__20_ <= r_n_508__20_;
      r_508__19_ <= r_n_508__19_;
      r_508__18_ <= r_n_508__18_;
      r_508__17_ <= r_n_508__17_;
      r_508__16_ <= r_n_508__16_;
      r_508__15_ <= r_n_508__15_;
      r_508__14_ <= r_n_508__14_;
      r_508__13_ <= r_n_508__13_;
      r_508__12_ <= r_n_508__12_;
      r_508__11_ <= r_n_508__11_;
      r_508__10_ <= r_n_508__10_;
      r_508__9_ <= r_n_508__9_;
      r_508__8_ <= r_n_508__8_;
      r_508__7_ <= r_n_508__7_;
      r_508__6_ <= r_n_508__6_;
      r_508__5_ <= r_n_508__5_;
      r_508__4_ <= r_n_508__4_;
      r_508__3_ <= r_n_508__3_;
      r_508__2_ <= r_n_508__2_;
      r_508__1_ <= r_n_508__1_;
      r_508__0_ <= r_n_508__0_;
    end 
    if(N4093) begin
      r_509__63_ <= r_n_509__63_;
      r_509__62_ <= r_n_509__62_;
      r_509__61_ <= r_n_509__61_;
      r_509__60_ <= r_n_509__60_;
      r_509__59_ <= r_n_509__59_;
      r_509__58_ <= r_n_509__58_;
      r_509__57_ <= r_n_509__57_;
      r_509__56_ <= r_n_509__56_;
      r_509__55_ <= r_n_509__55_;
      r_509__54_ <= r_n_509__54_;
      r_509__53_ <= r_n_509__53_;
      r_509__52_ <= r_n_509__52_;
      r_509__51_ <= r_n_509__51_;
      r_509__50_ <= r_n_509__50_;
      r_509__49_ <= r_n_509__49_;
      r_509__48_ <= r_n_509__48_;
      r_509__47_ <= r_n_509__47_;
      r_509__46_ <= r_n_509__46_;
      r_509__45_ <= r_n_509__45_;
      r_509__44_ <= r_n_509__44_;
      r_509__43_ <= r_n_509__43_;
      r_509__42_ <= r_n_509__42_;
      r_509__41_ <= r_n_509__41_;
      r_509__40_ <= r_n_509__40_;
      r_509__39_ <= r_n_509__39_;
      r_509__38_ <= r_n_509__38_;
      r_509__37_ <= r_n_509__37_;
      r_509__36_ <= r_n_509__36_;
      r_509__35_ <= r_n_509__35_;
      r_509__34_ <= r_n_509__34_;
      r_509__33_ <= r_n_509__33_;
      r_509__32_ <= r_n_509__32_;
      r_509__31_ <= r_n_509__31_;
      r_509__30_ <= r_n_509__30_;
      r_509__29_ <= r_n_509__29_;
      r_509__28_ <= r_n_509__28_;
      r_509__27_ <= r_n_509__27_;
      r_509__26_ <= r_n_509__26_;
      r_509__25_ <= r_n_509__25_;
      r_509__24_ <= r_n_509__24_;
      r_509__23_ <= r_n_509__23_;
      r_509__22_ <= r_n_509__22_;
      r_509__21_ <= r_n_509__21_;
      r_509__20_ <= r_n_509__20_;
      r_509__19_ <= r_n_509__19_;
      r_509__18_ <= r_n_509__18_;
      r_509__17_ <= r_n_509__17_;
      r_509__16_ <= r_n_509__16_;
      r_509__15_ <= r_n_509__15_;
      r_509__14_ <= r_n_509__14_;
      r_509__13_ <= r_n_509__13_;
      r_509__12_ <= r_n_509__12_;
      r_509__11_ <= r_n_509__11_;
      r_509__10_ <= r_n_509__10_;
      r_509__9_ <= r_n_509__9_;
      r_509__8_ <= r_n_509__8_;
      r_509__7_ <= r_n_509__7_;
      r_509__6_ <= r_n_509__6_;
      r_509__5_ <= r_n_509__5_;
      r_509__4_ <= r_n_509__4_;
      r_509__3_ <= r_n_509__3_;
      r_509__2_ <= r_n_509__2_;
      r_509__1_ <= r_n_509__1_;
      r_509__0_ <= r_n_509__0_;
    end 
    if(N4094) begin
      r_510__63_ <= r_n_510__63_;
      r_510__62_ <= r_n_510__62_;
      r_510__61_ <= r_n_510__61_;
      r_510__60_ <= r_n_510__60_;
      r_510__59_ <= r_n_510__59_;
      r_510__58_ <= r_n_510__58_;
      r_510__57_ <= r_n_510__57_;
      r_510__56_ <= r_n_510__56_;
      r_510__55_ <= r_n_510__55_;
      r_510__54_ <= r_n_510__54_;
      r_510__53_ <= r_n_510__53_;
      r_510__52_ <= r_n_510__52_;
      r_510__51_ <= r_n_510__51_;
      r_510__50_ <= r_n_510__50_;
      r_510__49_ <= r_n_510__49_;
      r_510__48_ <= r_n_510__48_;
      r_510__47_ <= r_n_510__47_;
      r_510__46_ <= r_n_510__46_;
      r_510__45_ <= r_n_510__45_;
      r_510__44_ <= r_n_510__44_;
      r_510__43_ <= r_n_510__43_;
      r_510__42_ <= r_n_510__42_;
      r_510__41_ <= r_n_510__41_;
      r_510__40_ <= r_n_510__40_;
      r_510__39_ <= r_n_510__39_;
      r_510__38_ <= r_n_510__38_;
      r_510__37_ <= r_n_510__37_;
      r_510__36_ <= r_n_510__36_;
      r_510__35_ <= r_n_510__35_;
      r_510__34_ <= r_n_510__34_;
      r_510__33_ <= r_n_510__33_;
      r_510__32_ <= r_n_510__32_;
      r_510__31_ <= r_n_510__31_;
      r_510__30_ <= r_n_510__30_;
      r_510__29_ <= r_n_510__29_;
      r_510__28_ <= r_n_510__28_;
      r_510__27_ <= r_n_510__27_;
      r_510__26_ <= r_n_510__26_;
      r_510__25_ <= r_n_510__25_;
      r_510__24_ <= r_n_510__24_;
      r_510__23_ <= r_n_510__23_;
      r_510__22_ <= r_n_510__22_;
      r_510__21_ <= r_n_510__21_;
      r_510__20_ <= r_n_510__20_;
      r_510__19_ <= r_n_510__19_;
      r_510__18_ <= r_n_510__18_;
      r_510__17_ <= r_n_510__17_;
      r_510__16_ <= r_n_510__16_;
      r_510__15_ <= r_n_510__15_;
      r_510__14_ <= r_n_510__14_;
      r_510__13_ <= r_n_510__13_;
      r_510__12_ <= r_n_510__12_;
      r_510__11_ <= r_n_510__11_;
      r_510__10_ <= r_n_510__10_;
      r_510__9_ <= r_n_510__9_;
      r_510__8_ <= r_n_510__8_;
      r_510__7_ <= r_n_510__7_;
      r_510__6_ <= r_n_510__6_;
      r_510__5_ <= r_n_510__5_;
      r_510__4_ <= r_n_510__4_;
      r_510__3_ <= r_n_510__3_;
      r_510__2_ <= r_n_510__2_;
      r_510__1_ <= r_n_510__1_;
      r_510__0_ <= r_n_510__0_;
    end 
    if(N4095) begin
      r_511__63_ <= r_n_511__63_;
      r_511__62_ <= r_n_511__62_;
      r_511__61_ <= r_n_511__61_;
      r_511__60_ <= r_n_511__60_;
      r_511__59_ <= r_n_511__59_;
      r_511__58_ <= r_n_511__58_;
      r_511__57_ <= r_n_511__57_;
      r_511__56_ <= r_n_511__56_;
      r_511__55_ <= r_n_511__55_;
      r_511__54_ <= r_n_511__54_;
      r_511__53_ <= r_n_511__53_;
      r_511__52_ <= r_n_511__52_;
      r_511__51_ <= r_n_511__51_;
      r_511__50_ <= r_n_511__50_;
      r_511__49_ <= r_n_511__49_;
      r_511__48_ <= r_n_511__48_;
      r_511__47_ <= r_n_511__47_;
      r_511__46_ <= r_n_511__46_;
      r_511__45_ <= r_n_511__45_;
      r_511__44_ <= r_n_511__44_;
      r_511__43_ <= r_n_511__43_;
      r_511__42_ <= r_n_511__42_;
      r_511__41_ <= r_n_511__41_;
      r_511__40_ <= r_n_511__40_;
      r_511__39_ <= r_n_511__39_;
      r_511__38_ <= r_n_511__38_;
      r_511__37_ <= r_n_511__37_;
      r_511__36_ <= r_n_511__36_;
      r_511__35_ <= r_n_511__35_;
      r_511__34_ <= r_n_511__34_;
      r_511__33_ <= r_n_511__33_;
      r_511__32_ <= r_n_511__32_;
      r_511__31_ <= r_n_511__31_;
      r_511__30_ <= r_n_511__30_;
      r_511__29_ <= r_n_511__29_;
      r_511__28_ <= r_n_511__28_;
      r_511__27_ <= r_n_511__27_;
      r_511__26_ <= r_n_511__26_;
      r_511__25_ <= r_n_511__25_;
      r_511__24_ <= r_n_511__24_;
      r_511__23_ <= r_n_511__23_;
      r_511__22_ <= r_n_511__22_;
      r_511__21_ <= r_n_511__21_;
      r_511__20_ <= r_n_511__20_;
      r_511__19_ <= r_n_511__19_;
      r_511__18_ <= r_n_511__18_;
      r_511__17_ <= r_n_511__17_;
      r_511__16_ <= r_n_511__16_;
      r_511__15_ <= r_n_511__15_;
      r_511__14_ <= r_n_511__14_;
      r_511__13_ <= r_n_511__13_;
      r_511__12_ <= r_n_511__12_;
      r_511__11_ <= r_n_511__11_;
      r_511__10_ <= r_n_511__10_;
      r_511__9_ <= r_n_511__9_;
      r_511__8_ <= r_n_511__8_;
      r_511__7_ <= r_n_511__7_;
      r_511__6_ <= r_n_511__6_;
      r_511__5_ <= r_n_511__5_;
      r_511__4_ <= r_n_511__4_;
      r_511__3_ <= r_n_511__3_;
      r_511__2_ <= r_n_511__2_;
      r_511__1_ <= r_n_511__1_;
      r_511__0_ <= r_n_511__0_;
    end 
  end


endmodule

