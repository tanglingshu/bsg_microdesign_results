

module top
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  yumi_o,
  v_o,
  data_o,
  tag_o,
  yumi_i
);

  input [4095:0] data_i;
  input [31:0] v_i;
  output [31:0] yumi_o;
  output [127:0] data_o;
  output [4:0] tag_o;
  input clk_i;
  input reset_i;
  input yumi_i;
  output v_o;

  bsg_round_robin_n_to_1
  wrapper
  (
    .data_i(data_i),
    .v_i(v_i),
    .yumi_o(yumi_o),
    .data_o(data_o),
    .tag_o(tag_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .yumi_i(yumi_i),
    .v_o(v_o)
  );


endmodule



module bsg_circular_ptr_slots_p32_max_add_p1
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [0:0] add_i;
  output [4:0] o;
  output [4:0] n_o;
  input clk;
  input reset_i;
  wire [4:0] n_o,genblk1_genblk1_ptr_r_p1;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;
  reg [4:0] o;
  assign genblk1_genblk1_ptr_r_p1 = o + 1'b1;
  assign { N9, N8, N7, N6, N5 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N1)? n_o : 1'b0;
  assign N0 = reset_i;
  assign N1 = N4;
  assign n_o = (N2)? genblk1_genblk1_ptr_r_p1 : 
               (N3)? o : 1'b0;
  assign N2 = add_i[0];
  assign N3 = N10;
  assign N4 = ~reset_i;
  assign N10 = ~add_i[0];

  always @(posedge clk) begin
    if(1'b1) begin
      { o[4:0] } <= { N9, N8, N7, N6, N5 };
    end 
  end


endmodule



module bsg_round_robin_n_to_1
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  yumi_o,
  v_o,
  data_o,
  tag_o,
  yumi_i
);

  input [4095:0] data_i;
  input [31:0] v_i;
  output [31:0] yumi_o;
  output [127:0] data_o;
  output [4:0] tag_o;
  input clk_i;
  input reset_i;
  input yumi_i;
  output v_o;
  wire [31:0] yumi_o;
  wire [127:0] data_o;
  wire [4:0] tag_o;
  wire v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,
  N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,
  N117,N118,N119,N120,N121,N122,N123,N124,SYNOPSYS_UNCONNECTED_1,
  SYNOPSYS_UNCONNECTED_2,SYNOPSYS_UNCONNECTED_3,SYNOPSYS_UNCONNECTED_4,SYNOPSYS_UNCONNECTED_5;

  bsg_circular_ptr_slots_p32_max_add_p1
  strict_circular_ptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(yumi_i),
    .o(tag_o),
    .n_o({ SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5 })
  );

  assign v_o = (N33)? v_i[0] : 
               (N35)? v_i[1] : 
               (N37)? v_i[2] : 
               (N39)? v_i[3] : 
               (N41)? v_i[4] : 
               (N43)? v_i[5] : 
               (N45)? v_i[6] : 
               (N47)? v_i[7] : 
               (N49)? v_i[8] : 
               (N51)? v_i[9] : 
               (N53)? v_i[10] : 
               (N55)? v_i[11] : 
               (N57)? v_i[12] : 
               (N59)? v_i[13] : 
               (N61)? v_i[14] : 
               (N63)? v_i[15] : 
               (N34)? v_i[16] : 
               (N36)? v_i[17] : 
               (N38)? v_i[18] : 
               (N40)? v_i[19] : 
               (N42)? v_i[20] : 
               (N44)? v_i[21] : 
               (N46)? v_i[22] : 
               (N48)? v_i[23] : 
               (N50)? v_i[24] : 
               (N52)? v_i[25] : 
               (N54)? v_i[26] : 
               (N56)? v_i[27] : 
               (N58)? v_i[28] : 
               (N60)? v_i[29] : 
               (N62)? v_i[30] : 
               (N64)? v_i[31] : 1'b0;
  assign data_o[127] = (N93)? data_i[127] : 
                       (N95)? data_i[255] : 
                       (N97)? data_i[383] : 
                       (N99)? data_i[511] : 
                       (N101)? data_i[639] : 
                       (N103)? data_i[767] : 
                       (N105)? data_i[895] : 
                       (N107)? data_i[1023] : 
                       (N109)? data_i[1151] : 
                       (N111)? data_i[1279] : 
                       (N113)? data_i[1407] : 
                       (N115)? data_i[1535] : 
                       (N117)? data_i[1663] : 
                       (N119)? data_i[1791] : 
                       (N121)? data_i[1919] : 
                       (N123)? data_i[2047] : 
                       (N94)? data_i[2175] : 
                       (N96)? data_i[2303] : 
                       (N98)? data_i[2431] : 
                       (N100)? data_i[2559] : 
                       (N102)? data_i[2687] : 
                       (N104)? data_i[2815] : 
                       (N106)? data_i[2943] : 
                       (N108)? data_i[3071] : 
                       (N110)? data_i[3199] : 
                       (N112)? data_i[3327] : 
                       (N114)? data_i[3455] : 
                       (N116)? data_i[3583] : 
                       (N118)? data_i[3711] : 
                       (N120)? data_i[3839] : 
                       (N122)? data_i[3967] : 
                       (N124)? data_i[4095] : 1'b0;
  assign data_o[126] = (N93)? data_i[126] : 
                       (N95)? data_i[254] : 
                       (N97)? data_i[382] : 
                       (N99)? data_i[510] : 
                       (N101)? data_i[638] : 
                       (N103)? data_i[766] : 
                       (N105)? data_i[894] : 
                       (N107)? data_i[1022] : 
                       (N109)? data_i[1150] : 
                       (N111)? data_i[1278] : 
                       (N113)? data_i[1406] : 
                       (N115)? data_i[1534] : 
                       (N117)? data_i[1662] : 
                       (N119)? data_i[1790] : 
                       (N121)? data_i[1918] : 
                       (N123)? data_i[2046] : 
                       (N94)? data_i[2174] : 
                       (N96)? data_i[2302] : 
                       (N98)? data_i[2430] : 
                       (N100)? data_i[2558] : 
                       (N102)? data_i[2686] : 
                       (N104)? data_i[2814] : 
                       (N106)? data_i[2942] : 
                       (N108)? data_i[3070] : 
                       (N110)? data_i[3198] : 
                       (N112)? data_i[3326] : 
                       (N114)? data_i[3454] : 
                       (N116)? data_i[3582] : 
                       (N118)? data_i[3710] : 
                       (N120)? data_i[3838] : 
                       (N122)? data_i[3966] : 
                       (N124)? data_i[4094] : 1'b0;
  assign data_o[125] = (N93)? data_i[125] : 
                       (N95)? data_i[253] : 
                       (N97)? data_i[381] : 
                       (N99)? data_i[509] : 
                       (N101)? data_i[637] : 
                       (N103)? data_i[765] : 
                       (N105)? data_i[893] : 
                       (N107)? data_i[1021] : 
                       (N109)? data_i[1149] : 
                       (N111)? data_i[1277] : 
                       (N113)? data_i[1405] : 
                       (N115)? data_i[1533] : 
                       (N117)? data_i[1661] : 
                       (N119)? data_i[1789] : 
                       (N121)? data_i[1917] : 
                       (N123)? data_i[2045] : 
                       (N94)? data_i[2173] : 
                       (N96)? data_i[2301] : 
                       (N98)? data_i[2429] : 
                       (N100)? data_i[2557] : 
                       (N102)? data_i[2685] : 
                       (N104)? data_i[2813] : 
                       (N106)? data_i[2941] : 
                       (N108)? data_i[3069] : 
                       (N110)? data_i[3197] : 
                       (N112)? data_i[3325] : 
                       (N114)? data_i[3453] : 
                       (N116)? data_i[3581] : 
                       (N118)? data_i[3709] : 
                       (N120)? data_i[3837] : 
                       (N122)? data_i[3965] : 
                       (N124)? data_i[4093] : 1'b0;
  assign data_o[124] = (N93)? data_i[124] : 
                       (N95)? data_i[252] : 
                       (N97)? data_i[380] : 
                       (N99)? data_i[508] : 
                       (N101)? data_i[636] : 
                       (N103)? data_i[764] : 
                       (N105)? data_i[892] : 
                       (N107)? data_i[1020] : 
                       (N109)? data_i[1148] : 
                       (N111)? data_i[1276] : 
                       (N113)? data_i[1404] : 
                       (N115)? data_i[1532] : 
                       (N117)? data_i[1660] : 
                       (N119)? data_i[1788] : 
                       (N121)? data_i[1916] : 
                       (N123)? data_i[2044] : 
                       (N94)? data_i[2172] : 
                       (N96)? data_i[2300] : 
                       (N98)? data_i[2428] : 
                       (N100)? data_i[2556] : 
                       (N102)? data_i[2684] : 
                       (N104)? data_i[2812] : 
                       (N106)? data_i[2940] : 
                       (N108)? data_i[3068] : 
                       (N110)? data_i[3196] : 
                       (N112)? data_i[3324] : 
                       (N114)? data_i[3452] : 
                       (N116)? data_i[3580] : 
                       (N118)? data_i[3708] : 
                       (N120)? data_i[3836] : 
                       (N122)? data_i[3964] : 
                       (N124)? data_i[4092] : 1'b0;
  assign data_o[123] = (N93)? data_i[123] : 
                       (N95)? data_i[251] : 
                       (N97)? data_i[379] : 
                       (N99)? data_i[507] : 
                       (N101)? data_i[635] : 
                       (N103)? data_i[763] : 
                       (N105)? data_i[891] : 
                       (N107)? data_i[1019] : 
                       (N109)? data_i[1147] : 
                       (N111)? data_i[1275] : 
                       (N113)? data_i[1403] : 
                       (N115)? data_i[1531] : 
                       (N117)? data_i[1659] : 
                       (N119)? data_i[1787] : 
                       (N121)? data_i[1915] : 
                       (N123)? data_i[2043] : 
                       (N94)? data_i[2171] : 
                       (N96)? data_i[2299] : 
                       (N98)? data_i[2427] : 
                       (N100)? data_i[2555] : 
                       (N102)? data_i[2683] : 
                       (N104)? data_i[2811] : 
                       (N106)? data_i[2939] : 
                       (N108)? data_i[3067] : 
                       (N110)? data_i[3195] : 
                       (N112)? data_i[3323] : 
                       (N114)? data_i[3451] : 
                       (N116)? data_i[3579] : 
                       (N118)? data_i[3707] : 
                       (N120)? data_i[3835] : 
                       (N122)? data_i[3963] : 
                       (N124)? data_i[4091] : 1'b0;
  assign data_o[122] = (N93)? data_i[122] : 
                       (N95)? data_i[250] : 
                       (N97)? data_i[378] : 
                       (N99)? data_i[506] : 
                       (N101)? data_i[634] : 
                       (N103)? data_i[762] : 
                       (N105)? data_i[890] : 
                       (N107)? data_i[1018] : 
                       (N109)? data_i[1146] : 
                       (N111)? data_i[1274] : 
                       (N113)? data_i[1402] : 
                       (N115)? data_i[1530] : 
                       (N117)? data_i[1658] : 
                       (N119)? data_i[1786] : 
                       (N121)? data_i[1914] : 
                       (N123)? data_i[2042] : 
                       (N94)? data_i[2170] : 
                       (N96)? data_i[2298] : 
                       (N98)? data_i[2426] : 
                       (N100)? data_i[2554] : 
                       (N102)? data_i[2682] : 
                       (N104)? data_i[2810] : 
                       (N106)? data_i[2938] : 
                       (N108)? data_i[3066] : 
                       (N110)? data_i[3194] : 
                       (N112)? data_i[3322] : 
                       (N114)? data_i[3450] : 
                       (N116)? data_i[3578] : 
                       (N118)? data_i[3706] : 
                       (N120)? data_i[3834] : 
                       (N122)? data_i[3962] : 
                       (N124)? data_i[4090] : 1'b0;
  assign data_o[121] = (N93)? data_i[121] : 
                       (N95)? data_i[249] : 
                       (N97)? data_i[377] : 
                       (N99)? data_i[505] : 
                       (N101)? data_i[633] : 
                       (N103)? data_i[761] : 
                       (N105)? data_i[889] : 
                       (N107)? data_i[1017] : 
                       (N109)? data_i[1145] : 
                       (N111)? data_i[1273] : 
                       (N113)? data_i[1401] : 
                       (N115)? data_i[1529] : 
                       (N117)? data_i[1657] : 
                       (N119)? data_i[1785] : 
                       (N121)? data_i[1913] : 
                       (N123)? data_i[2041] : 
                       (N94)? data_i[2169] : 
                       (N96)? data_i[2297] : 
                       (N98)? data_i[2425] : 
                       (N100)? data_i[2553] : 
                       (N102)? data_i[2681] : 
                       (N104)? data_i[2809] : 
                       (N106)? data_i[2937] : 
                       (N108)? data_i[3065] : 
                       (N110)? data_i[3193] : 
                       (N112)? data_i[3321] : 
                       (N114)? data_i[3449] : 
                       (N116)? data_i[3577] : 
                       (N118)? data_i[3705] : 
                       (N120)? data_i[3833] : 
                       (N122)? data_i[3961] : 
                       (N124)? data_i[4089] : 1'b0;
  assign data_o[120] = (N93)? data_i[120] : 
                       (N95)? data_i[248] : 
                       (N97)? data_i[376] : 
                       (N99)? data_i[504] : 
                       (N101)? data_i[632] : 
                       (N103)? data_i[760] : 
                       (N105)? data_i[888] : 
                       (N107)? data_i[1016] : 
                       (N109)? data_i[1144] : 
                       (N111)? data_i[1272] : 
                       (N113)? data_i[1400] : 
                       (N115)? data_i[1528] : 
                       (N117)? data_i[1656] : 
                       (N119)? data_i[1784] : 
                       (N121)? data_i[1912] : 
                       (N123)? data_i[2040] : 
                       (N94)? data_i[2168] : 
                       (N96)? data_i[2296] : 
                       (N98)? data_i[2424] : 
                       (N100)? data_i[2552] : 
                       (N102)? data_i[2680] : 
                       (N104)? data_i[2808] : 
                       (N106)? data_i[2936] : 
                       (N108)? data_i[3064] : 
                       (N110)? data_i[3192] : 
                       (N112)? data_i[3320] : 
                       (N114)? data_i[3448] : 
                       (N116)? data_i[3576] : 
                       (N118)? data_i[3704] : 
                       (N120)? data_i[3832] : 
                       (N122)? data_i[3960] : 
                       (N124)? data_i[4088] : 1'b0;
  assign data_o[119] = (N93)? data_i[119] : 
                       (N95)? data_i[247] : 
                       (N97)? data_i[375] : 
                       (N99)? data_i[503] : 
                       (N101)? data_i[631] : 
                       (N103)? data_i[759] : 
                       (N105)? data_i[887] : 
                       (N107)? data_i[1015] : 
                       (N109)? data_i[1143] : 
                       (N111)? data_i[1271] : 
                       (N113)? data_i[1399] : 
                       (N115)? data_i[1527] : 
                       (N117)? data_i[1655] : 
                       (N119)? data_i[1783] : 
                       (N121)? data_i[1911] : 
                       (N123)? data_i[2039] : 
                       (N94)? data_i[2167] : 
                       (N96)? data_i[2295] : 
                       (N98)? data_i[2423] : 
                       (N100)? data_i[2551] : 
                       (N102)? data_i[2679] : 
                       (N104)? data_i[2807] : 
                       (N106)? data_i[2935] : 
                       (N108)? data_i[3063] : 
                       (N110)? data_i[3191] : 
                       (N112)? data_i[3319] : 
                       (N114)? data_i[3447] : 
                       (N116)? data_i[3575] : 
                       (N118)? data_i[3703] : 
                       (N120)? data_i[3831] : 
                       (N122)? data_i[3959] : 
                       (N124)? data_i[4087] : 1'b0;
  assign data_o[118] = (N93)? data_i[118] : 
                       (N95)? data_i[246] : 
                       (N97)? data_i[374] : 
                       (N99)? data_i[502] : 
                       (N101)? data_i[630] : 
                       (N103)? data_i[758] : 
                       (N105)? data_i[886] : 
                       (N107)? data_i[1014] : 
                       (N109)? data_i[1142] : 
                       (N111)? data_i[1270] : 
                       (N113)? data_i[1398] : 
                       (N115)? data_i[1526] : 
                       (N117)? data_i[1654] : 
                       (N119)? data_i[1782] : 
                       (N121)? data_i[1910] : 
                       (N123)? data_i[2038] : 
                       (N94)? data_i[2166] : 
                       (N96)? data_i[2294] : 
                       (N98)? data_i[2422] : 
                       (N100)? data_i[2550] : 
                       (N102)? data_i[2678] : 
                       (N104)? data_i[2806] : 
                       (N106)? data_i[2934] : 
                       (N108)? data_i[3062] : 
                       (N110)? data_i[3190] : 
                       (N112)? data_i[3318] : 
                       (N114)? data_i[3446] : 
                       (N116)? data_i[3574] : 
                       (N118)? data_i[3702] : 
                       (N120)? data_i[3830] : 
                       (N122)? data_i[3958] : 
                       (N124)? data_i[4086] : 1'b0;
  assign data_o[117] = (N93)? data_i[117] : 
                       (N95)? data_i[245] : 
                       (N97)? data_i[373] : 
                       (N99)? data_i[501] : 
                       (N101)? data_i[629] : 
                       (N103)? data_i[757] : 
                       (N105)? data_i[885] : 
                       (N107)? data_i[1013] : 
                       (N109)? data_i[1141] : 
                       (N111)? data_i[1269] : 
                       (N113)? data_i[1397] : 
                       (N115)? data_i[1525] : 
                       (N117)? data_i[1653] : 
                       (N119)? data_i[1781] : 
                       (N121)? data_i[1909] : 
                       (N123)? data_i[2037] : 
                       (N94)? data_i[2165] : 
                       (N96)? data_i[2293] : 
                       (N98)? data_i[2421] : 
                       (N100)? data_i[2549] : 
                       (N102)? data_i[2677] : 
                       (N104)? data_i[2805] : 
                       (N106)? data_i[2933] : 
                       (N108)? data_i[3061] : 
                       (N110)? data_i[3189] : 
                       (N112)? data_i[3317] : 
                       (N114)? data_i[3445] : 
                       (N116)? data_i[3573] : 
                       (N118)? data_i[3701] : 
                       (N120)? data_i[3829] : 
                       (N122)? data_i[3957] : 
                       (N124)? data_i[4085] : 1'b0;
  assign data_o[116] = (N93)? data_i[116] : 
                       (N95)? data_i[244] : 
                       (N97)? data_i[372] : 
                       (N99)? data_i[500] : 
                       (N101)? data_i[628] : 
                       (N103)? data_i[756] : 
                       (N105)? data_i[884] : 
                       (N107)? data_i[1012] : 
                       (N109)? data_i[1140] : 
                       (N111)? data_i[1268] : 
                       (N113)? data_i[1396] : 
                       (N115)? data_i[1524] : 
                       (N117)? data_i[1652] : 
                       (N119)? data_i[1780] : 
                       (N121)? data_i[1908] : 
                       (N123)? data_i[2036] : 
                       (N94)? data_i[2164] : 
                       (N96)? data_i[2292] : 
                       (N98)? data_i[2420] : 
                       (N100)? data_i[2548] : 
                       (N102)? data_i[2676] : 
                       (N104)? data_i[2804] : 
                       (N106)? data_i[2932] : 
                       (N108)? data_i[3060] : 
                       (N110)? data_i[3188] : 
                       (N112)? data_i[3316] : 
                       (N114)? data_i[3444] : 
                       (N116)? data_i[3572] : 
                       (N118)? data_i[3700] : 
                       (N120)? data_i[3828] : 
                       (N122)? data_i[3956] : 
                       (N124)? data_i[4084] : 1'b0;
  assign data_o[115] = (N93)? data_i[115] : 
                       (N95)? data_i[243] : 
                       (N97)? data_i[371] : 
                       (N99)? data_i[499] : 
                       (N101)? data_i[627] : 
                       (N103)? data_i[755] : 
                       (N105)? data_i[883] : 
                       (N107)? data_i[1011] : 
                       (N109)? data_i[1139] : 
                       (N111)? data_i[1267] : 
                       (N113)? data_i[1395] : 
                       (N115)? data_i[1523] : 
                       (N117)? data_i[1651] : 
                       (N119)? data_i[1779] : 
                       (N121)? data_i[1907] : 
                       (N123)? data_i[2035] : 
                       (N94)? data_i[2163] : 
                       (N96)? data_i[2291] : 
                       (N98)? data_i[2419] : 
                       (N100)? data_i[2547] : 
                       (N102)? data_i[2675] : 
                       (N104)? data_i[2803] : 
                       (N106)? data_i[2931] : 
                       (N108)? data_i[3059] : 
                       (N110)? data_i[3187] : 
                       (N112)? data_i[3315] : 
                       (N114)? data_i[3443] : 
                       (N116)? data_i[3571] : 
                       (N118)? data_i[3699] : 
                       (N120)? data_i[3827] : 
                       (N122)? data_i[3955] : 
                       (N124)? data_i[4083] : 1'b0;
  assign data_o[114] = (N93)? data_i[114] : 
                       (N95)? data_i[242] : 
                       (N97)? data_i[370] : 
                       (N99)? data_i[498] : 
                       (N101)? data_i[626] : 
                       (N103)? data_i[754] : 
                       (N105)? data_i[882] : 
                       (N107)? data_i[1010] : 
                       (N109)? data_i[1138] : 
                       (N111)? data_i[1266] : 
                       (N113)? data_i[1394] : 
                       (N115)? data_i[1522] : 
                       (N117)? data_i[1650] : 
                       (N119)? data_i[1778] : 
                       (N121)? data_i[1906] : 
                       (N123)? data_i[2034] : 
                       (N94)? data_i[2162] : 
                       (N96)? data_i[2290] : 
                       (N98)? data_i[2418] : 
                       (N100)? data_i[2546] : 
                       (N102)? data_i[2674] : 
                       (N104)? data_i[2802] : 
                       (N106)? data_i[2930] : 
                       (N108)? data_i[3058] : 
                       (N110)? data_i[3186] : 
                       (N112)? data_i[3314] : 
                       (N114)? data_i[3442] : 
                       (N116)? data_i[3570] : 
                       (N118)? data_i[3698] : 
                       (N120)? data_i[3826] : 
                       (N122)? data_i[3954] : 
                       (N124)? data_i[4082] : 1'b0;
  assign data_o[113] = (N93)? data_i[113] : 
                       (N95)? data_i[241] : 
                       (N97)? data_i[369] : 
                       (N99)? data_i[497] : 
                       (N101)? data_i[625] : 
                       (N103)? data_i[753] : 
                       (N105)? data_i[881] : 
                       (N107)? data_i[1009] : 
                       (N109)? data_i[1137] : 
                       (N111)? data_i[1265] : 
                       (N113)? data_i[1393] : 
                       (N115)? data_i[1521] : 
                       (N117)? data_i[1649] : 
                       (N119)? data_i[1777] : 
                       (N121)? data_i[1905] : 
                       (N123)? data_i[2033] : 
                       (N94)? data_i[2161] : 
                       (N96)? data_i[2289] : 
                       (N98)? data_i[2417] : 
                       (N100)? data_i[2545] : 
                       (N102)? data_i[2673] : 
                       (N104)? data_i[2801] : 
                       (N106)? data_i[2929] : 
                       (N108)? data_i[3057] : 
                       (N110)? data_i[3185] : 
                       (N112)? data_i[3313] : 
                       (N114)? data_i[3441] : 
                       (N116)? data_i[3569] : 
                       (N118)? data_i[3697] : 
                       (N120)? data_i[3825] : 
                       (N122)? data_i[3953] : 
                       (N124)? data_i[4081] : 1'b0;
  assign data_o[112] = (N93)? data_i[112] : 
                       (N95)? data_i[240] : 
                       (N97)? data_i[368] : 
                       (N99)? data_i[496] : 
                       (N101)? data_i[624] : 
                       (N103)? data_i[752] : 
                       (N105)? data_i[880] : 
                       (N107)? data_i[1008] : 
                       (N109)? data_i[1136] : 
                       (N111)? data_i[1264] : 
                       (N113)? data_i[1392] : 
                       (N115)? data_i[1520] : 
                       (N117)? data_i[1648] : 
                       (N119)? data_i[1776] : 
                       (N121)? data_i[1904] : 
                       (N123)? data_i[2032] : 
                       (N94)? data_i[2160] : 
                       (N96)? data_i[2288] : 
                       (N98)? data_i[2416] : 
                       (N100)? data_i[2544] : 
                       (N102)? data_i[2672] : 
                       (N104)? data_i[2800] : 
                       (N106)? data_i[2928] : 
                       (N108)? data_i[3056] : 
                       (N110)? data_i[3184] : 
                       (N112)? data_i[3312] : 
                       (N114)? data_i[3440] : 
                       (N116)? data_i[3568] : 
                       (N118)? data_i[3696] : 
                       (N120)? data_i[3824] : 
                       (N122)? data_i[3952] : 
                       (N124)? data_i[4080] : 1'b0;
  assign data_o[111] = (N93)? data_i[111] : 
                       (N95)? data_i[239] : 
                       (N97)? data_i[367] : 
                       (N99)? data_i[495] : 
                       (N101)? data_i[623] : 
                       (N103)? data_i[751] : 
                       (N105)? data_i[879] : 
                       (N107)? data_i[1007] : 
                       (N109)? data_i[1135] : 
                       (N111)? data_i[1263] : 
                       (N113)? data_i[1391] : 
                       (N115)? data_i[1519] : 
                       (N117)? data_i[1647] : 
                       (N119)? data_i[1775] : 
                       (N121)? data_i[1903] : 
                       (N123)? data_i[2031] : 
                       (N94)? data_i[2159] : 
                       (N96)? data_i[2287] : 
                       (N98)? data_i[2415] : 
                       (N100)? data_i[2543] : 
                       (N102)? data_i[2671] : 
                       (N104)? data_i[2799] : 
                       (N106)? data_i[2927] : 
                       (N108)? data_i[3055] : 
                       (N110)? data_i[3183] : 
                       (N112)? data_i[3311] : 
                       (N114)? data_i[3439] : 
                       (N116)? data_i[3567] : 
                       (N118)? data_i[3695] : 
                       (N120)? data_i[3823] : 
                       (N122)? data_i[3951] : 
                       (N124)? data_i[4079] : 1'b0;
  assign data_o[110] = (N93)? data_i[110] : 
                       (N95)? data_i[238] : 
                       (N97)? data_i[366] : 
                       (N99)? data_i[494] : 
                       (N101)? data_i[622] : 
                       (N103)? data_i[750] : 
                       (N105)? data_i[878] : 
                       (N107)? data_i[1006] : 
                       (N109)? data_i[1134] : 
                       (N111)? data_i[1262] : 
                       (N113)? data_i[1390] : 
                       (N115)? data_i[1518] : 
                       (N117)? data_i[1646] : 
                       (N119)? data_i[1774] : 
                       (N121)? data_i[1902] : 
                       (N123)? data_i[2030] : 
                       (N94)? data_i[2158] : 
                       (N96)? data_i[2286] : 
                       (N98)? data_i[2414] : 
                       (N100)? data_i[2542] : 
                       (N102)? data_i[2670] : 
                       (N104)? data_i[2798] : 
                       (N106)? data_i[2926] : 
                       (N108)? data_i[3054] : 
                       (N110)? data_i[3182] : 
                       (N112)? data_i[3310] : 
                       (N114)? data_i[3438] : 
                       (N116)? data_i[3566] : 
                       (N118)? data_i[3694] : 
                       (N120)? data_i[3822] : 
                       (N122)? data_i[3950] : 
                       (N124)? data_i[4078] : 1'b0;
  assign data_o[109] = (N93)? data_i[109] : 
                       (N95)? data_i[237] : 
                       (N97)? data_i[365] : 
                       (N99)? data_i[493] : 
                       (N101)? data_i[621] : 
                       (N103)? data_i[749] : 
                       (N105)? data_i[877] : 
                       (N107)? data_i[1005] : 
                       (N109)? data_i[1133] : 
                       (N111)? data_i[1261] : 
                       (N113)? data_i[1389] : 
                       (N115)? data_i[1517] : 
                       (N117)? data_i[1645] : 
                       (N119)? data_i[1773] : 
                       (N121)? data_i[1901] : 
                       (N123)? data_i[2029] : 
                       (N94)? data_i[2157] : 
                       (N96)? data_i[2285] : 
                       (N98)? data_i[2413] : 
                       (N100)? data_i[2541] : 
                       (N102)? data_i[2669] : 
                       (N104)? data_i[2797] : 
                       (N106)? data_i[2925] : 
                       (N108)? data_i[3053] : 
                       (N110)? data_i[3181] : 
                       (N112)? data_i[3309] : 
                       (N114)? data_i[3437] : 
                       (N116)? data_i[3565] : 
                       (N118)? data_i[3693] : 
                       (N120)? data_i[3821] : 
                       (N122)? data_i[3949] : 
                       (N124)? data_i[4077] : 1'b0;
  assign data_o[108] = (N93)? data_i[108] : 
                       (N95)? data_i[236] : 
                       (N97)? data_i[364] : 
                       (N99)? data_i[492] : 
                       (N101)? data_i[620] : 
                       (N103)? data_i[748] : 
                       (N105)? data_i[876] : 
                       (N107)? data_i[1004] : 
                       (N109)? data_i[1132] : 
                       (N111)? data_i[1260] : 
                       (N113)? data_i[1388] : 
                       (N115)? data_i[1516] : 
                       (N117)? data_i[1644] : 
                       (N119)? data_i[1772] : 
                       (N121)? data_i[1900] : 
                       (N123)? data_i[2028] : 
                       (N94)? data_i[2156] : 
                       (N96)? data_i[2284] : 
                       (N98)? data_i[2412] : 
                       (N100)? data_i[2540] : 
                       (N102)? data_i[2668] : 
                       (N104)? data_i[2796] : 
                       (N106)? data_i[2924] : 
                       (N108)? data_i[3052] : 
                       (N110)? data_i[3180] : 
                       (N112)? data_i[3308] : 
                       (N114)? data_i[3436] : 
                       (N116)? data_i[3564] : 
                       (N118)? data_i[3692] : 
                       (N120)? data_i[3820] : 
                       (N122)? data_i[3948] : 
                       (N124)? data_i[4076] : 1'b0;
  assign data_o[107] = (N93)? data_i[107] : 
                       (N95)? data_i[235] : 
                       (N97)? data_i[363] : 
                       (N99)? data_i[491] : 
                       (N101)? data_i[619] : 
                       (N103)? data_i[747] : 
                       (N105)? data_i[875] : 
                       (N107)? data_i[1003] : 
                       (N109)? data_i[1131] : 
                       (N111)? data_i[1259] : 
                       (N113)? data_i[1387] : 
                       (N115)? data_i[1515] : 
                       (N117)? data_i[1643] : 
                       (N119)? data_i[1771] : 
                       (N121)? data_i[1899] : 
                       (N123)? data_i[2027] : 
                       (N94)? data_i[2155] : 
                       (N96)? data_i[2283] : 
                       (N98)? data_i[2411] : 
                       (N100)? data_i[2539] : 
                       (N102)? data_i[2667] : 
                       (N104)? data_i[2795] : 
                       (N106)? data_i[2923] : 
                       (N108)? data_i[3051] : 
                       (N110)? data_i[3179] : 
                       (N112)? data_i[3307] : 
                       (N114)? data_i[3435] : 
                       (N116)? data_i[3563] : 
                       (N118)? data_i[3691] : 
                       (N120)? data_i[3819] : 
                       (N122)? data_i[3947] : 
                       (N124)? data_i[4075] : 1'b0;
  assign data_o[106] = (N93)? data_i[106] : 
                       (N95)? data_i[234] : 
                       (N97)? data_i[362] : 
                       (N99)? data_i[490] : 
                       (N101)? data_i[618] : 
                       (N103)? data_i[746] : 
                       (N105)? data_i[874] : 
                       (N107)? data_i[1002] : 
                       (N109)? data_i[1130] : 
                       (N111)? data_i[1258] : 
                       (N113)? data_i[1386] : 
                       (N115)? data_i[1514] : 
                       (N117)? data_i[1642] : 
                       (N119)? data_i[1770] : 
                       (N121)? data_i[1898] : 
                       (N123)? data_i[2026] : 
                       (N94)? data_i[2154] : 
                       (N96)? data_i[2282] : 
                       (N98)? data_i[2410] : 
                       (N100)? data_i[2538] : 
                       (N102)? data_i[2666] : 
                       (N104)? data_i[2794] : 
                       (N106)? data_i[2922] : 
                       (N108)? data_i[3050] : 
                       (N110)? data_i[3178] : 
                       (N112)? data_i[3306] : 
                       (N114)? data_i[3434] : 
                       (N116)? data_i[3562] : 
                       (N118)? data_i[3690] : 
                       (N120)? data_i[3818] : 
                       (N122)? data_i[3946] : 
                       (N124)? data_i[4074] : 1'b0;
  assign data_o[105] = (N93)? data_i[105] : 
                       (N95)? data_i[233] : 
                       (N97)? data_i[361] : 
                       (N99)? data_i[489] : 
                       (N101)? data_i[617] : 
                       (N103)? data_i[745] : 
                       (N105)? data_i[873] : 
                       (N107)? data_i[1001] : 
                       (N109)? data_i[1129] : 
                       (N111)? data_i[1257] : 
                       (N113)? data_i[1385] : 
                       (N115)? data_i[1513] : 
                       (N117)? data_i[1641] : 
                       (N119)? data_i[1769] : 
                       (N121)? data_i[1897] : 
                       (N123)? data_i[2025] : 
                       (N94)? data_i[2153] : 
                       (N96)? data_i[2281] : 
                       (N98)? data_i[2409] : 
                       (N100)? data_i[2537] : 
                       (N102)? data_i[2665] : 
                       (N104)? data_i[2793] : 
                       (N106)? data_i[2921] : 
                       (N108)? data_i[3049] : 
                       (N110)? data_i[3177] : 
                       (N112)? data_i[3305] : 
                       (N114)? data_i[3433] : 
                       (N116)? data_i[3561] : 
                       (N118)? data_i[3689] : 
                       (N120)? data_i[3817] : 
                       (N122)? data_i[3945] : 
                       (N124)? data_i[4073] : 1'b0;
  assign data_o[104] = (N93)? data_i[104] : 
                       (N95)? data_i[232] : 
                       (N97)? data_i[360] : 
                       (N99)? data_i[488] : 
                       (N101)? data_i[616] : 
                       (N103)? data_i[744] : 
                       (N105)? data_i[872] : 
                       (N107)? data_i[1000] : 
                       (N109)? data_i[1128] : 
                       (N111)? data_i[1256] : 
                       (N113)? data_i[1384] : 
                       (N115)? data_i[1512] : 
                       (N117)? data_i[1640] : 
                       (N119)? data_i[1768] : 
                       (N121)? data_i[1896] : 
                       (N123)? data_i[2024] : 
                       (N94)? data_i[2152] : 
                       (N96)? data_i[2280] : 
                       (N98)? data_i[2408] : 
                       (N100)? data_i[2536] : 
                       (N102)? data_i[2664] : 
                       (N104)? data_i[2792] : 
                       (N106)? data_i[2920] : 
                       (N108)? data_i[3048] : 
                       (N110)? data_i[3176] : 
                       (N112)? data_i[3304] : 
                       (N114)? data_i[3432] : 
                       (N116)? data_i[3560] : 
                       (N118)? data_i[3688] : 
                       (N120)? data_i[3816] : 
                       (N122)? data_i[3944] : 
                       (N124)? data_i[4072] : 1'b0;
  assign data_o[103] = (N93)? data_i[103] : 
                       (N95)? data_i[231] : 
                       (N97)? data_i[359] : 
                       (N99)? data_i[487] : 
                       (N101)? data_i[615] : 
                       (N103)? data_i[743] : 
                       (N105)? data_i[871] : 
                       (N107)? data_i[999] : 
                       (N109)? data_i[1127] : 
                       (N111)? data_i[1255] : 
                       (N113)? data_i[1383] : 
                       (N115)? data_i[1511] : 
                       (N117)? data_i[1639] : 
                       (N119)? data_i[1767] : 
                       (N121)? data_i[1895] : 
                       (N123)? data_i[2023] : 
                       (N94)? data_i[2151] : 
                       (N96)? data_i[2279] : 
                       (N98)? data_i[2407] : 
                       (N100)? data_i[2535] : 
                       (N102)? data_i[2663] : 
                       (N104)? data_i[2791] : 
                       (N106)? data_i[2919] : 
                       (N108)? data_i[3047] : 
                       (N110)? data_i[3175] : 
                       (N112)? data_i[3303] : 
                       (N114)? data_i[3431] : 
                       (N116)? data_i[3559] : 
                       (N118)? data_i[3687] : 
                       (N120)? data_i[3815] : 
                       (N122)? data_i[3943] : 
                       (N124)? data_i[4071] : 1'b0;
  assign data_o[102] = (N93)? data_i[102] : 
                       (N95)? data_i[230] : 
                       (N97)? data_i[358] : 
                       (N99)? data_i[486] : 
                       (N101)? data_i[614] : 
                       (N103)? data_i[742] : 
                       (N105)? data_i[870] : 
                       (N107)? data_i[998] : 
                       (N109)? data_i[1126] : 
                       (N111)? data_i[1254] : 
                       (N113)? data_i[1382] : 
                       (N115)? data_i[1510] : 
                       (N117)? data_i[1638] : 
                       (N119)? data_i[1766] : 
                       (N121)? data_i[1894] : 
                       (N123)? data_i[2022] : 
                       (N94)? data_i[2150] : 
                       (N96)? data_i[2278] : 
                       (N98)? data_i[2406] : 
                       (N100)? data_i[2534] : 
                       (N102)? data_i[2662] : 
                       (N104)? data_i[2790] : 
                       (N106)? data_i[2918] : 
                       (N108)? data_i[3046] : 
                       (N110)? data_i[3174] : 
                       (N112)? data_i[3302] : 
                       (N114)? data_i[3430] : 
                       (N116)? data_i[3558] : 
                       (N118)? data_i[3686] : 
                       (N120)? data_i[3814] : 
                       (N122)? data_i[3942] : 
                       (N124)? data_i[4070] : 1'b0;
  assign data_o[101] = (N93)? data_i[101] : 
                       (N95)? data_i[229] : 
                       (N97)? data_i[357] : 
                       (N99)? data_i[485] : 
                       (N101)? data_i[613] : 
                       (N103)? data_i[741] : 
                       (N105)? data_i[869] : 
                       (N107)? data_i[997] : 
                       (N109)? data_i[1125] : 
                       (N111)? data_i[1253] : 
                       (N113)? data_i[1381] : 
                       (N115)? data_i[1509] : 
                       (N117)? data_i[1637] : 
                       (N119)? data_i[1765] : 
                       (N121)? data_i[1893] : 
                       (N123)? data_i[2021] : 
                       (N94)? data_i[2149] : 
                       (N96)? data_i[2277] : 
                       (N98)? data_i[2405] : 
                       (N100)? data_i[2533] : 
                       (N102)? data_i[2661] : 
                       (N104)? data_i[2789] : 
                       (N106)? data_i[2917] : 
                       (N108)? data_i[3045] : 
                       (N110)? data_i[3173] : 
                       (N112)? data_i[3301] : 
                       (N114)? data_i[3429] : 
                       (N116)? data_i[3557] : 
                       (N118)? data_i[3685] : 
                       (N120)? data_i[3813] : 
                       (N122)? data_i[3941] : 
                       (N124)? data_i[4069] : 1'b0;
  assign data_o[100] = (N93)? data_i[100] : 
                       (N95)? data_i[228] : 
                       (N97)? data_i[356] : 
                       (N99)? data_i[484] : 
                       (N101)? data_i[612] : 
                       (N103)? data_i[740] : 
                       (N105)? data_i[868] : 
                       (N107)? data_i[996] : 
                       (N109)? data_i[1124] : 
                       (N111)? data_i[1252] : 
                       (N113)? data_i[1380] : 
                       (N115)? data_i[1508] : 
                       (N117)? data_i[1636] : 
                       (N119)? data_i[1764] : 
                       (N121)? data_i[1892] : 
                       (N123)? data_i[2020] : 
                       (N94)? data_i[2148] : 
                       (N96)? data_i[2276] : 
                       (N98)? data_i[2404] : 
                       (N100)? data_i[2532] : 
                       (N102)? data_i[2660] : 
                       (N104)? data_i[2788] : 
                       (N106)? data_i[2916] : 
                       (N108)? data_i[3044] : 
                       (N110)? data_i[3172] : 
                       (N112)? data_i[3300] : 
                       (N114)? data_i[3428] : 
                       (N116)? data_i[3556] : 
                       (N118)? data_i[3684] : 
                       (N120)? data_i[3812] : 
                       (N122)? data_i[3940] : 
                       (N124)? data_i[4068] : 1'b0;
  assign data_o[99] = (N93)? data_i[99] : 
                      (N95)? data_i[227] : 
                      (N97)? data_i[355] : 
                      (N99)? data_i[483] : 
                      (N101)? data_i[611] : 
                      (N103)? data_i[739] : 
                      (N105)? data_i[867] : 
                      (N107)? data_i[995] : 
                      (N109)? data_i[1123] : 
                      (N111)? data_i[1251] : 
                      (N113)? data_i[1379] : 
                      (N115)? data_i[1507] : 
                      (N117)? data_i[1635] : 
                      (N119)? data_i[1763] : 
                      (N121)? data_i[1891] : 
                      (N123)? data_i[2019] : 
                      (N94)? data_i[2147] : 
                      (N96)? data_i[2275] : 
                      (N98)? data_i[2403] : 
                      (N100)? data_i[2531] : 
                      (N102)? data_i[2659] : 
                      (N104)? data_i[2787] : 
                      (N106)? data_i[2915] : 
                      (N108)? data_i[3043] : 
                      (N110)? data_i[3171] : 
                      (N112)? data_i[3299] : 
                      (N114)? data_i[3427] : 
                      (N116)? data_i[3555] : 
                      (N118)? data_i[3683] : 
                      (N120)? data_i[3811] : 
                      (N122)? data_i[3939] : 
                      (N124)? data_i[4067] : 1'b0;
  assign data_o[98] = (N93)? data_i[98] : 
                      (N95)? data_i[226] : 
                      (N97)? data_i[354] : 
                      (N99)? data_i[482] : 
                      (N101)? data_i[610] : 
                      (N103)? data_i[738] : 
                      (N105)? data_i[866] : 
                      (N107)? data_i[994] : 
                      (N109)? data_i[1122] : 
                      (N111)? data_i[1250] : 
                      (N113)? data_i[1378] : 
                      (N115)? data_i[1506] : 
                      (N117)? data_i[1634] : 
                      (N119)? data_i[1762] : 
                      (N121)? data_i[1890] : 
                      (N123)? data_i[2018] : 
                      (N94)? data_i[2146] : 
                      (N96)? data_i[2274] : 
                      (N98)? data_i[2402] : 
                      (N100)? data_i[2530] : 
                      (N102)? data_i[2658] : 
                      (N104)? data_i[2786] : 
                      (N106)? data_i[2914] : 
                      (N108)? data_i[3042] : 
                      (N110)? data_i[3170] : 
                      (N112)? data_i[3298] : 
                      (N114)? data_i[3426] : 
                      (N116)? data_i[3554] : 
                      (N118)? data_i[3682] : 
                      (N120)? data_i[3810] : 
                      (N122)? data_i[3938] : 
                      (N124)? data_i[4066] : 1'b0;
  assign data_o[97] = (N93)? data_i[97] : 
                      (N95)? data_i[225] : 
                      (N97)? data_i[353] : 
                      (N99)? data_i[481] : 
                      (N101)? data_i[609] : 
                      (N103)? data_i[737] : 
                      (N105)? data_i[865] : 
                      (N107)? data_i[993] : 
                      (N109)? data_i[1121] : 
                      (N111)? data_i[1249] : 
                      (N113)? data_i[1377] : 
                      (N115)? data_i[1505] : 
                      (N117)? data_i[1633] : 
                      (N119)? data_i[1761] : 
                      (N121)? data_i[1889] : 
                      (N123)? data_i[2017] : 
                      (N94)? data_i[2145] : 
                      (N96)? data_i[2273] : 
                      (N98)? data_i[2401] : 
                      (N100)? data_i[2529] : 
                      (N102)? data_i[2657] : 
                      (N104)? data_i[2785] : 
                      (N106)? data_i[2913] : 
                      (N108)? data_i[3041] : 
                      (N110)? data_i[3169] : 
                      (N112)? data_i[3297] : 
                      (N114)? data_i[3425] : 
                      (N116)? data_i[3553] : 
                      (N118)? data_i[3681] : 
                      (N120)? data_i[3809] : 
                      (N122)? data_i[3937] : 
                      (N124)? data_i[4065] : 1'b0;
  assign data_o[96] = (N93)? data_i[96] : 
                      (N95)? data_i[224] : 
                      (N97)? data_i[352] : 
                      (N99)? data_i[480] : 
                      (N101)? data_i[608] : 
                      (N103)? data_i[736] : 
                      (N105)? data_i[864] : 
                      (N107)? data_i[992] : 
                      (N109)? data_i[1120] : 
                      (N111)? data_i[1248] : 
                      (N113)? data_i[1376] : 
                      (N115)? data_i[1504] : 
                      (N117)? data_i[1632] : 
                      (N119)? data_i[1760] : 
                      (N121)? data_i[1888] : 
                      (N123)? data_i[2016] : 
                      (N94)? data_i[2144] : 
                      (N96)? data_i[2272] : 
                      (N98)? data_i[2400] : 
                      (N100)? data_i[2528] : 
                      (N102)? data_i[2656] : 
                      (N104)? data_i[2784] : 
                      (N106)? data_i[2912] : 
                      (N108)? data_i[3040] : 
                      (N110)? data_i[3168] : 
                      (N112)? data_i[3296] : 
                      (N114)? data_i[3424] : 
                      (N116)? data_i[3552] : 
                      (N118)? data_i[3680] : 
                      (N120)? data_i[3808] : 
                      (N122)? data_i[3936] : 
                      (N124)? data_i[4064] : 1'b0;
  assign data_o[95] = (N93)? data_i[95] : 
                      (N95)? data_i[223] : 
                      (N97)? data_i[351] : 
                      (N99)? data_i[479] : 
                      (N101)? data_i[607] : 
                      (N103)? data_i[735] : 
                      (N105)? data_i[863] : 
                      (N107)? data_i[991] : 
                      (N109)? data_i[1119] : 
                      (N111)? data_i[1247] : 
                      (N113)? data_i[1375] : 
                      (N115)? data_i[1503] : 
                      (N117)? data_i[1631] : 
                      (N119)? data_i[1759] : 
                      (N121)? data_i[1887] : 
                      (N123)? data_i[2015] : 
                      (N94)? data_i[2143] : 
                      (N96)? data_i[2271] : 
                      (N98)? data_i[2399] : 
                      (N100)? data_i[2527] : 
                      (N102)? data_i[2655] : 
                      (N104)? data_i[2783] : 
                      (N106)? data_i[2911] : 
                      (N108)? data_i[3039] : 
                      (N110)? data_i[3167] : 
                      (N112)? data_i[3295] : 
                      (N114)? data_i[3423] : 
                      (N116)? data_i[3551] : 
                      (N118)? data_i[3679] : 
                      (N120)? data_i[3807] : 
                      (N122)? data_i[3935] : 
                      (N124)? data_i[4063] : 1'b0;
  assign data_o[94] = (N93)? data_i[94] : 
                      (N95)? data_i[222] : 
                      (N97)? data_i[350] : 
                      (N99)? data_i[478] : 
                      (N101)? data_i[606] : 
                      (N103)? data_i[734] : 
                      (N105)? data_i[862] : 
                      (N107)? data_i[990] : 
                      (N109)? data_i[1118] : 
                      (N111)? data_i[1246] : 
                      (N113)? data_i[1374] : 
                      (N115)? data_i[1502] : 
                      (N117)? data_i[1630] : 
                      (N119)? data_i[1758] : 
                      (N121)? data_i[1886] : 
                      (N123)? data_i[2014] : 
                      (N94)? data_i[2142] : 
                      (N96)? data_i[2270] : 
                      (N98)? data_i[2398] : 
                      (N100)? data_i[2526] : 
                      (N102)? data_i[2654] : 
                      (N104)? data_i[2782] : 
                      (N106)? data_i[2910] : 
                      (N108)? data_i[3038] : 
                      (N110)? data_i[3166] : 
                      (N112)? data_i[3294] : 
                      (N114)? data_i[3422] : 
                      (N116)? data_i[3550] : 
                      (N118)? data_i[3678] : 
                      (N120)? data_i[3806] : 
                      (N122)? data_i[3934] : 
                      (N124)? data_i[4062] : 1'b0;
  assign data_o[93] = (N93)? data_i[93] : 
                      (N95)? data_i[221] : 
                      (N97)? data_i[349] : 
                      (N99)? data_i[477] : 
                      (N101)? data_i[605] : 
                      (N103)? data_i[733] : 
                      (N105)? data_i[861] : 
                      (N107)? data_i[989] : 
                      (N109)? data_i[1117] : 
                      (N111)? data_i[1245] : 
                      (N113)? data_i[1373] : 
                      (N115)? data_i[1501] : 
                      (N117)? data_i[1629] : 
                      (N119)? data_i[1757] : 
                      (N121)? data_i[1885] : 
                      (N123)? data_i[2013] : 
                      (N94)? data_i[2141] : 
                      (N96)? data_i[2269] : 
                      (N98)? data_i[2397] : 
                      (N100)? data_i[2525] : 
                      (N102)? data_i[2653] : 
                      (N104)? data_i[2781] : 
                      (N106)? data_i[2909] : 
                      (N108)? data_i[3037] : 
                      (N110)? data_i[3165] : 
                      (N112)? data_i[3293] : 
                      (N114)? data_i[3421] : 
                      (N116)? data_i[3549] : 
                      (N118)? data_i[3677] : 
                      (N120)? data_i[3805] : 
                      (N122)? data_i[3933] : 
                      (N124)? data_i[4061] : 1'b0;
  assign data_o[92] = (N93)? data_i[92] : 
                      (N95)? data_i[220] : 
                      (N97)? data_i[348] : 
                      (N99)? data_i[476] : 
                      (N101)? data_i[604] : 
                      (N103)? data_i[732] : 
                      (N105)? data_i[860] : 
                      (N107)? data_i[988] : 
                      (N109)? data_i[1116] : 
                      (N111)? data_i[1244] : 
                      (N113)? data_i[1372] : 
                      (N115)? data_i[1500] : 
                      (N117)? data_i[1628] : 
                      (N119)? data_i[1756] : 
                      (N121)? data_i[1884] : 
                      (N123)? data_i[2012] : 
                      (N94)? data_i[2140] : 
                      (N96)? data_i[2268] : 
                      (N98)? data_i[2396] : 
                      (N100)? data_i[2524] : 
                      (N102)? data_i[2652] : 
                      (N104)? data_i[2780] : 
                      (N106)? data_i[2908] : 
                      (N108)? data_i[3036] : 
                      (N110)? data_i[3164] : 
                      (N112)? data_i[3292] : 
                      (N114)? data_i[3420] : 
                      (N116)? data_i[3548] : 
                      (N118)? data_i[3676] : 
                      (N120)? data_i[3804] : 
                      (N122)? data_i[3932] : 
                      (N124)? data_i[4060] : 1'b0;
  assign data_o[91] = (N93)? data_i[91] : 
                      (N95)? data_i[219] : 
                      (N97)? data_i[347] : 
                      (N99)? data_i[475] : 
                      (N101)? data_i[603] : 
                      (N103)? data_i[731] : 
                      (N105)? data_i[859] : 
                      (N107)? data_i[987] : 
                      (N109)? data_i[1115] : 
                      (N111)? data_i[1243] : 
                      (N113)? data_i[1371] : 
                      (N115)? data_i[1499] : 
                      (N117)? data_i[1627] : 
                      (N119)? data_i[1755] : 
                      (N121)? data_i[1883] : 
                      (N123)? data_i[2011] : 
                      (N94)? data_i[2139] : 
                      (N96)? data_i[2267] : 
                      (N98)? data_i[2395] : 
                      (N100)? data_i[2523] : 
                      (N102)? data_i[2651] : 
                      (N104)? data_i[2779] : 
                      (N106)? data_i[2907] : 
                      (N108)? data_i[3035] : 
                      (N110)? data_i[3163] : 
                      (N112)? data_i[3291] : 
                      (N114)? data_i[3419] : 
                      (N116)? data_i[3547] : 
                      (N118)? data_i[3675] : 
                      (N120)? data_i[3803] : 
                      (N122)? data_i[3931] : 
                      (N124)? data_i[4059] : 1'b0;
  assign data_o[90] = (N93)? data_i[90] : 
                      (N95)? data_i[218] : 
                      (N97)? data_i[346] : 
                      (N99)? data_i[474] : 
                      (N101)? data_i[602] : 
                      (N103)? data_i[730] : 
                      (N105)? data_i[858] : 
                      (N107)? data_i[986] : 
                      (N109)? data_i[1114] : 
                      (N111)? data_i[1242] : 
                      (N113)? data_i[1370] : 
                      (N115)? data_i[1498] : 
                      (N117)? data_i[1626] : 
                      (N119)? data_i[1754] : 
                      (N121)? data_i[1882] : 
                      (N123)? data_i[2010] : 
                      (N94)? data_i[2138] : 
                      (N96)? data_i[2266] : 
                      (N98)? data_i[2394] : 
                      (N100)? data_i[2522] : 
                      (N102)? data_i[2650] : 
                      (N104)? data_i[2778] : 
                      (N106)? data_i[2906] : 
                      (N108)? data_i[3034] : 
                      (N110)? data_i[3162] : 
                      (N112)? data_i[3290] : 
                      (N114)? data_i[3418] : 
                      (N116)? data_i[3546] : 
                      (N118)? data_i[3674] : 
                      (N120)? data_i[3802] : 
                      (N122)? data_i[3930] : 
                      (N124)? data_i[4058] : 1'b0;
  assign data_o[89] = (N93)? data_i[89] : 
                      (N95)? data_i[217] : 
                      (N97)? data_i[345] : 
                      (N99)? data_i[473] : 
                      (N101)? data_i[601] : 
                      (N103)? data_i[729] : 
                      (N105)? data_i[857] : 
                      (N107)? data_i[985] : 
                      (N109)? data_i[1113] : 
                      (N111)? data_i[1241] : 
                      (N113)? data_i[1369] : 
                      (N115)? data_i[1497] : 
                      (N117)? data_i[1625] : 
                      (N119)? data_i[1753] : 
                      (N121)? data_i[1881] : 
                      (N123)? data_i[2009] : 
                      (N94)? data_i[2137] : 
                      (N96)? data_i[2265] : 
                      (N98)? data_i[2393] : 
                      (N100)? data_i[2521] : 
                      (N102)? data_i[2649] : 
                      (N104)? data_i[2777] : 
                      (N106)? data_i[2905] : 
                      (N108)? data_i[3033] : 
                      (N110)? data_i[3161] : 
                      (N112)? data_i[3289] : 
                      (N114)? data_i[3417] : 
                      (N116)? data_i[3545] : 
                      (N118)? data_i[3673] : 
                      (N120)? data_i[3801] : 
                      (N122)? data_i[3929] : 
                      (N124)? data_i[4057] : 1'b0;
  assign data_o[88] = (N93)? data_i[88] : 
                      (N95)? data_i[216] : 
                      (N97)? data_i[344] : 
                      (N99)? data_i[472] : 
                      (N101)? data_i[600] : 
                      (N103)? data_i[728] : 
                      (N105)? data_i[856] : 
                      (N107)? data_i[984] : 
                      (N109)? data_i[1112] : 
                      (N111)? data_i[1240] : 
                      (N113)? data_i[1368] : 
                      (N115)? data_i[1496] : 
                      (N117)? data_i[1624] : 
                      (N119)? data_i[1752] : 
                      (N121)? data_i[1880] : 
                      (N123)? data_i[2008] : 
                      (N94)? data_i[2136] : 
                      (N96)? data_i[2264] : 
                      (N98)? data_i[2392] : 
                      (N100)? data_i[2520] : 
                      (N102)? data_i[2648] : 
                      (N104)? data_i[2776] : 
                      (N106)? data_i[2904] : 
                      (N108)? data_i[3032] : 
                      (N110)? data_i[3160] : 
                      (N112)? data_i[3288] : 
                      (N114)? data_i[3416] : 
                      (N116)? data_i[3544] : 
                      (N118)? data_i[3672] : 
                      (N120)? data_i[3800] : 
                      (N122)? data_i[3928] : 
                      (N124)? data_i[4056] : 1'b0;
  assign data_o[87] = (N93)? data_i[87] : 
                      (N95)? data_i[215] : 
                      (N97)? data_i[343] : 
                      (N99)? data_i[471] : 
                      (N101)? data_i[599] : 
                      (N103)? data_i[727] : 
                      (N105)? data_i[855] : 
                      (N107)? data_i[983] : 
                      (N109)? data_i[1111] : 
                      (N111)? data_i[1239] : 
                      (N113)? data_i[1367] : 
                      (N115)? data_i[1495] : 
                      (N117)? data_i[1623] : 
                      (N119)? data_i[1751] : 
                      (N121)? data_i[1879] : 
                      (N123)? data_i[2007] : 
                      (N94)? data_i[2135] : 
                      (N96)? data_i[2263] : 
                      (N98)? data_i[2391] : 
                      (N100)? data_i[2519] : 
                      (N102)? data_i[2647] : 
                      (N104)? data_i[2775] : 
                      (N106)? data_i[2903] : 
                      (N108)? data_i[3031] : 
                      (N110)? data_i[3159] : 
                      (N112)? data_i[3287] : 
                      (N114)? data_i[3415] : 
                      (N116)? data_i[3543] : 
                      (N118)? data_i[3671] : 
                      (N120)? data_i[3799] : 
                      (N122)? data_i[3927] : 
                      (N124)? data_i[4055] : 1'b0;
  assign data_o[86] = (N93)? data_i[86] : 
                      (N95)? data_i[214] : 
                      (N97)? data_i[342] : 
                      (N99)? data_i[470] : 
                      (N101)? data_i[598] : 
                      (N103)? data_i[726] : 
                      (N105)? data_i[854] : 
                      (N107)? data_i[982] : 
                      (N109)? data_i[1110] : 
                      (N111)? data_i[1238] : 
                      (N113)? data_i[1366] : 
                      (N115)? data_i[1494] : 
                      (N117)? data_i[1622] : 
                      (N119)? data_i[1750] : 
                      (N121)? data_i[1878] : 
                      (N123)? data_i[2006] : 
                      (N94)? data_i[2134] : 
                      (N96)? data_i[2262] : 
                      (N98)? data_i[2390] : 
                      (N100)? data_i[2518] : 
                      (N102)? data_i[2646] : 
                      (N104)? data_i[2774] : 
                      (N106)? data_i[2902] : 
                      (N108)? data_i[3030] : 
                      (N110)? data_i[3158] : 
                      (N112)? data_i[3286] : 
                      (N114)? data_i[3414] : 
                      (N116)? data_i[3542] : 
                      (N118)? data_i[3670] : 
                      (N120)? data_i[3798] : 
                      (N122)? data_i[3926] : 
                      (N124)? data_i[4054] : 1'b0;
  assign data_o[85] = (N93)? data_i[85] : 
                      (N95)? data_i[213] : 
                      (N97)? data_i[341] : 
                      (N99)? data_i[469] : 
                      (N101)? data_i[597] : 
                      (N103)? data_i[725] : 
                      (N105)? data_i[853] : 
                      (N107)? data_i[981] : 
                      (N109)? data_i[1109] : 
                      (N111)? data_i[1237] : 
                      (N113)? data_i[1365] : 
                      (N115)? data_i[1493] : 
                      (N117)? data_i[1621] : 
                      (N119)? data_i[1749] : 
                      (N121)? data_i[1877] : 
                      (N123)? data_i[2005] : 
                      (N94)? data_i[2133] : 
                      (N96)? data_i[2261] : 
                      (N98)? data_i[2389] : 
                      (N100)? data_i[2517] : 
                      (N102)? data_i[2645] : 
                      (N104)? data_i[2773] : 
                      (N106)? data_i[2901] : 
                      (N108)? data_i[3029] : 
                      (N110)? data_i[3157] : 
                      (N112)? data_i[3285] : 
                      (N114)? data_i[3413] : 
                      (N116)? data_i[3541] : 
                      (N118)? data_i[3669] : 
                      (N120)? data_i[3797] : 
                      (N122)? data_i[3925] : 
                      (N124)? data_i[4053] : 1'b0;
  assign data_o[84] = (N93)? data_i[84] : 
                      (N95)? data_i[212] : 
                      (N97)? data_i[340] : 
                      (N99)? data_i[468] : 
                      (N101)? data_i[596] : 
                      (N103)? data_i[724] : 
                      (N105)? data_i[852] : 
                      (N107)? data_i[980] : 
                      (N109)? data_i[1108] : 
                      (N111)? data_i[1236] : 
                      (N113)? data_i[1364] : 
                      (N115)? data_i[1492] : 
                      (N117)? data_i[1620] : 
                      (N119)? data_i[1748] : 
                      (N121)? data_i[1876] : 
                      (N123)? data_i[2004] : 
                      (N94)? data_i[2132] : 
                      (N96)? data_i[2260] : 
                      (N98)? data_i[2388] : 
                      (N100)? data_i[2516] : 
                      (N102)? data_i[2644] : 
                      (N104)? data_i[2772] : 
                      (N106)? data_i[2900] : 
                      (N108)? data_i[3028] : 
                      (N110)? data_i[3156] : 
                      (N112)? data_i[3284] : 
                      (N114)? data_i[3412] : 
                      (N116)? data_i[3540] : 
                      (N118)? data_i[3668] : 
                      (N120)? data_i[3796] : 
                      (N122)? data_i[3924] : 
                      (N124)? data_i[4052] : 1'b0;
  assign data_o[83] = (N93)? data_i[83] : 
                      (N95)? data_i[211] : 
                      (N97)? data_i[339] : 
                      (N99)? data_i[467] : 
                      (N101)? data_i[595] : 
                      (N103)? data_i[723] : 
                      (N105)? data_i[851] : 
                      (N107)? data_i[979] : 
                      (N109)? data_i[1107] : 
                      (N111)? data_i[1235] : 
                      (N113)? data_i[1363] : 
                      (N115)? data_i[1491] : 
                      (N117)? data_i[1619] : 
                      (N119)? data_i[1747] : 
                      (N121)? data_i[1875] : 
                      (N123)? data_i[2003] : 
                      (N94)? data_i[2131] : 
                      (N96)? data_i[2259] : 
                      (N98)? data_i[2387] : 
                      (N100)? data_i[2515] : 
                      (N102)? data_i[2643] : 
                      (N104)? data_i[2771] : 
                      (N106)? data_i[2899] : 
                      (N108)? data_i[3027] : 
                      (N110)? data_i[3155] : 
                      (N112)? data_i[3283] : 
                      (N114)? data_i[3411] : 
                      (N116)? data_i[3539] : 
                      (N118)? data_i[3667] : 
                      (N120)? data_i[3795] : 
                      (N122)? data_i[3923] : 
                      (N124)? data_i[4051] : 1'b0;
  assign data_o[82] = (N93)? data_i[82] : 
                      (N95)? data_i[210] : 
                      (N97)? data_i[338] : 
                      (N99)? data_i[466] : 
                      (N101)? data_i[594] : 
                      (N103)? data_i[722] : 
                      (N105)? data_i[850] : 
                      (N107)? data_i[978] : 
                      (N109)? data_i[1106] : 
                      (N111)? data_i[1234] : 
                      (N113)? data_i[1362] : 
                      (N115)? data_i[1490] : 
                      (N117)? data_i[1618] : 
                      (N119)? data_i[1746] : 
                      (N121)? data_i[1874] : 
                      (N123)? data_i[2002] : 
                      (N94)? data_i[2130] : 
                      (N96)? data_i[2258] : 
                      (N98)? data_i[2386] : 
                      (N100)? data_i[2514] : 
                      (N102)? data_i[2642] : 
                      (N104)? data_i[2770] : 
                      (N106)? data_i[2898] : 
                      (N108)? data_i[3026] : 
                      (N110)? data_i[3154] : 
                      (N112)? data_i[3282] : 
                      (N114)? data_i[3410] : 
                      (N116)? data_i[3538] : 
                      (N118)? data_i[3666] : 
                      (N120)? data_i[3794] : 
                      (N122)? data_i[3922] : 
                      (N124)? data_i[4050] : 1'b0;
  assign data_o[81] = (N93)? data_i[81] : 
                      (N95)? data_i[209] : 
                      (N97)? data_i[337] : 
                      (N99)? data_i[465] : 
                      (N101)? data_i[593] : 
                      (N103)? data_i[721] : 
                      (N105)? data_i[849] : 
                      (N107)? data_i[977] : 
                      (N109)? data_i[1105] : 
                      (N111)? data_i[1233] : 
                      (N113)? data_i[1361] : 
                      (N115)? data_i[1489] : 
                      (N117)? data_i[1617] : 
                      (N119)? data_i[1745] : 
                      (N121)? data_i[1873] : 
                      (N123)? data_i[2001] : 
                      (N94)? data_i[2129] : 
                      (N96)? data_i[2257] : 
                      (N98)? data_i[2385] : 
                      (N100)? data_i[2513] : 
                      (N102)? data_i[2641] : 
                      (N104)? data_i[2769] : 
                      (N106)? data_i[2897] : 
                      (N108)? data_i[3025] : 
                      (N110)? data_i[3153] : 
                      (N112)? data_i[3281] : 
                      (N114)? data_i[3409] : 
                      (N116)? data_i[3537] : 
                      (N118)? data_i[3665] : 
                      (N120)? data_i[3793] : 
                      (N122)? data_i[3921] : 
                      (N124)? data_i[4049] : 1'b0;
  assign data_o[80] = (N93)? data_i[80] : 
                      (N95)? data_i[208] : 
                      (N97)? data_i[336] : 
                      (N99)? data_i[464] : 
                      (N101)? data_i[592] : 
                      (N103)? data_i[720] : 
                      (N105)? data_i[848] : 
                      (N107)? data_i[976] : 
                      (N109)? data_i[1104] : 
                      (N111)? data_i[1232] : 
                      (N113)? data_i[1360] : 
                      (N115)? data_i[1488] : 
                      (N117)? data_i[1616] : 
                      (N119)? data_i[1744] : 
                      (N121)? data_i[1872] : 
                      (N123)? data_i[2000] : 
                      (N94)? data_i[2128] : 
                      (N96)? data_i[2256] : 
                      (N98)? data_i[2384] : 
                      (N100)? data_i[2512] : 
                      (N102)? data_i[2640] : 
                      (N104)? data_i[2768] : 
                      (N106)? data_i[2896] : 
                      (N108)? data_i[3024] : 
                      (N110)? data_i[3152] : 
                      (N112)? data_i[3280] : 
                      (N114)? data_i[3408] : 
                      (N116)? data_i[3536] : 
                      (N118)? data_i[3664] : 
                      (N120)? data_i[3792] : 
                      (N122)? data_i[3920] : 
                      (N124)? data_i[4048] : 1'b0;
  assign data_o[79] = (N93)? data_i[79] : 
                      (N95)? data_i[207] : 
                      (N97)? data_i[335] : 
                      (N99)? data_i[463] : 
                      (N101)? data_i[591] : 
                      (N103)? data_i[719] : 
                      (N105)? data_i[847] : 
                      (N107)? data_i[975] : 
                      (N109)? data_i[1103] : 
                      (N111)? data_i[1231] : 
                      (N113)? data_i[1359] : 
                      (N115)? data_i[1487] : 
                      (N117)? data_i[1615] : 
                      (N119)? data_i[1743] : 
                      (N121)? data_i[1871] : 
                      (N123)? data_i[1999] : 
                      (N94)? data_i[2127] : 
                      (N96)? data_i[2255] : 
                      (N98)? data_i[2383] : 
                      (N100)? data_i[2511] : 
                      (N102)? data_i[2639] : 
                      (N104)? data_i[2767] : 
                      (N106)? data_i[2895] : 
                      (N108)? data_i[3023] : 
                      (N110)? data_i[3151] : 
                      (N112)? data_i[3279] : 
                      (N114)? data_i[3407] : 
                      (N116)? data_i[3535] : 
                      (N118)? data_i[3663] : 
                      (N120)? data_i[3791] : 
                      (N122)? data_i[3919] : 
                      (N124)? data_i[4047] : 1'b0;
  assign data_o[78] = (N93)? data_i[78] : 
                      (N95)? data_i[206] : 
                      (N97)? data_i[334] : 
                      (N99)? data_i[462] : 
                      (N101)? data_i[590] : 
                      (N103)? data_i[718] : 
                      (N105)? data_i[846] : 
                      (N107)? data_i[974] : 
                      (N109)? data_i[1102] : 
                      (N111)? data_i[1230] : 
                      (N113)? data_i[1358] : 
                      (N115)? data_i[1486] : 
                      (N117)? data_i[1614] : 
                      (N119)? data_i[1742] : 
                      (N121)? data_i[1870] : 
                      (N123)? data_i[1998] : 
                      (N94)? data_i[2126] : 
                      (N96)? data_i[2254] : 
                      (N98)? data_i[2382] : 
                      (N100)? data_i[2510] : 
                      (N102)? data_i[2638] : 
                      (N104)? data_i[2766] : 
                      (N106)? data_i[2894] : 
                      (N108)? data_i[3022] : 
                      (N110)? data_i[3150] : 
                      (N112)? data_i[3278] : 
                      (N114)? data_i[3406] : 
                      (N116)? data_i[3534] : 
                      (N118)? data_i[3662] : 
                      (N120)? data_i[3790] : 
                      (N122)? data_i[3918] : 
                      (N124)? data_i[4046] : 1'b0;
  assign data_o[77] = (N93)? data_i[77] : 
                      (N95)? data_i[205] : 
                      (N97)? data_i[333] : 
                      (N99)? data_i[461] : 
                      (N101)? data_i[589] : 
                      (N103)? data_i[717] : 
                      (N105)? data_i[845] : 
                      (N107)? data_i[973] : 
                      (N109)? data_i[1101] : 
                      (N111)? data_i[1229] : 
                      (N113)? data_i[1357] : 
                      (N115)? data_i[1485] : 
                      (N117)? data_i[1613] : 
                      (N119)? data_i[1741] : 
                      (N121)? data_i[1869] : 
                      (N123)? data_i[1997] : 
                      (N94)? data_i[2125] : 
                      (N96)? data_i[2253] : 
                      (N98)? data_i[2381] : 
                      (N100)? data_i[2509] : 
                      (N102)? data_i[2637] : 
                      (N104)? data_i[2765] : 
                      (N106)? data_i[2893] : 
                      (N108)? data_i[3021] : 
                      (N110)? data_i[3149] : 
                      (N112)? data_i[3277] : 
                      (N114)? data_i[3405] : 
                      (N116)? data_i[3533] : 
                      (N118)? data_i[3661] : 
                      (N120)? data_i[3789] : 
                      (N122)? data_i[3917] : 
                      (N124)? data_i[4045] : 1'b0;
  assign data_o[76] = (N93)? data_i[76] : 
                      (N95)? data_i[204] : 
                      (N97)? data_i[332] : 
                      (N99)? data_i[460] : 
                      (N101)? data_i[588] : 
                      (N103)? data_i[716] : 
                      (N105)? data_i[844] : 
                      (N107)? data_i[972] : 
                      (N109)? data_i[1100] : 
                      (N111)? data_i[1228] : 
                      (N113)? data_i[1356] : 
                      (N115)? data_i[1484] : 
                      (N117)? data_i[1612] : 
                      (N119)? data_i[1740] : 
                      (N121)? data_i[1868] : 
                      (N123)? data_i[1996] : 
                      (N94)? data_i[2124] : 
                      (N96)? data_i[2252] : 
                      (N98)? data_i[2380] : 
                      (N100)? data_i[2508] : 
                      (N102)? data_i[2636] : 
                      (N104)? data_i[2764] : 
                      (N106)? data_i[2892] : 
                      (N108)? data_i[3020] : 
                      (N110)? data_i[3148] : 
                      (N112)? data_i[3276] : 
                      (N114)? data_i[3404] : 
                      (N116)? data_i[3532] : 
                      (N118)? data_i[3660] : 
                      (N120)? data_i[3788] : 
                      (N122)? data_i[3916] : 
                      (N124)? data_i[4044] : 1'b0;
  assign data_o[75] = (N93)? data_i[75] : 
                      (N95)? data_i[203] : 
                      (N97)? data_i[331] : 
                      (N99)? data_i[459] : 
                      (N101)? data_i[587] : 
                      (N103)? data_i[715] : 
                      (N105)? data_i[843] : 
                      (N107)? data_i[971] : 
                      (N109)? data_i[1099] : 
                      (N111)? data_i[1227] : 
                      (N113)? data_i[1355] : 
                      (N115)? data_i[1483] : 
                      (N117)? data_i[1611] : 
                      (N119)? data_i[1739] : 
                      (N121)? data_i[1867] : 
                      (N123)? data_i[1995] : 
                      (N94)? data_i[2123] : 
                      (N96)? data_i[2251] : 
                      (N98)? data_i[2379] : 
                      (N100)? data_i[2507] : 
                      (N102)? data_i[2635] : 
                      (N104)? data_i[2763] : 
                      (N106)? data_i[2891] : 
                      (N108)? data_i[3019] : 
                      (N110)? data_i[3147] : 
                      (N112)? data_i[3275] : 
                      (N114)? data_i[3403] : 
                      (N116)? data_i[3531] : 
                      (N118)? data_i[3659] : 
                      (N120)? data_i[3787] : 
                      (N122)? data_i[3915] : 
                      (N124)? data_i[4043] : 1'b0;
  assign data_o[74] = (N93)? data_i[74] : 
                      (N95)? data_i[202] : 
                      (N97)? data_i[330] : 
                      (N99)? data_i[458] : 
                      (N101)? data_i[586] : 
                      (N103)? data_i[714] : 
                      (N105)? data_i[842] : 
                      (N107)? data_i[970] : 
                      (N109)? data_i[1098] : 
                      (N111)? data_i[1226] : 
                      (N113)? data_i[1354] : 
                      (N115)? data_i[1482] : 
                      (N117)? data_i[1610] : 
                      (N119)? data_i[1738] : 
                      (N121)? data_i[1866] : 
                      (N123)? data_i[1994] : 
                      (N94)? data_i[2122] : 
                      (N96)? data_i[2250] : 
                      (N98)? data_i[2378] : 
                      (N100)? data_i[2506] : 
                      (N102)? data_i[2634] : 
                      (N104)? data_i[2762] : 
                      (N106)? data_i[2890] : 
                      (N108)? data_i[3018] : 
                      (N110)? data_i[3146] : 
                      (N112)? data_i[3274] : 
                      (N114)? data_i[3402] : 
                      (N116)? data_i[3530] : 
                      (N118)? data_i[3658] : 
                      (N120)? data_i[3786] : 
                      (N122)? data_i[3914] : 
                      (N124)? data_i[4042] : 1'b0;
  assign data_o[73] = (N93)? data_i[73] : 
                      (N95)? data_i[201] : 
                      (N97)? data_i[329] : 
                      (N99)? data_i[457] : 
                      (N101)? data_i[585] : 
                      (N103)? data_i[713] : 
                      (N105)? data_i[841] : 
                      (N107)? data_i[969] : 
                      (N109)? data_i[1097] : 
                      (N111)? data_i[1225] : 
                      (N113)? data_i[1353] : 
                      (N115)? data_i[1481] : 
                      (N117)? data_i[1609] : 
                      (N119)? data_i[1737] : 
                      (N121)? data_i[1865] : 
                      (N123)? data_i[1993] : 
                      (N94)? data_i[2121] : 
                      (N96)? data_i[2249] : 
                      (N98)? data_i[2377] : 
                      (N100)? data_i[2505] : 
                      (N102)? data_i[2633] : 
                      (N104)? data_i[2761] : 
                      (N106)? data_i[2889] : 
                      (N108)? data_i[3017] : 
                      (N110)? data_i[3145] : 
                      (N112)? data_i[3273] : 
                      (N114)? data_i[3401] : 
                      (N116)? data_i[3529] : 
                      (N118)? data_i[3657] : 
                      (N120)? data_i[3785] : 
                      (N122)? data_i[3913] : 
                      (N124)? data_i[4041] : 1'b0;
  assign data_o[72] = (N93)? data_i[72] : 
                      (N95)? data_i[200] : 
                      (N97)? data_i[328] : 
                      (N99)? data_i[456] : 
                      (N101)? data_i[584] : 
                      (N103)? data_i[712] : 
                      (N105)? data_i[840] : 
                      (N107)? data_i[968] : 
                      (N109)? data_i[1096] : 
                      (N111)? data_i[1224] : 
                      (N113)? data_i[1352] : 
                      (N115)? data_i[1480] : 
                      (N117)? data_i[1608] : 
                      (N119)? data_i[1736] : 
                      (N121)? data_i[1864] : 
                      (N123)? data_i[1992] : 
                      (N94)? data_i[2120] : 
                      (N96)? data_i[2248] : 
                      (N98)? data_i[2376] : 
                      (N100)? data_i[2504] : 
                      (N102)? data_i[2632] : 
                      (N104)? data_i[2760] : 
                      (N106)? data_i[2888] : 
                      (N108)? data_i[3016] : 
                      (N110)? data_i[3144] : 
                      (N112)? data_i[3272] : 
                      (N114)? data_i[3400] : 
                      (N116)? data_i[3528] : 
                      (N118)? data_i[3656] : 
                      (N120)? data_i[3784] : 
                      (N122)? data_i[3912] : 
                      (N124)? data_i[4040] : 1'b0;
  assign data_o[71] = (N93)? data_i[71] : 
                      (N95)? data_i[199] : 
                      (N97)? data_i[327] : 
                      (N99)? data_i[455] : 
                      (N101)? data_i[583] : 
                      (N103)? data_i[711] : 
                      (N105)? data_i[839] : 
                      (N107)? data_i[967] : 
                      (N109)? data_i[1095] : 
                      (N111)? data_i[1223] : 
                      (N113)? data_i[1351] : 
                      (N115)? data_i[1479] : 
                      (N117)? data_i[1607] : 
                      (N119)? data_i[1735] : 
                      (N121)? data_i[1863] : 
                      (N123)? data_i[1991] : 
                      (N94)? data_i[2119] : 
                      (N96)? data_i[2247] : 
                      (N98)? data_i[2375] : 
                      (N100)? data_i[2503] : 
                      (N102)? data_i[2631] : 
                      (N104)? data_i[2759] : 
                      (N106)? data_i[2887] : 
                      (N108)? data_i[3015] : 
                      (N110)? data_i[3143] : 
                      (N112)? data_i[3271] : 
                      (N114)? data_i[3399] : 
                      (N116)? data_i[3527] : 
                      (N118)? data_i[3655] : 
                      (N120)? data_i[3783] : 
                      (N122)? data_i[3911] : 
                      (N124)? data_i[4039] : 1'b0;
  assign data_o[70] = (N93)? data_i[70] : 
                      (N95)? data_i[198] : 
                      (N97)? data_i[326] : 
                      (N99)? data_i[454] : 
                      (N101)? data_i[582] : 
                      (N103)? data_i[710] : 
                      (N105)? data_i[838] : 
                      (N107)? data_i[966] : 
                      (N109)? data_i[1094] : 
                      (N111)? data_i[1222] : 
                      (N113)? data_i[1350] : 
                      (N115)? data_i[1478] : 
                      (N117)? data_i[1606] : 
                      (N119)? data_i[1734] : 
                      (N121)? data_i[1862] : 
                      (N123)? data_i[1990] : 
                      (N94)? data_i[2118] : 
                      (N96)? data_i[2246] : 
                      (N98)? data_i[2374] : 
                      (N100)? data_i[2502] : 
                      (N102)? data_i[2630] : 
                      (N104)? data_i[2758] : 
                      (N106)? data_i[2886] : 
                      (N108)? data_i[3014] : 
                      (N110)? data_i[3142] : 
                      (N112)? data_i[3270] : 
                      (N114)? data_i[3398] : 
                      (N116)? data_i[3526] : 
                      (N118)? data_i[3654] : 
                      (N120)? data_i[3782] : 
                      (N122)? data_i[3910] : 
                      (N124)? data_i[4038] : 1'b0;
  assign data_o[69] = (N93)? data_i[69] : 
                      (N95)? data_i[197] : 
                      (N97)? data_i[325] : 
                      (N99)? data_i[453] : 
                      (N101)? data_i[581] : 
                      (N103)? data_i[709] : 
                      (N105)? data_i[837] : 
                      (N107)? data_i[965] : 
                      (N109)? data_i[1093] : 
                      (N111)? data_i[1221] : 
                      (N113)? data_i[1349] : 
                      (N115)? data_i[1477] : 
                      (N117)? data_i[1605] : 
                      (N119)? data_i[1733] : 
                      (N121)? data_i[1861] : 
                      (N123)? data_i[1989] : 
                      (N94)? data_i[2117] : 
                      (N96)? data_i[2245] : 
                      (N98)? data_i[2373] : 
                      (N100)? data_i[2501] : 
                      (N102)? data_i[2629] : 
                      (N104)? data_i[2757] : 
                      (N106)? data_i[2885] : 
                      (N108)? data_i[3013] : 
                      (N110)? data_i[3141] : 
                      (N112)? data_i[3269] : 
                      (N114)? data_i[3397] : 
                      (N116)? data_i[3525] : 
                      (N118)? data_i[3653] : 
                      (N120)? data_i[3781] : 
                      (N122)? data_i[3909] : 
                      (N124)? data_i[4037] : 1'b0;
  assign data_o[68] = (N93)? data_i[68] : 
                      (N95)? data_i[196] : 
                      (N97)? data_i[324] : 
                      (N99)? data_i[452] : 
                      (N101)? data_i[580] : 
                      (N103)? data_i[708] : 
                      (N105)? data_i[836] : 
                      (N107)? data_i[964] : 
                      (N109)? data_i[1092] : 
                      (N111)? data_i[1220] : 
                      (N113)? data_i[1348] : 
                      (N115)? data_i[1476] : 
                      (N117)? data_i[1604] : 
                      (N119)? data_i[1732] : 
                      (N121)? data_i[1860] : 
                      (N123)? data_i[1988] : 
                      (N94)? data_i[2116] : 
                      (N96)? data_i[2244] : 
                      (N98)? data_i[2372] : 
                      (N100)? data_i[2500] : 
                      (N102)? data_i[2628] : 
                      (N104)? data_i[2756] : 
                      (N106)? data_i[2884] : 
                      (N108)? data_i[3012] : 
                      (N110)? data_i[3140] : 
                      (N112)? data_i[3268] : 
                      (N114)? data_i[3396] : 
                      (N116)? data_i[3524] : 
                      (N118)? data_i[3652] : 
                      (N120)? data_i[3780] : 
                      (N122)? data_i[3908] : 
                      (N124)? data_i[4036] : 1'b0;
  assign data_o[67] = (N93)? data_i[67] : 
                      (N95)? data_i[195] : 
                      (N97)? data_i[323] : 
                      (N99)? data_i[451] : 
                      (N101)? data_i[579] : 
                      (N103)? data_i[707] : 
                      (N105)? data_i[835] : 
                      (N107)? data_i[963] : 
                      (N109)? data_i[1091] : 
                      (N111)? data_i[1219] : 
                      (N113)? data_i[1347] : 
                      (N115)? data_i[1475] : 
                      (N117)? data_i[1603] : 
                      (N119)? data_i[1731] : 
                      (N121)? data_i[1859] : 
                      (N123)? data_i[1987] : 
                      (N94)? data_i[2115] : 
                      (N96)? data_i[2243] : 
                      (N98)? data_i[2371] : 
                      (N100)? data_i[2499] : 
                      (N102)? data_i[2627] : 
                      (N104)? data_i[2755] : 
                      (N106)? data_i[2883] : 
                      (N108)? data_i[3011] : 
                      (N110)? data_i[3139] : 
                      (N112)? data_i[3267] : 
                      (N114)? data_i[3395] : 
                      (N116)? data_i[3523] : 
                      (N118)? data_i[3651] : 
                      (N120)? data_i[3779] : 
                      (N122)? data_i[3907] : 
                      (N124)? data_i[4035] : 1'b0;
  assign data_o[66] = (N93)? data_i[66] : 
                      (N95)? data_i[194] : 
                      (N97)? data_i[322] : 
                      (N99)? data_i[450] : 
                      (N101)? data_i[578] : 
                      (N103)? data_i[706] : 
                      (N105)? data_i[834] : 
                      (N107)? data_i[962] : 
                      (N109)? data_i[1090] : 
                      (N111)? data_i[1218] : 
                      (N113)? data_i[1346] : 
                      (N115)? data_i[1474] : 
                      (N117)? data_i[1602] : 
                      (N119)? data_i[1730] : 
                      (N121)? data_i[1858] : 
                      (N123)? data_i[1986] : 
                      (N94)? data_i[2114] : 
                      (N96)? data_i[2242] : 
                      (N98)? data_i[2370] : 
                      (N100)? data_i[2498] : 
                      (N102)? data_i[2626] : 
                      (N104)? data_i[2754] : 
                      (N106)? data_i[2882] : 
                      (N108)? data_i[3010] : 
                      (N110)? data_i[3138] : 
                      (N112)? data_i[3266] : 
                      (N114)? data_i[3394] : 
                      (N116)? data_i[3522] : 
                      (N118)? data_i[3650] : 
                      (N120)? data_i[3778] : 
                      (N122)? data_i[3906] : 
                      (N124)? data_i[4034] : 1'b0;
  assign data_o[65] = (N93)? data_i[65] : 
                      (N95)? data_i[193] : 
                      (N97)? data_i[321] : 
                      (N99)? data_i[449] : 
                      (N101)? data_i[577] : 
                      (N103)? data_i[705] : 
                      (N105)? data_i[833] : 
                      (N107)? data_i[961] : 
                      (N109)? data_i[1089] : 
                      (N111)? data_i[1217] : 
                      (N113)? data_i[1345] : 
                      (N115)? data_i[1473] : 
                      (N117)? data_i[1601] : 
                      (N119)? data_i[1729] : 
                      (N121)? data_i[1857] : 
                      (N123)? data_i[1985] : 
                      (N94)? data_i[2113] : 
                      (N96)? data_i[2241] : 
                      (N98)? data_i[2369] : 
                      (N100)? data_i[2497] : 
                      (N102)? data_i[2625] : 
                      (N104)? data_i[2753] : 
                      (N106)? data_i[2881] : 
                      (N108)? data_i[3009] : 
                      (N110)? data_i[3137] : 
                      (N112)? data_i[3265] : 
                      (N114)? data_i[3393] : 
                      (N116)? data_i[3521] : 
                      (N118)? data_i[3649] : 
                      (N120)? data_i[3777] : 
                      (N122)? data_i[3905] : 
                      (N124)? data_i[4033] : 1'b0;
  assign data_o[64] = (N93)? data_i[64] : 
                      (N95)? data_i[192] : 
                      (N97)? data_i[320] : 
                      (N99)? data_i[448] : 
                      (N101)? data_i[576] : 
                      (N103)? data_i[704] : 
                      (N105)? data_i[832] : 
                      (N107)? data_i[960] : 
                      (N109)? data_i[1088] : 
                      (N111)? data_i[1216] : 
                      (N113)? data_i[1344] : 
                      (N115)? data_i[1472] : 
                      (N117)? data_i[1600] : 
                      (N119)? data_i[1728] : 
                      (N121)? data_i[1856] : 
                      (N123)? data_i[1984] : 
                      (N94)? data_i[2112] : 
                      (N96)? data_i[2240] : 
                      (N98)? data_i[2368] : 
                      (N100)? data_i[2496] : 
                      (N102)? data_i[2624] : 
                      (N104)? data_i[2752] : 
                      (N106)? data_i[2880] : 
                      (N108)? data_i[3008] : 
                      (N110)? data_i[3136] : 
                      (N112)? data_i[3264] : 
                      (N114)? data_i[3392] : 
                      (N116)? data_i[3520] : 
                      (N118)? data_i[3648] : 
                      (N120)? data_i[3776] : 
                      (N122)? data_i[3904] : 
                      (N124)? data_i[4032] : 1'b0;
  assign data_o[63] = (N93)? data_i[63] : 
                      (N95)? data_i[191] : 
                      (N97)? data_i[319] : 
                      (N99)? data_i[447] : 
                      (N101)? data_i[575] : 
                      (N103)? data_i[703] : 
                      (N105)? data_i[831] : 
                      (N107)? data_i[959] : 
                      (N109)? data_i[1087] : 
                      (N111)? data_i[1215] : 
                      (N113)? data_i[1343] : 
                      (N115)? data_i[1471] : 
                      (N117)? data_i[1599] : 
                      (N119)? data_i[1727] : 
                      (N121)? data_i[1855] : 
                      (N123)? data_i[1983] : 
                      (N94)? data_i[2111] : 
                      (N96)? data_i[2239] : 
                      (N98)? data_i[2367] : 
                      (N100)? data_i[2495] : 
                      (N102)? data_i[2623] : 
                      (N104)? data_i[2751] : 
                      (N106)? data_i[2879] : 
                      (N108)? data_i[3007] : 
                      (N110)? data_i[3135] : 
                      (N112)? data_i[3263] : 
                      (N114)? data_i[3391] : 
                      (N116)? data_i[3519] : 
                      (N118)? data_i[3647] : 
                      (N120)? data_i[3775] : 
                      (N122)? data_i[3903] : 
                      (N124)? data_i[4031] : 1'b0;
  assign data_o[62] = (N93)? data_i[62] : 
                      (N95)? data_i[190] : 
                      (N97)? data_i[318] : 
                      (N99)? data_i[446] : 
                      (N101)? data_i[574] : 
                      (N103)? data_i[702] : 
                      (N105)? data_i[830] : 
                      (N107)? data_i[958] : 
                      (N109)? data_i[1086] : 
                      (N111)? data_i[1214] : 
                      (N113)? data_i[1342] : 
                      (N115)? data_i[1470] : 
                      (N117)? data_i[1598] : 
                      (N119)? data_i[1726] : 
                      (N121)? data_i[1854] : 
                      (N123)? data_i[1982] : 
                      (N94)? data_i[2110] : 
                      (N96)? data_i[2238] : 
                      (N98)? data_i[2366] : 
                      (N100)? data_i[2494] : 
                      (N102)? data_i[2622] : 
                      (N104)? data_i[2750] : 
                      (N106)? data_i[2878] : 
                      (N108)? data_i[3006] : 
                      (N110)? data_i[3134] : 
                      (N112)? data_i[3262] : 
                      (N114)? data_i[3390] : 
                      (N116)? data_i[3518] : 
                      (N118)? data_i[3646] : 
                      (N120)? data_i[3774] : 
                      (N122)? data_i[3902] : 
                      (N124)? data_i[4030] : 1'b0;
  assign data_o[61] = (N93)? data_i[61] : 
                      (N95)? data_i[189] : 
                      (N97)? data_i[317] : 
                      (N99)? data_i[445] : 
                      (N101)? data_i[573] : 
                      (N103)? data_i[701] : 
                      (N105)? data_i[829] : 
                      (N107)? data_i[957] : 
                      (N109)? data_i[1085] : 
                      (N111)? data_i[1213] : 
                      (N113)? data_i[1341] : 
                      (N115)? data_i[1469] : 
                      (N117)? data_i[1597] : 
                      (N119)? data_i[1725] : 
                      (N121)? data_i[1853] : 
                      (N123)? data_i[1981] : 
                      (N94)? data_i[2109] : 
                      (N96)? data_i[2237] : 
                      (N98)? data_i[2365] : 
                      (N100)? data_i[2493] : 
                      (N102)? data_i[2621] : 
                      (N104)? data_i[2749] : 
                      (N106)? data_i[2877] : 
                      (N108)? data_i[3005] : 
                      (N110)? data_i[3133] : 
                      (N112)? data_i[3261] : 
                      (N114)? data_i[3389] : 
                      (N116)? data_i[3517] : 
                      (N118)? data_i[3645] : 
                      (N120)? data_i[3773] : 
                      (N122)? data_i[3901] : 
                      (N124)? data_i[4029] : 1'b0;
  assign data_o[60] = (N93)? data_i[60] : 
                      (N95)? data_i[188] : 
                      (N97)? data_i[316] : 
                      (N99)? data_i[444] : 
                      (N101)? data_i[572] : 
                      (N103)? data_i[700] : 
                      (N105)? data_i[828] : 
                      (N107)? data_i[956] : 
                      (N109)? data_i[1084] : 
                      (N111)? data_i[1212] : 
                      (N113)? data_i[1340] : 
                      (N115)? data_i[1468] : 
                      (N117)? data_i[1596] : 
                      (N119)? data_i[1724] : 
                      (N121)? data_i[1852] : 
                      (N123)? data_i[1980] : 
                      (N94)? data_i[2108] : 
                      (N96)? data_i[2236] : 
                      (N98)? data_i[2364] : 
                      (N100)? data_i[2492] : 
                      (N102)? data_i[2620] : 
                      (N104)? data_i[2748] : 
                      (N106)? data_i[2876] : 
                      (N108)? data_i[3004] : 
                      (N110)? data_i[3132] : 
                      (N112)? data_i[3260] : 
                      (N114)? data_i[3388] : 
                      (N116)? data_i[3516] : 
                      (N118)? data_i[3644] : 
                      (N120)? data_i[3772] : 
                      (N122)? data_i[3900] : 
                      (N124)? data_i[4028] : 1'b0;
  assign data_o[59] = (N93)? data_i[59] : 
                      (N95)? data_i[187] : 
                      (N97)? data_i[315] : 
                      (N99)? data_i[443] : 
                      (N101)? data_i[571] : 
                      (N103)? data_i[699] : 
                      (N105)? data_i[827] : 
                      (N107)? data_i[955] : 
                      (N109)? data_i[1083] : 
                      (N111)? data_i[1211] : 
                      (N113)? data_i[1339] : 
                      (N115)? data_i[1467] : 
                      (N117)? data_i[1595] : 
                      (N119)? data_i[1723] : 
                      (N121)? data_i[1851] : 
                      (N123)? data_i[1979] : 
                      (N94)? data_i[2107] : 
                      (N96)? data_i[2235] : 
                      (N98)? data_i[2363] : 
                      (N100)? data_i[2491] : 
                      (N102)? data_i[2619] : 
                      (N104)? data_i[2747] : 
                      (N106)? data_i[2875] : 
                      (N108)? data_i[3003] : 
                      (N110)? data_i[3131] : 
                      (N112)? data_i[3259] : 
                      (N114)? data_i[3387] : 
                      (N116)? data_i[3515] : 
                      (N118)? data_i[3643] : 
                      (N120)? data_i[3771] : 
                      (N122)? data_i[3899] : 
                      (N124)? data_i[4027] : 1'b0;
  assign data_o[58] = (N93)? data_i[58] : 
                      (N95)? data_i[186] : 
                      (N97)? data_i[314] : 
                      (N99)? data_i[442] : 
                      (N101)? data_i[570] : 
                      (N103)? data_i[698] : 
                      (N105)? data_i[826] : 
                      (N107)? data_i[954] : 
                      (N109)? data_i[1082] : 
                      (N111)? data_i[1210] : 
                      (N113)? data_i[1338] : 
                      (N115)? data_i[1466] : 
                      (N117)? data_i[1594] : 
                      (N119)? data_i[1722] : 
                      (N121)? data_i[1850] : 
                      (N123)? data_i[1978] : 
                      (N94)? data_i[2106] : 
                      (N96)? data_i[2234] : 
                      (N98)? data_i[2362] : 
                      (N100)? data_i[2490] : 
                      (N102)? data_i[2618] : 
                      (N104)? data_i[2746] : 
                      (N106)? data_i[2874] : 
                      (N108)? data_i[3002] : 
                      (N110)? data_i[3130] : 
                      (N112)? data_i[3258] : 
                      (N114)? data_i[3386] : 
                      (N116)? data_i[3514] : 
                      (N118)? data_i[3642] : 
                      (N120)? data_i[3770] : 
                      (N122)? data_i[3898] : 
                      (N124)? data_i[4026] : 1'b0;
  assign data_o[57] = (N93)? data_i[57] : 
                      (N95)? data_i[185] : 
                      (N97)? data_i[313] : 
                      (N99)? data_i[441] : 
                      (N101)? data_i[569] : 
                      (N103)? data_i[697] : 
                      (N105)? data_i[825] : 
                      (N107)? data_i[953] : 
                      (N109)? data_i[1081] : 
                      (N111)? data_i[1209] : 
                      (N113)? data_i[1337] : 
                      (N115)? data_i[1465] : 
                      (N117)? data_i[1593] : 
                      (N119)? data_i[1721] : 
                      (N121)? data_i[1849] : 
                      (N123)? data_i[1977] : 
                      (N94)? data_i[2105] : 
                      (N96)? data_i[2233] : 
                      (N98)? data_i[2361] : 
                      (N100)? data_i[2489] : 
                      (N102)? data_i[2617] : 
                      (N104)? data_i[2745] : 
                      (N106)? data_i[2873] : 
                      (N108)? data_i[3001] : 
                      (N110)? data_i[3129] : 
                      (N112)? data_i[3257] : 
                      (N114)? data_i[3385] : 
                      (N116)? data_i[3513] : 
                      (N118)? data_i[3641] : 
                      (N120)? data_i[3769] : 
                      (N122)? data_i[3897] : 
                      (N124)? data_i[4025] : 1'b0;
  assign data_o[56] = (N93)? data_i[56] : 
                      (N95)? data_i[184] : 
                      (N97)? data_i[312] : 
                      (N99)? data_i[440] : 
                      (N101)? data_i[568] : 
                      (N103)? data_i[696] : 
                      (N105)? data_i[824] : 
                      (N107)? data_i[952] : 
                      (N109)? data_i[1080] : 
                      (N111)? data_i[1208] : 
                      (N113)? data_i[1336] : 
                      (N115)? data_i[1464] : 
                      (N117)? data_i[1592] : 
                      (N119)? data_i[1720] : 
                      (N121)? data_i[1848] : 
                      (N123)? data_i[1976] : 
                      (N94)? data_i[2104] : 
                      (N96)? data_i[2232] : 
                      (N98)? data_i[2360] : 
                      (N100)? data_i[2488] : 
                      (N102)? data_i[2616] : 
                      (N104)? data_i[2744] : 
                      (N106)? data_i[2872] : 
                      (N108)? data_i[3000] : 
                      (N110)? data_i[3128] : 
                      (N112)? data_i[3256] : 
                      (N114)? data_i[3384] : 
                      (N116)? data_i[3512] : 
                      (N118)? data_i[3640] : 
                      (N120)? data_i[3768] : 
                      (N122)? data_i[3896] : 
                      (N124)? data_i[4024] : 1'b0;
  assign data_o[55] = (N93)? data_i[55] : 
                      (N95)? data_i[183] : 
                      (N97)? data_i[311] : 
                      (N99)? data_i[439] : 
                      (N101)? data_i[567] : 
                      (N103)? data_i[695] : 
                      (N105)? data_i[823] : 
                      (N107)? data_i[951] : 
                      (N109)? data_i[1079] : 
                      (N111)? data_i[1207] : 
                      (N113)? data_i[1335] : 
                      (N115)? data_i[1463] : 
                      (N117)? data_i[1591] : 
                      (N119)? data_i[1719] : 
                      (N121)? data_i[1847] : 
                      (N123)? data_i[1975] : 
                      (N94)? data_i[2103] : 
                      (N96)? data_i[2231] : 
                      (N98)? data_i[2359] : 
                      (N100)? data_i[2487] : 
                      (N102)? data_i[2615] : 
                      (N104)? data_i[2743] : 
                      (N106)? data_i[2871] : 
                      (N108)? data_i[2999] : 
                      (N110)? data_i[3127] : 
                      (N112)? data_i[3255] : 
                      (N114)? data_i[3383] : 
                      (N116)? data_i[3511] : 
                      (N118)? data_i[3639] : 
                      (N120)? data_i[3767] : 
                      (N122)? data_i[3895] : 
                      (N124)? data_i[4023] : 1'b0;
  assign data_o[54] = (N93)? data_i[54] : 
                      (N95)? data_i[182] : 
                      (N97)? data_i[310] : 
                      (N99)? data_i[438] : 
                      (N101)? data_i[566] : 
                      (N103)? data_i[694] : 
                      (N105)? data_i[822] : 
                      (N107)? data_i[950] : 
                      (N109)? data_i[1078] : 
                      (N111)? data_i[1206] : 
                      (N113)? data_i[1334] : 
                      (N115)? data_i[1462] : 
                      (N117)? data_i[1590] : 
                      (N119)? data_i[1718] : 
                      (N121)? data_i[1846] : 
                      (N123)? data_i[1974] : 
                      (N94)? data_i[2102] : 
                      (N96)? data_i[2230] : 
                      (N98)? data_i[2358] : 
                      (N100)? data_i[2486] : 
                      (N102)? data_i[2614] : 
                      (N104)? data_i[2742] : 
                      (N106)? data_i[2870] : 
                      (N108)? data_i[2998] : 
                      (N110)? data_i[3126] : 
                      (N112)? data_i[3254] : 
                      (N114)? data_i[3382] : 
                      (N116)? data_i[3510] : 
                      (N118)? data_i[3638] : 
                      (N120)? data_i[3766] : 
                      (N122)? data_i[3894] : 
                      (N124)? data_i[4022] : 1'b0;
  assign data_o[53] = (N93)? data_i[53] : 
                      (N95)? data_i[181] : 
                      (N97)? data_i[309] : 
                      (N99)? data_i[437] : 
                      (N101)? data_i[565] : 
                      (N103)? data_i[693] : 
                      (N105)? data_i[821] : 
                      (N107)? data_i[949] : 
                      (N109)? data_i[1077] : 
                      (N111)? data_i[1205] : 
                      (N113)? data_i[1333] : 
                      (N115)? data_i[1461] : 
                      (N117)? data_i[1589] : 
                      (N119)? data_i[1717] : 
                      (N121)? data_i[1845] : 
                      (N123)? data_i[1973] : 
                      (N94)? data_i[2101] : 
                      (N96)? data_i[2229] : 
                      (N98)? data_i[2357] : 
                      (N100)? data_i[2485] : 
                      (N102)? data_i[2613] : 
                      (N104)? data_i[2741] : 
                      (N106)? data_i[2869] : 
                      (N108)? data_i[2997] : 
                      (N110)? data_i[3125] : 
                      (N112)? data_i[3253] : 
                      (N114)? data_i[3381] : 
                      (N116)? data_i[3509] : 
                      (N118)? data_i[3637] : 
                      (N120)? data_i[3765] : 
                      (N122)? data_i[3893] : 
                      (N124)? data_i[4021] : 1'b0;
  assign data_o[52] = (N93)? data_i[52] : 
                      (N95)? data_i[180] : 
                      (N97)? data_i[308] : 
                      (N99)? data_i[436] : 
                      (N101)? data_i[564] : 
                      (N103)? data_i[692] : 
                      (N105)? data_i[820] : 
                      (N107)? data_i[948] : 
                      (N109)? data_i[1076] : 
                      (N111)? data_i[1204] : 
                      (N113)? data_i[1332] : 
                      (N115)? data_i[1460] : 
                      (N117)? data_i[1588] : 
                      (N119)? data_i[1716] : 
                      (N121)? data_i[1844] : 
                      (N123)? data_i[1972] : 
                      (N94)? data_i[2100] : 
                      (N96)? data_i[2228] : 
                      (N98)? data_i[2356] : 
                      (N100)? data_i[2484] : 
                      (N102)? data_i[2612] : 
                      (N104)? data_i[2740] : 
                      (N106)? data_i[2868] : 
                      (N108)? data_i[2996] : 
                      (N110)? data_i[3124] : 
                      (N112)? data_i[3252] : 
                      (N114)? data_i[3380] : 
                      (N116)? data_i[3508] : 
                      (N118)? data_i[3636] : 
                      (N120)? data_i[3764] : 
                      (N122)? data_i[3892] : 
                      (N124)? data_i[4020] : 1'b0;
  assign data_o[51] = (N93)? data_i[51] : 
                      (N95)? data_i[179] : 
                      (N97)? data_i[307] : 
                      (N99)? data_i[435] : 
                      (N101)? data_i[563] : 
                      (N103)? data_i[691] : 
                      (N105)? data_i[819] : 
                      (N107)? data_i[947] : 
                      (N109)? data_i[1075] : 
                      (N111)? data_i[1203] : 
                      (N113)? data_i[1331] : 
                      (N115)? data_i[1459] : 
                      (N117)? data_i[1587] : 
                      (N119)? data_i[1715] : 
                      (N121)? data_i[1843] : 
                      (N123)? data_i[1971] : 
                      (N94)? data_i[2099] : 
                      (N96)? data_i[2227] : 
                      (N98)? data_i[2355] : 
                      (N100)? data_i[2483] : 
                      (N102)? data_i[2611] : 
                      (N104)? data_i[2739] : 
                      (N106)? data_i[2867] : 
                      (N108)? data_i[2995] : 
                      (N110)? data_i[3123] : 
                      (N112)? data_i[3251] : 
                      (N114)? data_i[3379] : 
                      (N116)? data_i[3507] : 
                      (N118)? data_i[3635] : 
                      (N120)? data_i[3763] : 
                      (N122)? data_i[3891] : 
                      (N124)? data_i[4019] : 1'b0;
  assign data_o[50] = (N93)? data_i[50] : 
                      (N95)? data_i[178] : 
                      (N97)? data_i[306] : 
                      (N99)? data_i[434] : 
                      (N101)? data_i[562] : 
                      (N103)? data_i[690] : 
                      (N105)? data_i[818] : 
                      (N107)? data_i[946] : 
                      (N109)? data_i[1074] : 
                      (N111)? data_i[1202] : 
                      (N113)? data_i[1330] : 
                      (N115)? data_i[1458] : 
                      (N117)? data_i[1586] : 
                      (N119)? data_i[1714] : 
                      (N121)? data_i[1842] : 
                      (N123)? data_i[1970] : 
                      (N94)? data_i[2098] : 
                      (N96)? data_i[2226] : 
                      (N98)? data_i[2354] : 
                      (N100)? data_i[2482] : 
                      (N102)? data_i[2610] : 
                      (N104)? data_i[2738] : 
                      (N106)? data_i[2866] : 
                      (N108)? data_i[2994] : 
                      (N110)? data_i[3122] : 
                      (N112)? data_i[3250] : 
                      (N114)? data_i[3378] : 
                      (N116)? data_i[3506] : 
                      (N118)? data_i[3634] : 
                      (N120)? data_i[3762] : 
                      (N122)? data_i[3890] : 
                      (N124)? data_i[4018] : 1'b0;
  assign data_o[49] = (N93)? data_i[49] : 
                      (N95)? data_i[177] : 
                      (N97)? data_i[305] : 
                      (N99)? data_i[433] : 
                      (N101)? data_i[561] : 
                      (N103)? data_i[689] : 
                      (N105)? data_i[817] : 
                      (N107)? data_i[945] : 
                      (N109)? data_i[1073] : 
                      (N111)? data_i[1201] : 
                      (N113)? data_i[1329] : 
                      (N115)? data_i[1457] : 
                      (N117)? data_i[1585] : 
                      (N119)? data_i[1713] : 
                      (N121)? data_i[1841] : 
                      (N123)? data_i[1969] : 
                      (N94)? data_i[2097] : 
                      (N96)? data_i[2225] : 
                      (N98)? data_i[2353] : 
                      (N100)? data_i[2481] : 
                      (N102)? data_i[2609] : 
                      (N104)? data_i[2737] : 
                      (N106)? data_i[2865] : 
                      (N108)? data_i[2993] : 
                      (N110)? data_i[3121] : 
                      (N112)? data_i[3249] : 
                      (N114)? data_i[3377] : 
                      (N116)? data_i[3505] : 
                      (N118)? data_i[3633] : 
                      (N120)? data_i[3761] : 
                      (N122)? data_i[3889] : 
                      (N124)? data_i[4017] : 1'b0;
  assign data_o[48] = (N93)? data_i[48] : 
                      (N95)? data_i[176] : 
                      (N97)? data_i[304] : 
                      (N99)? data_i[432] : 
                      (N101)? data_i[560] : 
                      (N103)? data_i[688] : 
                      (N105)? data_i[816] : 
                      (N107)? data_i[944] : 
                      (N109)? data_i[1072] : 
                      (N111)? data_i[1200] : 
                      (N113)? data_i[1328] : 
                      (N115)? data_i[1456] : 
                      (N117)? data_i[1584] : 
                      (N119)? data_i[1712] : 
                      (N121)? data_i[1840] : 
                      (N123)? data_i[1968] : 
                      (N94)? data_i[2096] : 
                      (N96)? data_i[2224] : 
                      (N98)? data_i[2352] : 
                      (N100)? data_i[2480] : 
                      (N102)? data_i[2608] : 
                      (N104)? data_i[2736] : 
                      (N106)? data_i[2864] : 
                      (N108)? data_i[2992] : 
                      (N110)? data_i[3120] : 
                      (N112)? data_i[3248] : 
                      (N114)? data_i[3376] : 
                      (N116)? data_i[3504] : 
                      (N118)? data_i[3632] : 
                      (N120)? data_i[3760] : 
                      (N122)? data_i[3888] : 
                      (N124)? data_i[4016] : 1'b0;
  assign data_o[47] = (N93)? data_i[47] : 
                      (N95)? data_i[175] : 
                      (N97)? data_i[303] : 
                      (N99)? data_i[431] : 
                      (N101)? data_i[559] : 
                      (N103)? data_i[687] : 
                      (N105)? data_i[815] : 
                      (N107)? data_i[943] : 
                      (N109)? data_i[1071] : 
                      (N111)? data_i[1199] : 
                      (N113)? data_i[1327] : 
                      (N115)? data_i[1455] : 
                      (N117)? data_i[1583] : 
                      (N119)? data_i[1711] : 
                      (N121)? data_i[1839] : 
                      (N123)? data_i[1967] : 
                      (N94)? data_i[2095] : 
                      (N96)? data_i[2223] : 
                      (N98)? data_i[2351] : 
                      (N100)? data_i[2479] : 
                      (N102)? data_i[2607] : 
                      (N104)? data_i[2735] : 
                      (N106)? data_i[2863] : 
                      (N108)? data_i[2991] : 
                      (N110)? data_i[3119] : 
                      (N112)? data_i[3247] : 
                      (N114)? data_i[3375] : 
                      (N116)? data_i[3503] : 
                      (N118)? data_i[3631] : 
                      (N120)? data_i[3759] : 
                      (N122)? data_i[3887] : 
                      (N124)? data_i[4015] : 1'b0;
  assign data_o[46] = (N93)? data_i[46] : 
                      (N95)? data_i[174] : 
                      (N97)? data_i[302] : 
                      (N99)? data_i[430] : 
                      (N101)? data_i[558] : 
                      (N103)? data_i[686] : 
                      (N105)? data_i[814] : 
                      (N107)? data_i[942] : 
                      (N109)? data_i[1070] : 
                      (N111)? data_i[1198] : 
                      (N113)? data_i[1326] : 
                      (N115)? data_i[1454] : 
                      (N117)? data_i[1582] : 
                      (N119)? data_i[1710] : 
                      (N121)? data_i[1838] : 
                      (N123)? data_i[1966] : 
                      (N94)? data_i[2094] : 
                      (N96)? data_i[2222] : 
                      (N98)? data_i[2350] : 
                      (N100)? data_i[2478] : 
                      (N102)? data_i[2606] : 
                      (N104)? data_i[2734] : 
                      (N106)? data_i[2862] : 
                      (N108)? data_i[2990] : 
                      (N110)? data_i[3118] : 
                      (N112)? data_i[3246] : 
                      (N114)? data_i[3374] : 
                      (N116)? data_i[3502] : 
                      (N118)? data_i[3630] : 
                      (N120)? data_i[3758] : 
                      (N122)? data_i[3886] : 
                      (N124)? data_i[4014] : 1'b0;
  assign data_o[45] = (N93)? data_i[45] : 
                      (N95)? data_i[173] : 
                      (N97)? data_i[301] : 
                      (N99)? data_i[429] : 
                      (N101)? data_i[557] : 
                      (N103)? data_i[685] : 
                      (N105)? data_i[813] : 
                      (N107)? data_i[941] : 
                      (N109)? data_i[1069] : 
                      (N111)? data_i[1197] : 
                      (N113)? data_i[1325] : 
                      (N115)? data_i[1453] : 
                      (N117)? data_i[1581] : 
                      (N119)? data_i[1709] : 
                      (N121)? data_i[1837] : 
                      (N123)? data_i[1965] : 
                      (N94)? data_i[2093] : 
                      (N96)? data_i[2221] : 
                      (N98)? data_i[2349] : 
                      (N100)? data_i[2477] : 
                      (N102)? data_i[2605] : 
                      (N104)? data_i[2733] : 
                      (N106)? data_i[2861] : 
                      (N108)? data_i[2989] : 
                      (N110)? data_i[3117] : 
                      (N112)? data_i[3245] : 
                      (N114)? data_i[3373] : 
                      (N116)? data_i[3501] : 
                      (N118)? data_i[3629] : 
                      (N120)? data_i[3757] : 
                      (N122)? data_i[3885] : 
                      (N124)? data_i[4013] : 1'b0;
  assign data_o[44] = (N93)? data_i[44] : 
                      (N95)? data_i[172] : 
                      (N97)? data_i[300] : 
                      (N99)? data_i[428] : 
                      (N101)? data_i[556] : 
                      (N103)? data_i[684] : 
                      (N105)? data_i[812] : 
                      (N107)? data_i[940] : 
                      (N109)? data_i[1068] : 
                      (N111)? data_i[1196] : 
                      (N113)? data_i[1324] : 
                      (N115)? data_i[1452] : 
                      (N117)? data_i[1580] : 
                      (N119)? data_i[1708] : 
                      (N121)? data_i[1836] : 
                      (N123)? data_i[1964] : 
                      (N94)? data_i[2092] : 
                      (N96)? data_i[2220] : 
                      (N98)? data_i[2348] : 
                      (N100)? data_i[2476] : 
                      (N102)? data_i[2604] : 
                      (N104)? data_i[2732] : 
                      (N106)? data_i[2860] : 
                      (N108)? data_i[2988] : 
                      (N110)? data_i[3116] : 
                      (N112)? data_i[3244] : 
                      (N114)? data_i[3372] : 
                      (N116)? data_i[3500] : 
                      (N118)? data_i[3628] : 
                      (N120)? data_i[3756] : 
                      (N122)? data_i[3884] : 
                      (N124)? data_i[4012] : 1'b0;
  assign data_o[43] = (N93)? data_i[43] : 
                      (N95)? data_i[171] : 
                      (N97)? data_i[299] : 
                      (N99)? data_i[427] : 
                      (N101)? data_i[555] : 
                      (N103)? data_i[683] : 
                      (N105)? data_i[811] : 
                      (N107)? data_i[939] : 
                      (N109)? data_i[1067] : 
                      (N111)? data_i[1195] : 
                      (N113)? data_i[1323] : 
                      (N115)? data_i[1451] : 
                      (N117)? data_i[1579] : 
                      (N119)? data_i[1707] : 
                      (N121)? data_i[1835] : 
                      (N123)? data_i[1963] : 
                      (N94)? data_i[2091] : 
                      (N96)? data_i[2219] : 
                      (N98)? data_i[2347] : 
                      (N100)? data_i[2475] : 
                      (N102)? data_i[2603] : 
                      (N104)? data_i[2731] : 
                      (N106)? data_i[2859] : 
                      (N108)? data_i[2987] : 
                      (N110)? data_i[3115] : 
                      (N112)? data_i[3243] : 
                      (N114)? data_i[3371] : 
                      (N116)? data_i[3499] : 
                      (N118)? data_i[3627] : 
                      (N120)? data_i[3755] : 
                      (N122)? data_i[3883] : 
                      (N124)? data_i[4011] : 1'b0;
  assign data_o[42] = (N93)? data_i[42] : 
                      (N95)? data_i[170] : 
                      (N97)? data_i[298] : 
                      (N99)? data_i[426] : 
                      (N101)? data_i[554] : 
                      (N103)? data_i[682] : 
                      (N105)? data_i[810] : 
                      (N107)? data_i[938] : 
                      (N109)? data_i[1066] : 
                      (N111)? data_i[1194] : 
                      (N113)? data_i[1322] : 
                      (N115)? data_i[1450] : 
                      (N117)? data_i[1578] : 
                      (N119)? data_i[1706] : 
                      (N121)? data_i[1834] : 
                      (N123)? data_i[1962] : 
                      (N94)? data_i[2090] : 
                      (N96)? data_i[2218] : 
                      (N98)? data_i[2346] : 
                      (N100)? data_i[2474] : 
                      (N102)? data_i[2602] : 
                      (N104)? data_i[2730] : 
                      (N106)? data_i[2858] : 
                      (N108)? data_i[2986] : 
                      (N110)? data_i[3114] : 
                      (N112)? data_i[3242] : 
                      (N114)? data_i[3370] : 
                      (N116)? data_i[3498] : 
                      (N118)? data_i[3626] : 
                      (N120)? data_i[3754] : 
                      (N122)? data_i[3882] : 
                      (N124)? data_i[4010] : 1'b0;
  assign data_o[41] = (N93)? data_i[41] : 
                      (N95)? data_i[169] : 
                      (N97)? data_i[297] : 
                      (N99)? data_i[425] : 
                      (N101)? data_i[553] : 
                      (N103)? data_i[681] : 
                      (N105)? data_i[809] : 
                      (N107)? data_i[937] : 
                      (N109)? data_i[1065] : 
                      (N111)? data_i[1193] : 
                      (N113)? data_i[1321] : 
                      (N115)? data_i[1449] : 
                      (N117)? data_i[1577] : 
                      (N119)? data_i[1705] : 
                      (N121)? data_i[1833] : 
                      (N123)? data_i[1961] : 
                      (N94)? data_i[2089] : 
                      (N96)? data_i[2217] : 
                      (N98)? data_i[2345] : 
                      (N100)? data_i[2473] : 
                      (N102)? data_i[2601] : 
                      (N104)? data_i[2729] : 
                      (N106)? data_i[2857] : 
                      (N108)? data_i[2985] : 
                      (N110)? data_i[3113] : 
                      (N112)? data_i[3241] : 
                      (N114)? data_i[3369] : 
                      (N116)? data_i[3497] : 
                      (N118)? data_i[3625] : 
                      (N120)? data_i[3753] : 
                      (N122)? data_i[3881] : 
                      (N124)? data_i[4009] : 1'b0;
  assign data_o[40] = (N93)? data_i[40] : 
                      (N95)? data_i[168] : 
                      (N97)? data_i[296] : 
                      (N99)? data_i[424] : 
                      (N101)? data_i[552] : 
                      (N103)? data_i[680] : 
                      (N105)? data_i[808] : 
                      (N107)? data_i[936] : 
                      (N109)? data_i[1064] : 
                      (N111)? data_i[1192] : 
                      (N113)? data_i[1320] : 
                      (N115)? data_i[1448] : 
                      (N117)? data_i[1576] : 
                      (N119)? data_i[1704] : 
                      (N121)? data_i[1832] : 
                      (N123)? data_i[1960] : 
                      (N94)? data_i[2088] : 
                      (N96)? data_i[2216] : 
                      (N98)? data_i[2344] : 
                      (N100)? data_i[2472] : 
                      (N102)? data_i[2600] : 
                      (N104)? data_i[2728] : 
                      (N106)? data_i[2856] : 
                      (N108)? data_i[2984] : 
                      (N110)? data_i[3112] : 
                      (N112)? data_i[3240] : 
                      (N114)? data_i[3368] : 
                      (N116)? data_i[3496] : 
                      (N118)? data_i[3624] : 
                      (N120)? data_i[3752] : 
                      (N122)? data_i[3880] : 
                      (N124)? data_i[4008] : 1'b0;
  assign data_o[39] = (N93)? data_i[39] : 
                      (N95)? data_i[167] : 
                      (N97)? data_i[295] : 
                      (N99)? data_i[423] : 
                      (N101)? data_i[551] : 
                      (N103)? data_i[679] : 
                      (N105)? data_i[807] : 
                      (N107)? data_i[935] : 
                      (N109)? data_i[1063] : 
                      (N111)? data_i[1191] : 
                      (N113)? data_i[1319] : 
                      (N115)? data_i[1447] : 
                      (N117)? data_i[1575] : 
                      (N119)? data_i[1703] : 
                      (N121)? data_i[1831] : 
                      (N123)? data_i[1959] : 
                      (N94)? data_i[2087] : 
                      (N96)? data_i[2215] : 
                      (N98)? data_i[2343] : 
                      (N100)? data_i[2471] : 
                      (N102)? data_i[2599] : 
                      (N104)? data_i[2727] : 
                      (N106)? data_i[2855] : 
                      (N108)? data_i[2983] : 
                      (N110)? data_i[3111] : 
                      (N112)? data_i[3239] : 
                      (N114)? data_i[3367] : 
                      (N116)? data_i[3495] : 
                      (N118)? data_i[3623] : 
                      (N120)? data_i[3751] : 
                      (N122)? data_i[3879] : 
                      (N124)? data_i[4007] : 1'b0;
  assign data_o[38] = (N93)? data_i[38] : 
                      (N95)? data_i[166] : 
                      (N97)? data_i[294] : 
                      (N99)? data_i[422] : 
                      (N101)? data_i[550] : 
                      (N103)? data_i[678] : 
                      (N105)? data_i[806] : 
                      (N107)? data_i[934] : 
                      (N109)? data_i[1062] : 
                      (N111)? data_i[1190] : 
                      (N113)? data_i[1318] : 
                      (N115)? data_i[1446] : 
                      (N117)? data_i[1574] : 
                      (N119)? data_i[1702] : 
                      (N121)? data_i[1830] : 
                      (N123)? data_i[1958] : 
                      (N94)? data_i[2086] : 
                      (N96)? data_i[2214] : 
                      (N98)? data_i[2342] : 
                      (N100)? data_i[2470] : 
                      (N102)? data_i[2598] : 
                      (N104)? data_i[2726] : 
                      (N106)? data_i[2854] : 
                      (N108)? data_i[2982] : 
                      (N110)? data_i[3110] : 
                      (N112)? data_i[3238] : 
                      (N114)? data_i[3366] : 
                      (N116)? data_i[3494] : 
                      (N118)? data_i[3622] : 
                      (N120)? data_i[3750] : 
                      (N122)? data_i[3878] : 
                      (N124)? data_i[4006] : 1'b0;
  assign data_o[37] = (N93)? data_i[37] : 
                      (N95)? data_i[165] : 
                      (N97)? data_i[293] : 
                      (N99)? data_i[421] : 
                      (N101)? data_i[549] : 
                      (N103)? data_i[677] : 
                      (N105)? data_i[805] : 
                      (N107)? data_i[933] : 
                      (N109)? data_i[1061] : 
                      (N111)? data_i[1189] : 
                      (N113)? data_i[1317] : 
                      (N115)? data_i[1445] : 
                      (N117)? data_i[1573] : 
                      (N119)? data_i[1701] : 
                      (N121)? data_i[1829] : 
                      (N123)? data_i[1957] : 
                      (N94)? data_i[2085] : 
                      (N96)? data_i[2213] : 
                      (N98)? data_i[2341] : 
                      (N100)? data_i[2469] : 
                      (N102)? data_i[2597] : 
                      (N104)? data_i[2725] : 
                      (N106)? data_i[2853] : 
                      (N108)? data_i[2981] : 
                      (N110)? data_i[3109] : 
                      (N112)? data_i[3237] : 
                      (N114)? data_i[3365] : 
                      (N116)? data_i[3493] : 
                      (N118)? data_i[3621] : 
                      (N120)? data_i[3749] : 
                      (N122)? data_i[3877] : 
                      (N124)? data_i[4005] : 1'b0;
  assign data_o[36] = (N93)? data_i[36] : 
                      (N95)? data_i[164] : 
                      (N97)? data_i[292] : 
                      (N99)? data_i[420] : 
                      (N101)? data_i[548] : 
                      (N103)? data_i[676] : 
                      (N105)? data_i[804] : 
                      (N107)? data_i[932] : 
                      (N109)? data_i[1060] : 
                      (N111)? data_i[1188] : 
                      (N113)? data_i[1316] : 
                      (N115)? data_i[1444] : 
                      (N117)? data_i[1572] : 
                      (N119)? data_i[1700] : 
                      (N121)? data_i[1828] : 
                      (N123)? data_i[1956] : 
                      (N94)? data_i[2084] : 
                      (N96)? data_i[2212] : 
                      (N98)? data_i[2340] : 
                      (N100)? data_i[2468] : 
                      (N102)? data_i[2596] : 
                      (N104)? data_i[2724] : 
                      (N106)? data_i[2852] : 
                      (N108)? data_i[2980] : 
                      (N110)? data_i[3108] : 
                      (N112)? data_i[3236] : 
                      (N114)? data_i[3364] : 
                      (N116)? data_i[3492] : 
                      (N118)? data_i[3620] : 
                      (N120)? data_i[3748] : 
                      (N122)? data_i[3876] : 
                      (N124)? data_i[4004] : 1'b0;
  assign data_o[35] = (N93)? data_i[35] : 
                      (N95)? data_i[163] : 
                      (N97)? data_i[291] : 
                      (N99)? data_i[419] : 
                      (N101)? data_i[547] : 
                      (N103)? data_i[675] : 
                      (N105)? data_i[803] : 
                      (N107)? data_i[931] : 
                      (N109)? data_i[1059] : 
                      (N111)? data_i[1187] : 
                      (N113)? data_i[1315] : 
                      (N115)? data_i[1443] : 
                      (N117)? data_i[1571] : 
                      (N119)? data_i[1699] : 
                      (N121)? data_i[1827] : 
                      (N123)? data_i[1955] : 
                      (N94)? data_i[2083] : 
                      (N96)? data_i[2211] : 
                      (N98)? data_i[2339] : 
                      (N100)? data_i[2467] : 
                      (N102)? data_i[2595] : 
                      (N104)? data_i[2723] : 
                      (N106)? data_i[2851] : 
                      (N108)? data_i[2979] : 
                      (N110)? data_i[3107] : 
                      (N112)? data_i[3235] : 
                      (N114)? data_i[3363] : 
                      (N116)? data_i[3491] : 
                      (N118)? data_i[3619] : 
                      (N120)? data_i[3747] : 
                      (N122)? data_i[3875] : 
                      (N124)? data_i[4003] : 1'b0;
  assign data_o[34] = (N93)? data_i[34] : 
                      (N95)? data_i[162] : 
                      (N97)? data_i[290] : 
                      (N99)? data_i[418] : 
                      (N101)? data_i[546] : 
                      (N103)? data_i[674] : 
                      (N105)? data_i[802] : 
                      (N107)? data_i[930] : 
                      (N109)? data_i[1058] : 
                      (N111)? data_i[1186] : 
                      (N113)? data_i[1314] : 
                      (N115)? data_i[1442] : 
                      (N117)? data_i[1570] : 
                      (N119)? data_i[1698] : 
                      (N121)? data_i[1826] : 
                      (N123)? data_i[1954] : 
                      (N94)? data_i[2082] : 
                      (N96)? data_i[2210] : 
                      (N98)? data_i[2338] : 
                      (N100)? data_i[2466] : 
                      (N102)? data_i[2594] : 
                      (N104)? data_i[2722] : 
                      (N106)? data_i[2850] : 
                      (N108)? data_i[2978] : 
                      (N110)? data_i[3106] : 
                      (N112)? data_i[3234] : 
                      (N114)? data_i[3362] : 
                      (N116)? data_i[3490] : 
                      (N118)? data_i[3618] : 
                      (N120)? data_i[3746] : 
                      (N122)? data_i[3874] : 
                      (N124)? data_i[4002] : 1'b0;
  assign data_o[33] = (N93)? data_i[33] : 
                      (N95)? data_i[161] : 
                      (N97)? data_i[289] : 
                      (N99)? data_i[417] : 
                      (N101)? data_i[545] : 
                      (N103)? data_i[673] : 
                      (N105)? data_i[801] : 
                      (N107)? data_i[929] : 
                      (N109)? data_i[1057] : 
                      (N111)? data_i[1185] : 
                      (N113)? data_i[1313] : 
                      (N115)? data_i[1441] : 
                      (N117)? data_i[1569] : 
                      (N119)? data_i[1697] : 
                      (N121)? data_i[1825] : 
                      (N123)? data_i[1953] : 
                      (N94)? data_i[2081] : 
                      (N96)? data_i[2209] : 
                      (N98)? data_i[2337] : 
                      (N100)? data_i[2465] : 
                      (N102)? data_i[2593] : 
                      (N104)? data_i[2721] : 
                      (N106)? data_i[2849] : 
                      (N108)? data_i[2977] : 
                      (N110)? data_i[3105] : 
                      (N112)? data_i[3233] : 
                      (N114)? data_i[3361] : 
                      (N116)? data_i[3489] : 
                      (N118)? data_i[3617] : 
                      (N120)? data_i[3745] : 
                      (N122)? data_i[3873] : 
                      (N124)? data_i[4001] : 1'b0;
  assign data_o[32] = (N93)? data_i[32] : 
                      (N95)? data_i[160] : 
                      (N97)? data_i[288] : 
                      (N99)? data_i[416] : 
                      (N101)? data_i[544] : 
                      (N103)? data_i[672] : 
                      (N105)? data_i[800] : 
                      (N107)? data_i[928] : 
                      (N109)? data_i[1056] : 
                      (N111)? data_i[1184] : 
                      (N113)? data_i[1312] : 
                      (N115)? data_i[1440] : 
                      (N117)? data_i[1568] : 
                      (N119)? data_i[1696] : 
                      (N121)? data_i[1824] : 
                      (N123)? data_i[1952] : 
                      (N94)? data_i[2080] : 
                      (N96)? data_i[2208] : 
                      (N98)? data_i[2336] : 
                      (N100)? data_i[2464] : 
                      (N102)? data_i[2592] : 
                      (N104)? data_i[2720] : 
                      (N106)? data_i[2848] : 
                      (N108)? data_i[2976] : 
                      (N110)? data_i[3104] : 
                      (N112)? data_i[3232] : 
                      (N114)? data_i[3360] : 
                      (N116)? data_i[3488] : 
                      (N118)? data_i[3616] : 
                      (N120)? data_i[3744] : 
                      (N122)? data_i[3872] : 
                      (N124)? data_i[4000] : 1'b0;
  assign data_o[31] = (N93)? data_i[31] : 
                      (N95)? data_i[159] : 
                      (N97)? data_i[287] : 
                      (N99)? data_i[415] : 
                      (N101)? data_i[543] : 
                      (N103)? data_i[671] : 
                      (N105)? data_i[799] : 
                      (N107)? data_i[927] : 
                      (N109)? data_i[1055] : 
                      (N111)? data_i[1183] : 
                      (N113)? data_i[1311] : 
                      (N115)? data_i[1439] : 
                      (N117)? data_i[1567] : 
                      (N119)? data_i[1695] : 
                      (N121)? data_i[1823] : 
                      (N123)? data_i[1951] : 
                      (N94)? data_i[2079] : 
                      (N96)? data_i[2207] : 
                      (N98)? data_i[2335] : 
                      (N100)? data_i[2463] : 
                      (N102)? data_i[2591] : 
                      (N104)? data_i[2719] : 
                      (N106)? data_i[2847] : 
                      (N108)? data_i[2975] : 
                      (N110)? data_i[3103] : 
                      (N112)? data_i[3231] : 
                      (N114)? data_i[3359] : 
                      (N116)? data_i[3487] : 
                      (N118)? data_i[3615] : 
                      (N120)? data_i[3743] : 
                      (N122)? data_i[3871] : 
                      (N124)? data_i[3999] : 1'b0;
  assign data_o[30] = (N93)? data_i[30] : 
                      (N95)? data_i[158] : 
                      (N97)? data_i[286] : 
                      (N99)? data_i[414] : 
                      (N101)? data_i[542] : 
                      (N103)? data_i[670] : 
                      (N105)? data_i[798] : 
                      (N107)? data_i[926] : 
                      (N109)? data_i[1054] : 
                      (N111)? data_i[1182] : 
                      (N113)? data_i[1310] : 
                      (N115)? data_i[1438] : 
                      (N117)? data_i[1566] : 
                      (N119)? data_i[1694] : 
                      (N121)? data_i[1822] : 
                      (N123)? data_i[1950] : 
                      (N94)? data_i[2078] : 
                      (N96)? data_i[2206] : 
                      (N98)? data_i[2334] : 
                      (N100)? data_i[2462] : 
                      (N102)? data_i[2590] : 
                      (N104)? data_i[2718] : 
                      (N106)? data_i[2846] : 
                      (N108)? data_i[2974] : 
                      (N110)? data_i[3102] : 
                      (N112)? data_i[3230] : 
                      (N114)? data_i[3358] : 
                      (N116)? data_i[3486] : 
                      (N118)? data_i[3614] : 
                      (N120)? data_i[3742] : 
                      (N122)? data_i[3870] : 
                      (N124)? data_i[3998] : 1'b0;
  assign data_o[29] = (N93)? data_i[29] : 
                      (N95)? data_i[157] : 
                      (N97)? data_i[285] : 
                      (N99)? data_i[413] : 
                      (N101)? data_i[541] : 
                      (N103)? data_i[669] : 
                      (N105)? data_i[797] : 
                      (N107)? data_i[925] : 
                      (N109)? data_i[1053] : 
                      (N111)? data_i[1181] : 
                      (N113)? data_i[1309] : 
                      (N115)? data_i[1437] : 
                      (N117)? data_i[1565] : 
                      (N119)? data_i[1693] : 
                      (N121)? data_i[1821] : 
                      (N123)? data_i[1949] : 
                      (N94)? data_i[2077] : 
                      (N96)? data_i[2205] : 
                      (N98)? data_i[2333] : 
                      (N100)? data_i[2461] : 
                      (N102)? data_i[2589] : 
                      (N104)? data_i[2717] : 
                      (N106)? data_i[2845] : 
                      (N108)? data_i[2973] : 
                      (N110)? data_i[3101] : 
                      (N112)? data_i[3229] : 
                      (N114)? data_i[3357] : 
                      (N116)? data_i[3485] : 
                      (N118)? data_i[3613] : 
                      (N120)? data_i[3741] : 
                      (N122)? data_i[3869] : 
                      (N124)? data_i[3997] : 1'b0;
  assign data_o[28] = (N93)? data_i[28] : 
                      (N95)? data_i[156] : 
                      (N97)? data_i[284] : 
                      (N99)? data_i[412] : 
                      (N101)? data_i[540] : 
                      (N103)? data_i[668] : 
                      (N105)? data_i[796] : 
                      (N107)? data_i[924] : 
                      (N109)? data_i[1052] : 
                      (N111)? data_i[1180] : 
                      (N113)? data_i[1308] : 
                      (N115)? data_i[1436] : 
                      (N117)? data_i[1564] : 
                      (N119)? data_i[1692] : 
                      (N121)? data_i[1820] : 
                      (N123)? data_i[1948] : 
                      (N94)? data_i[2076] : 
                      (N96)? data_i[2204] : 
                      (N98)? data_i[2332] : 
                      (N100)? data_i[2460] : 
                      (N102)? data_i[2588] : 
                      (N104)? data_i[2716] : 
                      (N106)? data_i[2844] : 
                      (N108)? data_i[2972] : 
                      (N110)? data_i[3100] : 
                      (N112)? data_i[3228] : 
                      (N114)? data_i[3356] : 
                      (N116)? data_i[3484] : 
                      (N118)? data_i[3612] : 
                      (N120)? data_i[3740] : 
                      (N122)? data_i[3868] : 
                      (N124)? data_i[3996] : 1'b0;
  assign data_o[27] = (N93)? data_i[27] : 
                      (N95)? data_i[155] : 
                      (N97)? data_i[283] : 
                      (N99)? data_i[411] : 
                      (N101)? data_i[539] : 
                      (N103)? data_i[667] : 
                      (N105)? data_i[795] : 
                      (N107)? data_i[923] : 
                      (N109)? data_i[1051] : 
                      (N111)? data_i[1179] : 
                      (N113)? data_i[1307] : 
                      (N115)? data_i[1435] : 
                      (N117)? data_i[1563] : 
                      (N119)? data_i[1691] : 
                      (N121)? data_i[1819] : 
                      (N123)? data_i[1947] : 
                      (N94)? data_i[2075] : 
                      (N96)? data_i[2203] : 
                      (N98)? data_i[2331] : 
                      (N100)? data_i[2459] : 
                      (N102)? data_i[2587] : 
                      (N104)? data_i[2715] : 
                      (N106)? data_i[2843] : 
                      (N108)? data_i[2971] : 
                      (N110)? data_i[3099] : 
                      (N112)? data_i[3227] : 
                      (N114)? data_i[3355] : 
                      (N116)? data_i[3483] : 
                      (N118)? data_i[3611] : 
                      (N120)? data_i[3739] : 
                      (N122)? data_i[3867] : 
                      (N124)? data_i[3995] : 1'b0;
  assign data_o[26] = (N93)? data_i[26] : 
                      (N95)? data_i[154] : 
                      (N97)? data_i[282] : 
                      (N99)? data_i[410] : 
                      (N101)? data_i[538] : 
                      (N103)? data_i[666] : 
                      (N105)? data_i[794] : 
                      (N107)? data_i[922] : 
                      (N109)? data_i[1050] : 
                      (N111)? data_i[1178] : 
                      (N113)? data_i[1306] : 
                      (N115)? data_i[1434] : 
                      (N117)? data_i[1562] : 
                      (N119)? data_i[1690] : 
                      (N121)? data_i[1818] : 
                      (N123)? data_i[1946] : 
                      (N94)? data_i[2074] : 
                      (N96)? data_i[2202] : 
                      (N98)? data_i[2330] : 
                      (N100)? data_i[2458] : 
                      (N102)? data_i[2586] : 
                      (N104)? data_i[2714] : 
                      (N106)? data_i[2842] : 
                      (N108)? data_i[2970] : 
                      (N110)? data_i[3098] : 
                      (N112)? data_i[3226] : 
                      (N114)? data_i[3354] : 
                      (N116)? data_i[3482] : 
                      (N118)? data_i[3610] : 
                      (N120)? data_i[3738] : 
                      (N122)? data_i[3866] : 
                      (N124)? data_i[3994] : 1'b0;
  assign data_o[25] = (N93)? data_i[25] : 
                      (N95)? data_i[153] : 
                      (N97)? data_i[281] : 
                      (N99)? data_i[409] : 
                      (N101)? data_i[537] : 
                      (N103)? data_i[665] : 
                      (N105)? data_i[793] : 
                      (N107)? data_i[921] : 
                      (N109)? data_i[1049] : 
                      (N111)? data_i[1177] : 
                      (N113)? data_i[1305] : 
                      (N115)? data_i[1433] : 
                      (N117)? data_i[1561] : 
                      (N119)? data_i[1689] : 
                      (N121)? data_i[1817] : 
                      (N123)? data_i[1945] : 
                      (N94)? data_i[2073] : 
                      (N96)? data_i[2201] : 
                      (N98)? data_i[2329] : 
                      (N100)? data_i[2457] : 
                      (N102)? data_i[2585] : 
                      (N104)? data_i[2713] : 
                      (N106)? data_i[2841] : 
                      (N108)? data_i[2969] : 
                      (N110)? data_i[3097] : 
                      (N112)? data_i[3225] : 
                      (N114)? data_i[3353] : 
                      (N116)? data_i[3481] : 
                      (N118)? data_i[3609] : 
                      (N120)? data_i[3737] : 
                      (N122)? data_i[3865] : 
                      (N124)? data_i[3993] : 1'b0;
  assign data_o[24] = (N93)? data_i[24] : 
                      (N95)? data_i[152] : 
                      (N97)? data_i[280] : 
                      (N99)? data_i[408] : 
                      (N101)? data_i[536] : 
                      (N103)? data_i[664] : 
                      (N105)? data_i[792] : 
                      (N107)? data_i[920] : 
                      (N109)? data_i[1048] : 
                      (N111)? data_i[1176] : 
                      (N113)? data_i[1304] : 
                      (N115)? data_i[1432] : 
                      (N117)? data_i[1560] : 
                      (N119)? data_i[1688] : 
                      (N121)? data_i[1816] : 
                      (N123)? data_i[1944] : 
                      (N94)? data_i[2072] : 
                      (N96)? data_i[2200] : 
                      (N98)? data_i[2328] : 
                      (N100)? data_i[2456] : 
                      (N102)? data_i[2584] : 
                      (N104)? data_i[2712] : 
                      (N106)? data_i[2840] : 
                      (N108)? data_i[2968] : 
                      (N110)? data_i[3096] : 
                      (N112)? data_i[3224] : 
                      (N114)? data_i[3352] : 
                      (N116)? data_i[3480] : 
                      (N118)? data_i[3608] : 
                      (N120)? data_i[3736] : 
                      (N122)? data_i[3864] : 
                      (N124)? data_i[3992] : 1'b0;
  assign data_o[23] = (N93)? data_i[23] : 
                      (N95)? data_i[151] : 
                      (N97)? data_i[279] : 
                      (N99)? data_i[407] : 
                      (N101)? data_i[535] : 
                      (N103)? data_i[663] : 
                      (N105)? data_i[791] : 
                      (N107)? data_i[919] : 
                      (N109)? data_i[1047] : 
                      (N111)? data_i[1175] : 
                      (N113)? data_i[1303] : 
                      (N115)? data_i[1431] : 
                      (N117)? data_i[1559] : 
                      (N119)? data_i[1687] : 
                      (N121)? data_i[1815] : 
                      (N123)? data_i[1943] : 
                      (N94)? data_i[2071] : 
                      (N96)? data_i[2199] : 
                      (N98)? data_i[2327] : 
                      (N100)? data_i[2455] : 
                      (N102)? data_i[2583] : 
                      (N104)? data_i[2711] : 
                      (N106)? data_i[2839] : 
                      (N108)? data_i[2967] : 
                      (N110)? data_i[3095] : 
                      (N112)? data_i[3223] : 
                      (N114)? data_i[3351] : 
                      (N116)? data_i[3479] : 
                      (N118)? data_i[3607] : 
                      (N120)? data_i[3735] : 
                      (N122)? data_i[3863] : 
                      (N124)? data_i[3991] : 1'b0;
  assign data_o[22] = (N93)? data_i[22] : 
                      (N95)? data_i[150] : 
                      (N97)? data_i[278] : 
                      (N99)? data_i[406] : 
                      (N101)? data_i[534] : 
                      (N103)? data_i[662] : 
                      (N105)? data_i[790] : 
                      (N107)? data_i[918] : 
                      (N109)? data_i[1046] : 
                      (N111)? data_i[1174] : 
                      (N113)? data_i[1302] : 
                      (N115)? data_i[1430] : 
                      (N117)? data_i[1558] : 
                      (N119)? data_i[1686] : 
                      (N121)? data_i[1814] : 
                      (N123)? data_i[1942] : 
                      (N94)? data_i[2070] : 
                      (N96)? data_i[2198] : 
                      (N98)? data_i[2326] : 
                      (N100)? data_i[2454] : 
                      (N102)? data_i[2582] : 
                      (N104)? data_i[2710] : 
                      (N106)? data_i[2838] : 
                      (N108)? data_i[2966] : 
                      (N110)? data_i[3094] : 
                      (N112)? data_i[3222] : 
                      (N114)? data_i[3350] : 
                      (N116)? data_i[3478] : 
                      (N118)? data_i[3606] : 
                      (N120)? data_i[3734] : 
                      (N122)? data_i[3862] : 
                      (N124)? data_i[3990] : 1'b0;
  assign data_o[21] = (N93)? data_i[21] : 
                      (N95)? data_i[149] : 
                      (N97)? data_i[277] : 
                      (N99)? data_i[405] : 
                      (N101)? data_i[533] : 
                      (N103)? data_i[661] : 
                      (N105)? data_i[789] : 
                      (N107)? data_i[917] : 
                      (N109)? data_i[1045] : 
                      (N111)? data_i[1173] : 
                      (N113)? data_i[1301] : 
                      (N115)? data_i[1429] : 
                      (N117)? data_i[1557] : 
                      (N119)? data_i[1685] : 
                      (N121)? data_i[1813] : 
                      (N123)? data_i[1941] : 
                      (N94)? data_i[2069] : 
                      (N96)? data_i[2197] : 
                      (N98)? data_i[2325] : 
                      (N100)? data_i[2453] : 
                      (N102)? data_i[2581] : 
                      (N104)? data_i[2709] : 
                      (N106)? data_i[2837] : 
                      (N108)? data_i[2965] : 
                      (N110)? data_i[3093] : 
                      (N112)? data_i[3221] : 
                      (N114)? data_i[3349] : 
                      (N116)? data_i[3477] : 
                      (N118)? data_i[3605] : 
                      (N120)? data_i[3733] : 
                      (N122)? data_i[3861] : 
                      (N124)? data_i[3989] : 1'b0;
  assign data_o[20] = (N93)? data_i[20] : 
                      (N95)? data_i[148] : 
                      (N97)? data_i[276] : 
                      (N99)? data_i[404] : 
                      (N101)? data_i[532] : 
                      (N103)? data_i[660] : 
                      (N105)? data_i[788] : 
                      (N107)? data_i[916] : 
                      (N109)? data_i[1044] : 
                      (N111)? data_i[1172] : 
                      (N113)? data_i[1300] : 
                      (N115)? data_i[1428] : 
                      (N117)? data_i[1556] : 
                      (N119)? data_i[1684] : 
                      (N121)? data_i[1812] : 
                      (N123)? data_i[1940] : 
                      (N94)? data_i[2068] : 
                      (N96)? data_i[2196] : 
                      (N98)? data_i[2324] : 
                      (N100)? data_i[2452] : 
                      (N102)? data_i[2580] : 
                      (N104)? data_i[2708] : 
                      (N106)? data_i[2836] : 
                      (N108)? data_i[2964] : 
                      (N110)? data_i[3092] : 
                      (N112)? data_i[3220] : 
                      (N114)? data_i[3348] : 
                      (N116)? data_i[3476] : 
                      (N118)? data_i[3604] : 
                      (N120)? data_i[3732] : 
                      (N122)? data_i[3860] : 
                      (N124)? data_i[3988] : 1'b0;
  assign data_o[19] = (N93)? data_i[19] : 
                      (N95)? data_i[147] : 
                      (N97)? data_i[275] : 
                      (N99)? data_i[403] : 
                      (N101)? data_i[531] : 
                      (N103)? data_i[659] : 
                      (N105)? data_i[787] : 
                      (N107)? data_i[915] : 
                      (N109)? data_i[1043] : 
                      (N111)? data_i[1171] : 
                      (N113)? data_i[1299] : 
                      (N115)? data_i[1427] : 
                      (N117)? data_i[1555] : 
                      (N119)? data_i[1683] : 
                      (N121)? data_i[1811] : 
                      (N123)? data_i[1939] : 
                      (N94)? data_i[2067] : 
                      (N96)? data_i[2195] : 
                      (N98)? data_i[2323] : 
                      (N100)? data_i[2451] : 
                      (N102)? data_i[2579] : 
                      (N104)? data_i[2707] : 
                      (N106)? data_i[2835] : 
                      (N108)? data_i[2963] : 
                      (N110)? data_i[3091] : 
                      (N112)? data_i[3219] : 
                      (N114)? data_i[3347] : 
                      (N116)? data_i[3475] : 
                      (N118)? data_i[3603] : 
                      (N120)? data_i[3731] : 
                      (N122)? data_i[3859] : 
                      (N124)? data_i[3987] : 1'b0;
  assign data_o[18] = (N93)? data_i[18] : 
                      (N95)? data_i[146] : 
                      (N97)? data_i[274] : 
                      (N99)? data_i[402] : 
                      (N101)? data_i[530] : 
                      (N103)? data_i[658] : 
                      (N105)? data_i[786] : 
                      (N107)? data_i[914] : 
                      (N109)? data_i[1042] : 
                      (N111)? data_i[1170] : 
                      (N113)? data_i[1298] : 
                      (N115)? data_i[1426] : 
                      (N117)? data_i[1554] : 
                      (N119)? data_i[1682] : 
                      (N121)? data_i[1810] : 
                      (N123)? data_i[1938] : 
                      (N94)? data_i[2066] : 
                      (N96)? data_i[2194] : 
                      (N98)? data_i[2322] : 
                      (N100)? data_i[2450] : 
                      (N102)? data_i[2578] : 
                      (N104)? data_i[2706] : 
                      (N106)? data_i[2834] : 
                      (N108)? data_i[2962] : 
                      (N110)? data_i[3090] : 
                      (N112)? data_i[3218] : 
                      (N114)? data_i[3346] : 
                      (N116)? data_i[3474] : 
                      (N118)? data_i[3602] : 
                      (N120)? data_i[3730] : 
                      (N122)? data_i[3858] : 
                      (N124)? data_i[3986] : 1'b0;
  assign data_o[17] = (N93)? data_i[17] : 
                      (N95)? data_i[145] : 
                      (N97)? data_i[273] : 
                      (N99)? data_i[401] : 
                      (N101)? data_i[529] : 
                      (N103)? data_i[657] : 
                      (N105)? data_i[785] : 
                      (N107)? data_i[913] : 
                      (N109)? data_i[1041] : 
                      (N111)? data_i[1169] : 
                      (N113)? data_i[1297] : 
                      (N115)? data_i[1425] : 
                      (N117)? data_i[1553] : 
                      (N119)? data_i[1681] : 
                      (N121)? data_i[1809] : 
                      (N123)? data_i[1937] : 
                      (N94)? data_i[2065] : 
                      (N96)? data_i[2193] : 
                      (N98)? data_i[2321] : 
                      (N100)? data_i[2449] : 
                      (N102)? data_i[2577] : 
                      (N104)? data_i[2705] : 
                      (N106)? data_i[2833] : 
                      (N108)? data_i[2961] : 
                      (N110)? data_i[3089] : 
                      (N112)? data_i[3217] : 
                      (N114)? data_i[3345] : 
                      (N116)? data_i[3473] : 
                      (N118)? data_i[3601] : 
                      (N120)? data_i[3729] : 
                      (N122)? data_i[3857] : 
                      (N124)? data_i[3985] : 1'b0;
  assign data_o[16] = (N93)? data_i[16] : 
                      (N95)? data_i[144] : 
                      (N97)? data_i[272] : 
                      (N99)? data_i[400] : 
                      (N101)? data_i[528] : 
                      (N103)? data_i[656] : 
                      (N105)? data_i[784] : 
                      (N107)? data_i[912] : 
                      (N109)? data_i[1040] : 
                      (N111)? data_i[1168] : 
                      (N113)? data_i[1296] : 
                      (N115)? data_i[1424] : 
                      (N117)? data_i[1552] : 
                      (N119)? data_i[1680] : 
                      (N121)? data_i[1808] : 
                      (N123)? data_i[1936] : 
                      (N94)? data_i[2064] : 
                      (N96)? data_i[2192] : 
                      (N98)? data_i[2320] : 
                      (N100)? data_i[2448] : 
                      (N102)? data_i[2576] : 
                      (N104)? data_i[2704] : 
                      (N106)? data_i[2832] : 
                      (N108)? data_i[2960] : 
                      (N110)? data_i[3088] : 
                      (N112)? data_i[3216] : 
                      (N114)? data_i[3344] : 
                      (N116)? data_i[3472] : 
                      (N118)? data_i[3600] : 
                      (N120)? data_i[3728] : 
                      (N122)? data_i[3856] : 
                      (N124)? data_i[3984] : 1'b0;
  assign data_o[15] = (N93)? data_i[15] : 
                      (N95)? data_i[143] : 
                      (N97)? data_i[271] : 
                      (N99)? data_i[399] : 
                      (N101)? data_i[527] : 
                      (N103)? data_i[655] : 
                      (N105)? data_i[783] : 
                      (N107)? data_i[911] : 
                      (N109)? data_i[1039] : 
                      (N111)? data_i[1167] : 
                      (N113)? data_i[1295] : 
                      (N115)? data_i[1423] : 
                      (N117)? data_i[1551] : 
                      (N119)? data_i[1679] : 
                      (N121)? data_i[1807] : 
                      (N123)? data_i[1935] : 
                      (N94)? data_i[2063] : 
                      (N96)? data_i[2191] : 
                      (N98)? data_i[2319] : 
                      (N100)? data_i[2447] : 
                      (N102)? data_i[2575] : 
                      (N104)? data_i[2703] : 
                      (N106)? data_i[2831] : 
                      (N108)? data_i[2959] : 
                      (N110)? data_i[3087] : 
                      (N112)? data_i[3215] : 
                      (N114)? data_i[3343] : 
                      (N116)? data_i[3471] : 
                      (N118)? data_i[3599] : 
                      (N120)? data_i[3727] : 
                      (N122)? data_i[3855] : 
                      (N124)? data_i[3983] : 1'b0;
  assign data_o[14] = (N93)? data_i[14] : 
                      (N95)? data_i[142] : 
                      (N97)? data_i[270] : 
                      (N99)? data_i[398] : 
                      (N101)? data_i[526] : 
                      (N103)? data_i[654] : 
                      (N105)? data_i[782] : 
                      (N107)? data_i[910] : 
                      (N109)? data_i[1038] : 
                      (N111)? data_i[1166] : 
                      (N113)? data_i[1294] : 
                      (N115)? data_i[1422] : 
                      (N117)? data_i[1550] : 
                      (N119)? data_i[1678] : 
                      (N121)? data_i[1806] : 
                      (N123)? data_i[1934] : 
                      (N94)? data_i[2062] : 
                      (N96)? data_i[2190] : 
                      (N98)? data_i[2318] : 
                      (N100)? data_i[2446] : 
                      (N102)? data_i[2574] : 
                      (N104)? data_i[2702] : 
                      (N106)? data_i[2830] : 
                      (N108)? data_i[2958] : 
                      (N110)? data_i[3086] : 
                      (N112)? data_i[3214] : 
                      (N114)? data_i[3342] : 
                      (N116)? data_i[3470] : 
                      (N118)? data_i[3598] : 
                      (N120)? data_i[3726] : 
                      (N122)? data_i[3854] : 
                      (N124)? data_i[3982] : 1'b0;
  assign data_o[13] = (N93)? data_i[13] : 
                      (N95)? data_i[141] : 
                      (N97)? data_i[269] : 
                      (N99)? data_i[397] : 
                      (N101)? data_i[525] : 
                      (N103)? data_i[653] : 
                      (N105)? data_i[781] : 
                      (N107)? data_i[909] : 
                      (N109)? data_i[1037] : 
                      (N111)? data_i[1165] : 
                      (N113)? data_i[1293] : 
                      (N115)? data_i[1421] : 
                      (N117)? data_i[1549] : 
                      (N119)? data_i[1677] : 
                      (N121)? data_i[1805] : 
                      (N123)? data_i[1933] : 
                      (N94)? data_i[2061] : 
                      (N96)? data_i[2189] : 
                      (N98)? data_i[2317] : 
                      (N100)? data_i[2445] : 
                      (N102)? data_i[2573] : 
                      (N104)? data_i[2701] : 
                      (N106)? data_i[2829] : 
                      (N108)? data_i[2957] : 
                      (N110)? data_i[3085] : 
                      (N112)? data_i[3213] : 
                      (N114)? data_i[3341] : 
                      (N116)? data_i[3469] : 
                      (N118)? data_i[3597] : 
                      (N120)? data_i[3725] : 
                      (N122)? data_i[3853] : 
                      (N124)? data_i[3981] : 1'b0;
  assign data_o[12] = (N93)? data_i[12] : 
                      (N95)? data_i[140] : 
                      (N97)? data_i[268] : 
                      (N99)? data_i[396] : 
                      (N101)? data_i[524] : 
                      (N103)? data_i[652] : 
                      (N105)? data_i[780] : 
                      (N107)? data_i[908] : 
                      (N109)? data_i[1036] : 
                      (N111)? data_i[1164] : 
                      (N113)? data_i[1292] : 
                      (N115)? data_i[1420] : 
                      (N117)? data_i[1548] : 
                      (N119)? data_i[1676] : 
                      (N121)? data_i[1804] : 
                      (N123)? data_i[1932] : 
                      (N94)? data_i[2060] : 
                      (N96)? data_i[2188] : 
                      (N98)? data_i[2316] : 
                      (N100)? data_i[2444] : 
                      (N102)? data_i[2572] : 
                      (N104)? data_i[2700] : 
                      (N106)? data_i[2828] : 
                      (N108)? data_i[2956] : 
                      (N110)? data_i[3084] : 
                      (N112)? data_i[3212] : 
                      (N114)? data_i[3340] : 
                      (N116)? data_i[3468] : 
                      (N118)? data_i[3596] : 
                      (N120)? data_i[3724] : 
                      (N122)? data_i[3852] : 
                      (N124)? data_i[3980] : 1'b0;
  assign data_o[11] = (N93)? data_i[11] : 
                      (N95)? data_i[139] : 
                      (N97)? data_i[267] : 
                      (N99)? data_i[395] : 
                      (N101)? data_i[523] : 
                      (N103)? data_i[651] : 
                      (N105)? data_i[779] : 
                      (N107)? data_i[907] : 
                      (N109)? data_i[1035] : 
                      (N111)? data_i[1163] : 
                      (N113)? data_i[1291] : 
                      (N115)? data_i[1419] : 
                      (N117)? data_i[1547] : 
                      (N119)? data_i[1675] : 
                      (N121)? data_i[1803] : 
                      (N123)? data_i[1931] : 
                      (N94)? data_i[2059] : 
                      (N96)? data_i[2187] : 
                      (N98)? data_i[2315] : 
                      (N100)? data_i[2443] : 
                      (N102)? data_i[2571] : 
                      (N104)? data_i[2699] : 
                      (N106)? data_i[2827] : 
                      (N108)? data_i[2955] : 
                      (N110)? data_i[3083] : 
                      (N112)? data_i[3211] : 
                      (N114)? data_i[3339] : 
                      (N116)? data_i[3467] : 
                      (N118)? data_i[3595] : 
                      (N120)? data_i[3723] : 
                      (N122)? data_i[3851] : 
                      (N124)? data_i[3979] : 1'b0;
  assign data_o[10] = (N93)? data_i[10] : 
                      (N95)? data_i[138] : 
                      (N97)? data_i[266] : 
                      (N99)? data_i[394] : 
                      (N101)? data_i[522] : 
                      (N103)? data_i[650] : 
                      (N105)? data_i[778] : 
                      (N107)? data_i[906] : 
                      (N109)? data_i[1034] : 
                      (N111)? data_i[1162] : 
                      (N113)? data_i[1290] : 
                      (N115)? data_i[1418] : 
                      (N117)? data_i[1546] : 
                      (N119)? data_i[1674] : 
                      (N121)? data_i[1802] : 
                      (N123)? data_i[1930] : 
                      (N94)? data_i[2058] : 
                      (N96)? data_i[2186] : 
                      (N98)? data_i[2314] : 
                      (N100)? data_i[2442] : 
                      (N102)? data_i[2570] : 
                      (N104)? data_i[2698] : 
                      (N106)? data_i[2826] : 
                      (N108)? data_i[2954] : 
                      (N110)? data_i[3082] : 
                      (N112)? data_i[3210] : 
                      (N114)? data_i[3338] : 
                      (N116)? data_i[3466] : 
                      (N118)? data_i[3594] : 
                      (N120)? data_i[3722] : 
                      (N122)? data_i[3850] : 
                      (N124)? data_i[3978] : 1'b0;
  assign data_o[9] = (N93)? data_i[9] : 
                     (N95)? data_i[137] : 
                     (N97)? data_i[265] : 
                     (N99)? data_i[393] : 
                     (N101)? data_i[521] : 
                     (N103)? data_i[649] : 
                     (N105)? data_i[777] : 
                     (N107)? data_i[905] : 
                     (N109)? data_i[1033] : 
                     (N111)? data_i[1161] : 
                     (N113)? data_i[1289] : 
                     (N115)? data_i[1417] : 
                     (N117)? data_i[1545] : 
                     (N119)? data_i[1673] : 
                     (N121)? data_i[1801] : 
                     (N123)? data_i[1929] : 
                     (N94)? data_i[2057] : 
                     (N96)? data_i[2185] : 
                     (N98)? data_i[2313] : 
                     (N100)? data_i[2441] : 
                     (N102)? data_i[2569] : 
                     (N104)? data_i[2697] : 
                     (N106)? data_i[2825] : 
                     (N108)? data_i[2953] : 
                     (N110)? data_i[3081] : 
                     (N112)? data_i[3209] : 
                     (N114)? data_i[3337] : 
                     (N116)? data_i[3465] : 
                     (N118)? data_i[3593] : 
                     (N120)? data_i[3721] : 
                     (N122)? data_i[3849] : 
                     (N124)? data_i[3977] : 1'b0;
  assign data_o[8] = (N93)? data_i[8] : 
                     (N95)? data_i[136] : 
                     (N97)? data_i[264] : 
                     (N99)? data_i[392] : 
                     (N101)? data_i[520] : 
                     (N103)? data_i[648] : 
                     (N105)? data_i[776] : 
                     (N107)? data_i[904] : 
                     (N109)? data_i[1032] : 
                     (N111)? data_i[1160] : 
                     (N113)? data_i[1288] : 
                     (N115)? data_i[1416] : 
                     (N117)? data_i[1544] : 
                     (N119)? data_i[1672] : 
                     (N121)? data_i[1800] : 
                     (N123)? data_i[1928] : 
                     (N94)? data_i[2056] : 
                     (N96)? data_i[2184] : 
                     (N98)? data_i[2312] : 
                     (N100)? data_i[2440] : 
                     (N102)? data_i[2568] : 
                     (N104)? data_i[2696] : 
                     (N106)? data_i[2824] : 
                     (N108)? data_i[2952] : 
                     (N110)? data_i[3080] : 
                     (N112)? data_i[3208] : 
                     (N114)? data_i[3336] : 
                     (N116)? data_i[3464] : 
                     (N118)? data_i[3592] : 
                     (N120)? data_i[3720] : 
                     (N122)? data_i[3848] : 
                     (N124)? data_i[3976] : 1'b0;
  assign data_o[7] = (N93)? data_i[7] : 
                     (N95)? data_i[135] : 
                     (N97)? data_i[263] : 
                     (N99)? data_i[391] : 
                     (N101)? data_i[519] : 
                     (N103)? data_i[647] : 
                     (N105)? data_i[775] : 
                     (N107)? data_i[903] : 
                     (N109)? data_i[1031] : 
                     (N111)? data_i[1159] : 
                     (N113)? data_i[1287] : 
                     (N115)? data_i[1415] : 
                     (N117)? data_i[1543] : 
                     (N119)? data_i[1671] : 
                     (N121)? data_i[1799] : 
                     (N123)? data_i[1927] : 
                     (N94)? data_i[2055] : 
                     (N96)? data_i[2183] : 
                     (N98)? data_i[2311] : 
                     (N100)? data_i[2439] : 
                     (N102)? data_i[2567] : 
                     (N104)? data_i[2695] : 
                     (N106)? data_i[2823] : 
                     (N108)? data_i[2951] : 
                     (N110)? data_i[3079] : 
                     (N112)? data_i[3207] : 
                     (N114)? data_i[3335] : 
                     (N116)? data_i[3463] : 
                     (N118)? data_i[3591] : 
                     (N120)? data_i[3719] : 
                     (N122)? data_i[3847] : 
                     (N124)? data_i[3975] : 1'b0;
  assign data_o[6] = (N93)? data_i[6] : 
                     (N95)? data_i[134] : 
                     (N97)? data_i[262] : 
                     (N99)? data_i[390] : 
                     (N101)? data_i[518] : 
                     (N103)? data_i[646] : 
                     (N105)? data_i[774] : 
                     (N107)? data_i[902] : 
                     (N109)? data_i[1030] : 
                     (N111)? data_i[1158] : 
                     (N113)? data_i[1286] : 
                     (N115)? data_i[1414] : 
                     (N117)? data_i[1542] : 
                     (N119)? data_i[1670] : 
                     (N121)? data_i[1798] : 
                     (N123)? data_i[1926] : 
                     (N94)? data_i[2054] : 
                     (N96)? data_i[2182] : 
                     (N98)? data_i[2310] : 
                     (N100)? data_i[2438] : 
                     (N102)? data_i[2566] : 
                     (N104)? data_i[2694] : 
                     (N106)? data_i[2822] : 
                     (N108)? data_i[2950] : 
                     (N110)? data_i[3078] : 
                     (N112)? data_i[3206] : 
                     (N114)? data_i[3334] : 
                     (N116)? data_i[3462] : 
                     (N118)? data_i[3590] : 
                     (N120)? data_i[3718] : 
                     (N122)? data_i[3846] : 
                     (N124)? data_i[3974] : 1'b0;
  assign data_o[5] = (N93)? data_i[5] : 
                     (N95)? data_i[133] : 
                     (N97)? data_i[261] : 
                     (N99)? data_i[389] : 
                     (N101)? data_i[517] : 
                     (N103)? data_i[645] : 
                     (N105)? data_i[773] : 
                     (N107)? data_i[901] : 
                     (N109)? data_i[1029] : 
                     (N111)? data_i[1157] : 
                     (N113)? data_i[1285] : 
                     (N115)? data_i[1413] : 
                     (N117)? data_i[1541] : 
                     (N119)? data_i[1669] : 
                     (N121)? data_i[1797] : 
                     (N123)? data_i[1925] : 
                     (N94)? data_i[2053] : 
                     (N96)? data_i[2181] : 
                     (N98)? data_i[2309] : 
                     (N100)? data_i[2437] : 
                     (N102)? data_i[2565] : 
                     (N104)? data_i[2693] : 
                     (N106)? data_i[2821] : 
                     (N108)? data_i[2949] : 
                     (N110)? data_i[3077] : 
                     (N112)? data_i[3205] : 
                     (N114)? data_i[3333] : 
                     (N116)? data_i[3461] : 
                     (N118)? data_i[3589] : 
                     (N120)? data_i[3717] : 
                     (N122)? data_i[3845] : 
                     (N124)? data_i[3973] : 1'b0;
  assign data_o[4] = (N93)? data_i[4] : 
                     (N95)? data_i[132] : 
                     (N97)? data_i[260] : 
                     (N99)? data_i[388] : 
                     (N101)? data_i[516] : 
                     (N103)? data_i[644] : 
                     (N105)? data_i[772] : 
                     (N107)? data_i[900] : 
                     (N109)? data_i[1028] : 
                     (N111)? data_i[1156] : 
                     (N113)? data_i[1284] : 
                     (N115)? data_i[1412] : 
                     (N117)? data_i[1540] : 
                     (N119)? data_i[1668] : 
                     (N121)? data_i[1796] : 
                     (N123)? data_i[1924] : 
                     (N94)? data_i[2052] : 
                     (N96)? data_i[2180] : 
                     (N98)? data_i[2308] : 
                     (N100)? data_i[2436] : 
                     (N102)? data_i[2564] : 
                     (N104)? data_i[2692] : 
                     (N106)? data_i[2820] : 
                     (N108)? data_i[2948] : 
                     (N110)? data_i[3076] : 
                     (N112)? data_i[3204] : 
                     (N114)? data_i[3332] : 
                     (N116)? data_i[3460] : 
                     (N118)? data_i[3588] : 
                     (N120)? data_i[3716] : 
                     (N122)? data_i[3844] : 
                     (N124)? data_i[3972] : 1'b0;
  assign data_o[3] = (N93)? data_i[3] : 
                     (N95)? data_i[131] : 
                     (N97)? data_i[259] : 
                     (N99)? data_i[387] : 
                     (N101)? data_i[515] : 
                     (N103)? data_i[643] : 
                     (N105)? data_i[771] : 
                     (N107)? data_i[899] : 
                     (N109)? data_i[1027] : 
                     (N111)? data_i[1155] : 
                     (N113)? data_i[1283] : 
                     (N115)? data_i[1411] : 
                     (N117)? data_i[1539] : 
                     (N119)? data_i[1667] : 
                     (N121)? data_i[1795] : 
                     (N123)? data_i[1923] : 
                     (N94)? data_i[2051] : 
                     (N96)? data_i[2179] : 
                     (N98)? data_i[2307] : 
                     (N100)? data_i[2435] : 
                     (N102)? data_i[2563] : 
                     (N104)? data_i[2691] : 
                     (N106)? data_i[2819] : 
                     (N108)? data_i[2947] : 
                     (N110)? data_i[3075] : 
                     (N112)? data_i[3203] : 
                     (N114)? data_i[3331] : 
                     (N116)? data_i[3459] : 
                     (N118)? data_i[3587] : 
                     (N120)? data_i[3715] : 
                     (N122)? data_i[3843] : 
                     (N124)? data_i[3971] : 1'b0;
  assign data_o[2] = (N93)? data_i[2] : 
                     (N95)? data_i[130] : 
                     (N97)? data_i[258] : 
                     (N99)? data_i[386] : 
                     (N101)? data_i[514] : 
                     (N103)? data_i[642] : 
                     (N105)? data_i[770] : 
                     (N107)? data_i[898] : 
                     (N109)? data_i[1026] : 
                     (N111)? data_i[1154] : 
                     (N113)? data_i[1282] : 
                     (N115)? data_i[1410] : 
                     (N117)? data_i[1538] : 
                     (N119)? data_i[1666] : 
                     (N121)? data_i[1794] : 
                     (N123)? data_i[1922] : 
                     (N94)? data_i[2050] : 
                     (N96)? data_i[2178] : 
                     (N98)? data_i[2306] : 
                     (N100)? data_i[2434] : 
                     (N102)? data_i[2562] : 
                     (N104)? data_i[2690] : 
                     (N106)? data_i[2818] : 
                     (N108)? data_i[2946] : 
                     (N110)? data_i[3074] : 
                     (N112)? data_i[3202] : 
                     (N114)? data_i[3330] : 
                     (N116)? data_i[3458] : 
                     (N118)? data_i[3586] : 
                     (N120)? data_i[3714] : 
                     (N122)? data_i[3842] : 
                     (N124)? data_i[3970] : 1'b0;
  assign data_o[1] = (N93)? data_i[1] : 
                     (N95)? data_i[129] : 
                     (N97)? data_i[257] : 
                     (N99)? data_i[385] : 
                     (N101)? data_i[513] : 
                     (N103)? data_i[641] : 
                     (N105)? data_i[769] : 
                     (N107)? data_i[897] : 
                     (N109)? data_i[1025] : 
                     (N111)? data_i[1153] : 
                     (N113)? data_i[1281] : 
                     (N115)? data_i[1409] : 
                     (N117)? data_i[1537] : 
                     (N119)? data_i[1665] : 
                     (N121)? data_i[1793] : 
                     (N123)? data_i[1921] : 
                     (N94)? data_i[2049] : 
                     (N96)? data_i[2177] : 
                     (N98)? data_i[2305] : 
                     (N100)? data_i[2433] : 
                     (N102)? data_i[2561] : 
                     (N104)? data_i[2689] : 
                     (N106)? data_i[2817] : 
                     (N108)? data_i[2945] : 
                     (N110)? data_i[3073] : 
                     (N112)? data_i[3201] : 
                     (N114)? data_i[3329] : 
                     (N116)? data_i[3457] : 
                     (N118)? data_i[3585] : 
                     (N120)? data_i[3713] : 
                     (N122)? data_i[3841] : 
                     (N124)? data_i[3969] : 1'b0;
  assign data_o[0] = (N93)? data_i[0] : 
                     (N95)? data_i[128] : 
                     (N97)? data_i[256] : 
                     (N99)? data_i[384] : 
                     (N101)? data_i[512] : 
                     (N103)? data_i[640] : 
                     (N105)? data_i[768] : 
                     (N107)? data_i[896] : 
                     (N109)? data_i[1024] : 
                     (N111)? data_i[1152] : 
                     (N113)? data_i[1280] : 
                     (N115)? data_i[1408] : 
                     (N117)? data_i[1536] : 
                     (N119)? data_i[1664] : 
                     (N121)? data_i[1792] : 
                     (N123)? data_i[1920] : 
                     (N94)? data_i[2048] : 
                     (N96)? data_i[2176] : 
                     (N98)? data_i[2304] : 
                     (N100)? data_i[2432] : 
                     (N102)? data_i[2560] : 
                     (N104)? data_i[2688] : 
                     (N106)? data_i[2816] : 
                     (N108)? data_i[2944] : 
                     (N110)? data_i[3072] : 
                     (N112)? data_i[3200] : 
                     (N114)? data_i[3328] : 
                     (N116)? data_i[3456] : 
                     (N118)? data_i[3584] : 
                     (N120)? data_i[3712] : 
                     (N122)? data_i[3840] : 
                     (N124)? data_i[3968] : 1'b0;
  assign yumi_o = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, yumi_i } << tag_o;
  assign N0 = ~tag_o[0];
  assign N1 = ~tag_o[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & tag_o[1];
  assign N4 = tag_o[0] & N1;
  assign N5 = tag_o[0] & tag_o[1];
  assign N6 = ~tag_o[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & tag_o[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & tag_o[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & tag_o[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & tag_o[2];
  assign N15 = ~tag_o[3];
  assign N16 = N7 & N15;
  assign N17 = N7 & tag_o[3];
  assign N18 = N9 & N15;
  assign N19 = N9 & tag_o[3];
  assign N20 = N11 & N15;
  assign N21 = N11 & tag_o[3];
  assign N22 = N13 & N15;
  assign N23 = N13 & tag_o[3];
  assign N24 = N8 & N15;
  assign N25 = N8 & tag_o[3];
  assign N26 = N10 & N15;
  assign N27 = N10 & tag_o[3];
  assign N28 = N12 & N15;
  assign N29 = N12 & tag_o[3];
  assign N30 = N14 & N15;
  assign N31 = N14 & tag_o[3];
  assign N32 = ~tag_o[4];
  assign N33 = N16 & N32;
  assign N34 = N16 & tag_o[4];
  assign N35 = N18 & N32;
  assign N36 = N18 & tag_o[4];
  assign N37 = N20 & N32;
  assign N38 = N20 & tag_o[4];
  assign N39 = N22 & N32;
  assign N40 = N22 & tag_o[4];
  assign N41 = N24 & N32;
  assign N42 = N24 & tag_o[4];
  assign N43 = N26 & N32;
  assign N44 = N26 & tag_o[4];
  assign N45 = N28 & N32;
  assign N46 = N28 & tag_o[4];
  assign N47 = N30 & N32;
  assign N48 = N30 & tag_o[4];
  assign N49 = N17 & N32;
  assign N50 = N17 & tag_o[4];
  assign N51 = N19 & N32;
  assign N52 = N19 & tag_o[4];
  assign N53 = N21 & N32;
  assign N54 = N21 & tag_o[4];
  assign N55 = N23 & N32;
  assign N56 = N23 & tag_o[4];
  assign N57 = N25 & N32;
  assign N58 = N25 & tag_o[4];
  assign N59 = N27 & N32;
  assign N60 = N27 & tag_o[4];
  assign N61 = N29 & N32;
  assign N62 = N29 & tag_o[4];
  assign N63 = N31 & N32;
  assign N64 = N31 & tag_o[4];
  assign N65 = N0 & N1;
  assign N66 = N0 & tag_o[1];
  assign N67 = tag_o[0] & N1;
  assign N68 = tag_o[0] & tag_o[1];
  assign N69 = N65 & N6;
  assign N70 = N65 & tag_o[2];
  assign N71 = N67 & N6;
  assign N72 = N67 & tag_o[2];
  assign N73 = N66 & N6;
  assign N74 = N66 & tag_o[2];
  assign N75 = N68 & N6;
  assign N76 = N68 & tag_o[2];
  assign N77 = N69 & N15;
  assign N78 = N69 & tag_o[3];
  assign N79 = N71 & N15;
  assign N80 = N71 & tag_o[3];
  assign N81 = N73 & N15;
  assign N82 = N73 & tag_o[3];
  assign N83 = N75 & N15;
  assign N84 = N75 & tag_o[3];
  assign N85 = N70 & N15;
  assign N86 = N70 & tag_o[3];
  assign N87 = N72 & N15;
  assign N88 = N72 & tag_o[3];
  assign N89 = N74 & N15;
  assign N90 = N74 & tag_o[3];
  assign N91 = N76 & N15;
  assign N92 = N76 & tag_o[3];
  assign N93 = N77 & N32;
  assign N94 = N77 & tag_o[4];
  assign N95 = N79 & N32;
  assign N96 = N79 & tag_o[4];
  assign N97 = N81 & N32;
  assign N98 = N81 & tag_o[4];
  assign N99 = N83 & N32;
  assign N100 = N83 & tag_o[4];
  assign N101 = N85 & N32;
  assign N102 = N85 & tag_o[4];
  assign N103 = N87 & N32;
  assign N104 = N87 & tag_o[4];
  assign N105 = N89 & N32;
  assign N106 = N89 & tag_o[4];
  assign N107 = N91 & N32;
  assign N108 = N91 & tag_o[4];
  assign N109 = N78 & N32;
  assign N110 = N78 & tag_o[4];
  assign N111 = N80 & N32;
  assign N112 = N80 & tag_o[4];
  assign N113 = N82 & N32;
  assign N114 = N82 & tag_o[4];
  assign N115 = N84 & N32;
  assign N116 = N84 & tag_o[4];
  assign N117 = N86 & N32;
  assign N118 = N86 & tag_o[4];
  assign N119 = N88 & N32;
  assign N120 = N88 & tag_o[4];
  assign N121 = N90 & N32;
  assign N122 = N90 & tag_o[4];
  assign N123 = N92 & N32;
  assign N124 = N92 & tag_o[4];

endmodule

