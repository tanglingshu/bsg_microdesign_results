

module top
(
  lru_i,
  way_id_o
);

  input [126:0] lru_i;
  output [6:0] way_id_o;

  bsg_lru_pseudo_tree_encode
  wrapper
  (
    .lru_i(lru_i),
    .way_id_o(way_id_o)
  );


endmodule



module bsg_lru_pseudo_tree_encode
(
  lru_i,
  way_id_o
);

  input [126:0] lru_i;
  output [6:0] way_id_o;
  wire [6:0] way_id_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
  N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,
  N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,
  N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,
  N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,
  N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,
  N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,
  N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,
  N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,
  N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,
  N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,
  N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,
  N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,
  N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,
  N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,
  N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,
  N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,
  N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
  N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,
  N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,
  N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,
  N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,
  N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,
  N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,
  N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,
  N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,
  N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,
  N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,
  N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,
  N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,
  N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,
  N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,
  N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,
  N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,
  N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,
  N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,
  N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,
  N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,
  N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,
  N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,
  N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,
  N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,
  N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,
  N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,
  N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,
  N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,
  N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,
  N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,
  N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,
  N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,
  N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,
  N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,
  N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,
  N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,
  N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,
  N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,
  N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,
  N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,
  N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,
  N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,
  N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,
  N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,
  N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,
  N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,
  N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,
  N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,
  N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,
  N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,
  N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,
  N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,
  N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,
  N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,
  N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,
  N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,
  N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,
  N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,
  N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,
  N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,
  N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,
  N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,
  N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,
  N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,
  N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,
  N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144,
  N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,
  N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,N2170,
  N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,N2184,
  N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197,
  N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,N2210,
  N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,N2224,
  N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,
  N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,
  N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,N2264,
  N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,
  N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290,
  N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302,N2303,N2304,
  N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,
  N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,
  N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,
  N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,
  N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2369,N2370,
  N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382,N2383,N2384,
  N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,N2394,N2395,N2396,N2397,
  N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407,N2408,N2409,N2410,
  N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422,N2423,N2424,
  N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,
  N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447,N2448,N2449,N2450,
  N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,N2460,N2461,N2462,N2463,N2464,
  N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,N2474,N2475,N2476,N2477,
  N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,N2488,N2489,N2490,
  N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,N2500,N2501,N2502,N2503,N2504,
  N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,N2514,N2515,N2516,N2517,
  N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528,N2529,N2530,
  N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539,N2540,N2541,N2542,N2543,N2544,
  N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2554,N2555,N2556,N2557,
  N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,N2567,N2568,N2569,N2570,
  N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579,N2580,N2581,N2582,N2583,N2584,
  N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,N2594,N2595,N2596,N2597,
  N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,N2609,N2610,
  N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,N2620,N2621,N2622,N2623,N2624,
  N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2637,
  N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,N2649,N2650,
  N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662,N2663,N2664,
  N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,
  N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,N2687,N2688,N2689,N2690,
  N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2704,
  N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,N2714,N2715,N2716,N2717,
  N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,N2727,N2728,N2729,N2730,
  N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,
  N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,N2754,N2755,N2756,N2757,
  N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,N2767,N2768,N2769,N2770,
  N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2779,N2780,N2781,N2782,N2783,N2784,
  N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793,N2794,N2795,N2796,N2797,
  N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,N2807,N2808,N2809,N2810,
  N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,N2819,N2820,N2821,N2822,N2823,N2824,
  N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,N2834,N2835,N2836,N2837,
  N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,N2847,N2848,N2849,N2850,
  N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,N2859,N2860,N2861,N2862,N2863,N2864,
  N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877,
  N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,N2887,N2888,N2889,N2890,
  N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,N2899,N2900,N2901,N2902,N2903,N2904,
  N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,N2917,
  N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,N2930,
  N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,N2939,N2940,N2941,N2942,N2943,N2944,
  N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952,N2953,N2954,N2955,N2956,N2957,
  N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2965,N2966,N2967,N2968,N2969,N2970,
  N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980,N2981,N2982,N2983,N2984,
  N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,
  N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,N3010,
  N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022,N3023,N3024,
  N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3036,N3037,
  N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,N3050,
  N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3062,N3063,N3064,
  N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,N3076,N3077,
  N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,N3090,
  N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,N3101,N3102,N3103,N3104,
  N3105,N3106,N3107,N3108,N3109,N3110,N3111,N3112,N3113,N3114,N3115,N3116,N3117,
  N3118,N3119,N3120,N3121,N3122,N3123,N3124,N3125,N3126,N3127,N3128,N3129,N3130,
  N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,N3139,N3140,N3141,N3142,N3143,N3144,
  N3145,N3146,N3147,N3148,N3149,N3150,N3151,N3152,N3153,N3154,N3155,N3156,N3157,
  N3158,N3159,N3160,N3161,N3162,N3163,N3164,N3165,N3166,N3167,N3168,N3169,N3170,
  N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,N3179,N3180,N3181,N3182,N3183,N3184,
  N3185,N3186,N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194,N3195,N3196,N3197,
  N3198,N3199,N3200,N3201,N3202,N3203,N3204,N3205,N3206,N3207,N3208,N3209,N3210,
  N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,N3220,N3221,N3222,N3223,N3224,
  N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,
  N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,N3249,N3250,
  N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,N3260,N3261,N3262,N3263,N3264,
  N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,
  N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,N3290,
  N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,N3300,N3301,N3302,N3303,N3304,
  N3305,N3306,N3307,N3308,N3309,N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,
  N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,N3330,
  N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,N3339,N3340,N3341,N3342,N3343,N3344,
  N3345,N3346,N3347,N3348,N3349,N3350,N3351,N3352,N3353,N3354,N3355,N3356,N3357,
  N3358,N3359,N3360,N3361,N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,N3370,
  N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,N3379,N3380,N3381,N3382,N3383,N3384,
  N3385,N3386,N3387,N3388,N3389,N3390,N3391,N3392,N3393,N3394,N3395,N3396,N3397,
  N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3408,N3409,N3410,
  N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,N3419,N3420,N3421,N3422,N3423,N3424,
  N3425,N3426,N3427,N3428,N3429,N3430,N3431,N3432,N3433,N3434,N3435,N3436,N3437,
  N3438,N3439,N3440,N3441,N3442,N3443,N3444,N3445,N3446,N3447,N3448,N3449,N3450,
  N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,N3459,N3460,N3461,N3462,N3463,N3464,
  N3465,N3466,N3467,N3468,N3469,N3470,N3471,N3472,N3473,N3474,N3475,N3476,N3477,
  N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,N3487,N3488,N3489,N3490,
  N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,N3499,N3500,N3501,N3502,N3503,N3504,
  N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,N3513,N3514,N3515,N3516,N3517,
  N3518,N3519,N3520,N3521,N3522,N3523,N3524,N3525,N3526,N3527,N3528,N3529,N3530,
  N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,N3539,N3540,N3541,N3542,N3543,N3544,
  N3545,N3546,N3547,N3548,N3549,N3550,N3551,N3552,N3553,N3554,N3555,N3556,N3557,
  N3558,N3559,N3560,N3561,N3562,N3563,N3564,N3565,N3566,N3567,N3568,N3569,N3570,
  N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,N3579,N3580,N3581,N3582,N3583,N3584,
  N3585,N3586,N3587,N3588,N3589,N3590,N3591,N3592,N3593,N3594,N3595,N3596,N3597,
  N3598,N3599,N3600,N3601,N3602,N3603,N3604,N3605,N3606,N3607,N3608,N3609,N3610,
  N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,N3619,N3620,N3621,N3622,N3623,N3624,
  N3625,N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3636,N3637,
  N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3646,N3647,N3648,N3649,N3650,
  N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,N3659,N3660,N3661,N3662,N3663,N3664,
  N3665,N3666,N3667,N3668,N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3676,N3677,
  N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685,N3686,N3687,N3688,N3689,N3690,
  N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,N3699,N3700,N3701,N3702,N3703,N3704,
  N3705,N3706,N3707,N3708,N3709,N3710,N3711,N3712,N3713,N3714,N3715,N3716,N3717,
  N3718,N3719,N3720,N3721,N3722,N3723,N3724,N3725,N3726,N3727,N3728,N3729,N3730,
  N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,N3739,N3740,N3741,N3742,N3743,N3744,
  N3745,N3746,N3747,N3748,N3749,N3750,N3751,N3752,N3753,N3754,N3755,N3756,N3757,
  N3758,N3759,N3760,N3761,N3762,N3763,N3764,N3765,N3766,N3767,N3768,N3769,N3770,
  N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,N3779,N3780,N3781,N3782,N3783,N3784,
  N3785,N3786,N3787,N3788,N3789,N3790,N3791,N3792,N3793,N3794,N3795,N3796,N3797,
  N3798,N3799,N3800,N3801,N3802,N3803,N3804,N3805,N3806,N3807,N3808,N3809,N3810,
  N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,N3819,N3820,N3821,N3822,N3823,N3824,
  N3825,N3826,N3827,N3828,N3829,N3830,N3831,N3832,N3833,N3834,N3835,N3836,N3837,
  N3838,N3839,N3840,N3841,N3842,N3843,N3844,N3845,N3846,N3847,N3848,N3849,N3850,
  N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,N3859,N3860,N3861,N3862,N3863,N3864,
  N3865,N3866,N3867,N3868,N3869,N3870,N3871,N3872,N3873,N3874,N3875,N3876,N3877,
  N3878,N3879,N3880,N3881,N3882,N3883,N3884,N3885,N3886,N3887,N3888,N3889,N3890,
  N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,N3899,N3900,N3901,N3902,N3903,N3904,
  N3905,N3906,N3907,N3908,N3909,N3910,N3911,N3912,N3913,N3914,N3915,N3916,N3917,
  N3918,N3919,N3920,N3921,N3922,N3923,N3924,N3925,N3926,N3927,N3928,N3929,N3930,
  N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,N3939,N3940,N3941,N3942,N3943,N3944,
  N3945,N3946,N3947,N3948,N3949,N3950,N3951,N3952,N3953,N3954,N3955,N3956,N3957,
  N3958,N3959,N3960,N3961,N3962,N3963,N3964,N3965,N3966,N3967,N3968,N3969,N3970,
  N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978,N3979,N3980,N3981,N3982,N3983,N3984,
  N3985,N3986,N3987,N3988,N3989,N3990,N3991,N3992,N3993,N3994,N3995,N3996,N3997,
  N3998,N3999,N4000,N4001,N4002,N4003,N4004,N4005,N4006,N4007,N4008,N4009,N4010,
  N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,N4019,N4020,N4021,N4022,N4023,N4024,
  N4025,N4026,N4027,N4028,N4029,N4030,N4031,N4032,N4033,N4034,N4035,N4036,N4037,
  N4038,N4039,N4040,N4041,N4042,N4043,N4044,N4045,N4046,N4047,N4048,N4049,N4050,
  N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,N4059,N4060,N4061,N4062,N4063,N4064,
  N4065,N4066,N4067,N4068,N4069,N4070,N4071,N4072,N4073,N4074,N4075,N4076,N4077,
  N4078,N4079,N4080,N4081,N4082,N4083,N4084,N4085,N4086,N4087,N4088,N4089,N4090,
  N4091,N4092,N4093,N4094,N4095,N4096,N4097,N4098,N4099,N4100,N4101,N4102,N4103,N4104,
  N4105,N4106,N4107,N4108,N4109,N4110,N4111,N4112,N4113,N4114,N4115,N4116,N4117,
  N4118,N4119,N4120,N4121,N4122,N4123,N4124,N4125,N4126,N4127,N4128,N4129,N4130,
  N4131,N4132,N4133,N4134,N4135,N4136,N4137,N4138,N4139,N4140,N4141,N4142,N4143,N4144,
  N4145,N4146,N4147,N4148,N4149,N4150,N4151,N4152,N4153,N4154,N4155,N4156,N4157,
  N4158,N4159,N4160,N4161,N4162,N4163,N4164,N4165,N4166,N4167,N4168,N4169,N4170,
  N4171,N4172,N4173,N4174,N4175,N4176,N4177,N4178,N4179,N4180,N4181,N4182,N4183,N4184,
  N4185,N4186,N4187,N4188,N4189,N4190,N4191,N4192,N4193,N4194,N4195,N4196,N4197,
  N4198,N4199,N4200,N4201,N4202,N4203,N4204,N4205,N4206,N4207,N4208,N4209,N4210,
  N4211,N4212,N4213,N4214,N4215,N4216,N4217,N4218,N4219,N4220,N4221,N4222,N4223,N4224,
  N4225,N4226,N4227,N4228,N4229,N4230,N4231,N4232,N4233,N4234,N4235,N4236,N4237,
  N4238,N4239,N4240,N4241,N4242,N4243,N4244,N4245,N4246,N4247,N4248,N4249,N4250,
  N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,N4259,N4260,N4261,N4262,N4263,N4264,
  N4265,N4266,N4267,N4268,N4269,N4270,N4271,N4272,N4273,N4274,N4275,N4276,N4277,
  N4278,N4279,N4280,N4281,N4282,N4283,N4284,N4285,N4286,N4287,N4288,N4289,N4290,
  N4291,N4292,N4293,N4294,N4295,N4296,N4297,N4298,N4299,N4300,N4301,N4302,N4303,N4304,
  N4305,N4306,N4307,N4308,N4309,N4310,N4311,N4312,N4313,N4314,N4315,N4316,N4317,
  N4318,N4319,N4320,N4321,N4322,N4323,N4324,N4325,N4326,N4327,N4328,N4329,N4330,
  N4331,N4332,N4333,N4334,N4335,N4336,N4337,N4338,N4339,N4340,N4341,N4342,N4343,N4344,
  N4345,N4346,N4347,N4348,N4349,N4350,N4351,N4352,N4353,N4354,N4355,N4356,N4357,
  N4358,N4359,N4360,N4361,N4362,N4363,N4364,N4365,N4366,N4367,N4368,N4369,N4370,
  N4371,N4372,N4373,N4374,N4375,N4376,N4377,N4378,N4379,N4380,N4381,N4382,N4383,N4384,
  N4385,N4386,N4387,N4388,N4389,N4390,N4391,N4392,N4393,N4394,N4395,N4396,N4397,
  N4398,N4399,N4400,N4401,N4402,N4403,N4404,N4405,N4406,N4407,N4408,N4409,N4410,
  N4411,N4412,N4413,N4414,N4415,N4416,N4417,N4418,N4419,N4420,N4421,N4422,N4423,N4424,
  N4425,N4426,N4427,N4428,N4429,N4430,N4431,N4432,N4433,N4434,N4435,N4436,N4437,
  N4438,N4439,N4440,N4441,N4442,N4443,N4444,N4445,N4446,N4447,N4448,N4449,N4450,
  N4451,N4452,N4453,N4454,N4455,N4456,N4457,N4458,N4459,N4460,N4461,N4462,N4463,N4464,
  N4465,N4466,N4467,N4468,N4469,N4470,N4471,N4472,N4473,N4474,N4475,N4476,N4477,
  N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,N4487,N4488,N4489,N4490,
  N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,N4499,N4500,N4501,N4502,N4503,N4504,
  N4505,N4506,N4507,N4508,N4509,N4510,N4511,N4512,N4513,N4514,N4515,N4516,N4517,
  N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,N4527,N4528,N4529,N4530,
  N4531,N4532,N4533,N4534,N4535,N4536,N4537,N4538,N4539,N4540,N4541,N4542,N4543,N4544,
  N4545,N4546,N4547,N4548,N4549,N4550,N4551,N4552,N4553,N4554,N4555,N4556,N4557,
  N4558,N4559,N4560,N4561,N4562,N4563,N4564,N4565,N4566,N4567,N4568,N4569,N4570,
  N4571,N4572,N4573,N4574,N4575,N4576,N4577,N4578,N4579,N4580,N4581,N4582,N4583,N4584,
  N4585,N4586,N4587,N4588,N4589,N4590,N4591,N4592,N4593,N4594,N4595,N4596,N4597,
  N4598,N4599,N4600,N4601,N4602,N4603,N4604,N4605,N4606,N4607,N4608,N4609,N4610,
  N4611,N4612,N4613,N4614,N4615,N4616,N4617,N4618,N4619,N4620,N4621,N4622,N4623,N4624,
  N4625,N4626,N4627,N4628,N4629,N4630,N4631,N4632,N4633,N4634,N4635,N4636,N4637,
  N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,N4647,N4648,N4649,N4650,
  N4651,N4652,N4653,N4654,N4655,N4656,N4657,N4658,N4659,N4660,N4661,N4662,N4663,N4664,
  N4665,N4666,N4667,N4668,N4669,N4670,N4671,N4672,N4673,N4674,N4675,N4676,N4677,
  N4678,N4679,N4680,N4681,N4682,N4683,N4684,N4685,N4686,N4687,N4688,N4689,N4690,
  N4691,N4692,N4693,N4694,N4695,N4696,N4697,N4698,N4699,N4700,N4701,N4702,N4703,N4704,
  N4705,N4706,N4707,N4708,N4709,N4710,N4711,N4712,N4713,N4714,N4715,N4716,N4717,
  N4718,N4719,N4720,N4721,N4722,N4723,N4724,N4725,N4726,N4727,N4728,N4729,N4730,
  N4731,N4732,N4733,N4734,N4735,N4736,N4737,N4738,N4739,N4740,N4741,N4742,N4743,N4744,
  N4745,N4746,N4747,N4748,N4749,N4750,N4751,N4752,N4753,N4754,N4755,N4756,N4757,
  N4758,N4759,N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,N4768,N4769,N4770,
  N4771,N4772,N4773,N4774,N4775,N4776,N4777,N4778,N4779,N4780,N4781,N4782,N4783,N4784,
  N4785,N4786,N4787,N4788,N4789,N4790,N4791,N4792,N4793,N4794,N4795,N4796,N4797,
  N4798,N4799,N4800,N4801,N4802,N4803,N4804,N4805,N4806,N4807,N4808,N4809,N4810,
  N4811,N4812,N4813,N4814,N4815,N4816,N4817,N4818,N4819,N4820,N4821,N4822,N4823,N4824,
  N4825,N4826,N4827,N4828,N4829,N4830,N4831,N4832,N4833,N4834,N4835,N4836,N4837,
  N4838,N4839,N4840,N4841,N4842,N4843,N4844,N4845,N4846,N4847,N4848,N4849,N4850,
  N4851,N4852,N4853,N4854,N4855,N4856,N4857,N4858,N4859,N4860,N4861,N4862,N4863,N4864,
  N4865,N4866,N4867,N4868,N4869,N4870,N4871,N4872,N4873,N4874,N4875,N4876,N4877,
  N4878,N4879,N4880,N4881,N4882,N4883,N4884,N4885,N4886,N4887,N4888,N4889,N4890,
  N4891,N4892,N4893,N4894,N4895,N4896,N4897,N4898,N4899,N4900,N4901,N4902,N4903,N4904,
  N4905,N4906,N4907,N4908,N4909,N4910,N4911,N4912,N4913,N4914,N4915,N4916,N4917,
  N4918,N4919,N4920,N4921,N4922,N4923,N4924,N4925,N4926,N4927,N4928,N4929,N4930,
  N4931,N4932,N4933,N4934,N4935,N4936,N4937,N4938,N4939,N4940,N4941,N4942,N4943,N4944,
  N4945,N4946,N4947,N4948,N4949,N4950,N4951,N4952,N4953,N4954,N4955,N4956,N4957,
  N4958,N4959,N4960,N4961,N4962,N4963,N4964,N4965,N4966,N4967,N4968,N4969,N4970,
  N4971,N4972,N4973,N4974,N4975,N4976,N4977,N4978,N4979,N4980,N4981,N4982,N4983,N4984,
  N4985,N4986,N4987,N4988,N4989,N4990,N4991,N4992,N4993,N4994,N4995,N4996,N4997,
  N4998,N4999,N5000,N5001,N5002,N5003,N5004,N5005,N5006,N5007,N5008,N5009,N5010,
  N5011,N5012,N5013,N5014,N5015,N5016,N5017,N5018,N5019,N5020,N5021,N5022,N5023,N5024,
  N5025,N5026,N5027,N5028,N5029,N5030,N5031,N5032,N5033,N5034,N5035,N5036,N5037,
  N5038,N5039,N5040,N5041,N5042,N5043,N5044,N5045,N5046,N5047,N5048,N5049,N5050,
  N5051,N5052,N5053,N5054,N5055,N5056,N5057,N5058,N5059,N5060,N5061,N5062,N5063,N5064,
  N5065,N5066,N5067,N5068,N5069,N5070,N5071,N5072,N5073,N5074,N5075,N5076,N5077,
  N5078,N5079,N5080,N5081,N5082,N5083,N5084,N5085,N5086,N5087,N5088,N5089,N5090,
  N5091,N5092,N5093,N5094,N5095,N5096,N5097,N5098,N5099,N5100,N5101,N5102,N5103,N5104,
  N5105,N5106,N5107,N5108,N5109,N5110,N5111,N5112,N5113,N5114,N5115,N5116,N5117,
  N5118,N5119,N5120,N5121,N5122,N5123,N5124,N5125,N5126,N5127,N5128,N5129,N5130,
  N5131,N5132,N5133,N5134,N5135,N5136,N5137,N5138,N5139,N5140,N5141,N5142,N5143,N5144,
  N5145,N5146,N5147,N5148,N5149,N5150,N5151,N5152,N5153,N5154,N5155,N5156,N5157,
  N5158,N5159,N5160,N5161,N5162,N5163,N5164,N5165,N5166,N5167,N5168,N5169,N5170,
  N5171,N5172,N5173,N5174,N5175,N5176,N5177,N5178,N5179,N5180,N5181,N5182,N5183,N5184,
  N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,N5193,N5194,N5195,N5196,N5197,
  N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,N5207,N5208,N5209,N5210,
  N5211,N5212,N5213,N5214,N5215,N5216,N5217,N5218,N5219,N5220,N5221,N5222,N5223,N5224,
  N5225,N5226,N5227,N5228,N5229,N5230,N5231,N5232,N5233,N5234,N5235,N5236,N5237,
  N5238,N5239,N5240,N5241,N5242,N5243,N5244,N5245,N5246,N5247,N5248,N5249,N5250,
  N5251,N5252,N5253,N5254,N5255,N5256,N5257,N5258,N5259,N5260,N5261,N5262,N5263,N5264,
  N5265,N5266,N5267,N5268,N5269,N5270,N5271,N5272,N5273,N5274,N5275,N5276,N5277,
  N5278,N5279,N5280,N5281,N5282,N5283,N5284,N5285,N5286,N5287,N5288,N5289,N5290,
  N5291,N5292,N5293,N5294,N5295,N5296,N5297,N5298,N5299,N5300,N5301,N5302,N5303,N5304,
  N5305,N5306,N5307,N5308,N5309,N5310,N5311,N5312,N5313,N5314,N5315,N5316,N5317,
  N5318,N5319,N5320,N5321,N5322,N5323,N5324,N5325,N5326,N5327,N5328,N5329,N5330,
  N5331,N5332,N5333,N5334,N5335,N5336,N5337,N5338,N5339,N5340,N5341,N5342,N5343,N5344,
  N5345,N5346,N5347,N5348,N5349,N5350,N5351,N5352,N5353,N5354,N5355,N5356,N5357,
  N5358,N5359,N5360,N5361,N5362,N5363,N5364,N5365,N5366,N5367,N5368,N5369,N5370,
  N5371,N5372,N5373,N5374,N5375,N5376,N5377,N5378,N5379,N5380,N5381,N5382,N5383,N5384,
  N5385,N5386,N5387,N5388,N5389,N5390,N5391,N5392,N5393,N5394,N5395,N5396,N5397,
  N5398,N5399,N5400,N5401,N5402,N5403,N5404,N5405,N5406,N5407,N5408,N5409,N5410,
  N5411,N5412,N5413,N5414,N5415,N5416,N5417,N5418,N5419,N5420,N5421,N5422,N5423,N5424,
  N5425,N5426,N5427,N5428,N5429,N5430,N5431,N5432,N5433,N5434,N5435,N5436,N5437,
  N5438,N5439,N5440,N5441,N5442,N5443,N5444,N5445,N5446,N5447,N5448,N5449,N5450,
  N5451,N5452,N5453,N5454,N5455,N5456,N5457,N5458,N5459,N5460,N5461,N5462,N5463,N5464,
  N5465,N5466,N5467,N5468,N5469,N5470,N5471,N5472,N5473,N5474,N5475,N5476,N5477,
  N5478,N5479,N5480,N5481,N5482,N5483,N5484,N5485,N5486,N5487,N5488,N5489,N5490,
  N5491,N5492,N5493,N5494,N5495,N5496,N5497,N5498,N5499,N5500,N5501,N5502,N5503,N5504,
  N5505,N5506,N5507,N5508,N5509,N5510,N5511,N5512,N5513,N5514,N5515,N5516,N5517,
  N5518,N5519,N5520,N5521,N5522,N5523,N5524,N5525,N5526,N5527,N5528,N5529,N5530,
  N5531,N5532,N5533,N5534,N5535,N5536,N5537,N5538,N5539,N5540,N5541,N5542,N5543,N5544,
  N5545,N5546,N5547,N5548,N5549,N5550,N5551,N5552,N5553,N5554,N5555,N5556,N5557,
  N5558,N5559,N5560,N5561,N5562,N5563,N5564,N5565,N5566,N5567,N5568,N5569,N5570,
  N5571,N5572,N5573,N5574,N5575,N5576,N5577,N5578,N5579,N5580,N5581,N5582,N5583,N5584,
  N5585,N5586,N5587,N5588,N5589,N5590,N5591,N5592,N5593,N5594,N5595,N5596,N5597,
  N5598,N5599,N5600,N5601,N5602,N5603,N5604,N5605,N5606,N5607,N5608,N5609,N5610,
  N5611,N5612,N5613,N5614,N5615,N5616,N5617,N5618,N5619,N5620,N5621,N5622,N5623,N5624,
  N5625,N5626,N5627,N5628,N5629,N5630,N5631,N5632,N5633,N5634,N5635,N5636,N5637,
  N5638,N5639,N5640,N5641,N5642,N5643,N5644,N5645,N5646,N5647,N5648,N5649,N5650,
  N5651,N5652,N5653,N5654,N5655,N5656,N5657,N5658,N5659,N5660,N5661,N5662,N5663,N5664,
  N5665,N5666,N5667,N5668,N5669,N5670,N5671,N5672,N5673,N5674,N5675,N5676,N5677,
  N5678,N5679,N5680,N5681,N5682,N5683,N5684,N5685,N5686,N5687,N5688,N5689,N5690,
  N5691,N5692,N5693,N5694,N5695,N5696,N5697,N5698,N5699,N5700,N5701,N5702,N5703,N5704,
  N5705,N5706,N5707,N5708,N5709,N5710,N5711,N5712,N5713,N5714,N5715,N5716,N5717,
  N5718,N5719,N5720,N5721,N5722,N5723,N5724,N5725,N5726,N5727,N5728,N5729,N5730,
  N5731,N5732,N5733,N5734,N5735,N5736,N5737,N5738,N5739,N5740,N5741,N5742,N5743,N5744,
  N5745,N5746,N5747,N5748,N5749,N5750,N5751,N5752,N5753,N5754,N5755,N5756,N5757,
  N5758,N5759,N5760,N5761,N5762,N5763,N5764,N5765,N5766,N5767,N5768,N5769,N5770,
  N5771,N5772,N5773,N5774,N5775,N5776,N5777,N5778,N5779,N5780,N5781,N5782,N5783,N5784,
  N5785,N5786,N5787,N5788,N5789,N5790,N5791,N5792,N5793,N5794,N5795,N5796,N5797,
  N5798,N5799,N5800,N5801,N5802,N5803,N5804,N5805,N5806,N5807,N5808,N5809,N5810,
  N5811,N5812,N5813,N5814,N5815,N5816,N5817,N5818,N5819,N5820,N5821,N5822,N5823,N5824,
  N5825,N5826,N5827,N5828,N5829,N5830,N5831,N5832,N5833,N5834,N5835,N5836,N5837,
  N5838,N5839,N5840,N5841,N5842,N5843,N5844,N5845,N5846,N5847,N5848,N5849,N5850,
  N5851,N5852,N5853,N5854,N5855,N5856,N5857,N5858,N5859,N5860,N5861,N5862,N5863,N5864,
  N5865,N5866,N5867,N5868,N5869,N5870,N5871,N5872,N5873,N5874,N5875,N5876,N5877,
  N5878,N5879,N5880,N5881,N5882,N5883,N5884,N5885,N5886,N5887,N5888,N5889,N5890,
  N5891,N5892,N5893,N5894,N5895,N5896,N5897,N5898,N5899,N5900,N5901,N5902,N5903,N5904,
  N5905,N5906,N5907,N5908,N5909,N5910,N5911,N5912,N5913,N5914,N5915,N5916,N5917,
  N5918,N5919,N5920,N5921,N5922,N5923,N5924,N5925,N5926,N5927,N5928,N5929,N5930,
  N5931,N5932,N5933,N5934,N5935,N5936,N5937,N5938,N5939,N5940,N5941,N5942,N5943,N5944,
  N5945,N5946,N5947,N5948,N5949,N5950,N5951,N5952,N5953,N5954,N5955,N5956,N5957,
  N5958,N5959,N5960,N5961,N5962,N5963,N5964,N5965,N5966,N5967,N5968,N5969,N5970,
  N5971,N5972,N5973,N5974,N5975,N5976,N5977,N5978,N5979,N5980,N5981,N5982,N5983,N5984,
  N5985,N5986,N5987,N5988,N5989,N5990,N5991,N5992,N5993,N5994,N5995,N5996,N5997,
  N5998,N5999,N6000,N6001,N6002,N6003,N6004,N6005,N6006,N6007,N6008,N6009,N6010,
  N6011,N6012,N6013,N6014,N6015,N6016,N6017,N6018,N6019,N6020,N6021,N6022,N6023,N6024,
  N6025,N6026,N6027,N6028,N6029,N6030,N6031,N6032,N6033,N6034,N6035,N6036,N6037,
  N6038,N6039,N6040,N6041,N6042,N6043,N6044,N6045,N6046,N6047,N6048,N6049,N6050,
  N6051,N6052,N6053,N6054,N6055,N6056,N6057,N6058,N6059,N6060,N6061,N6062,N6063,N6064,
  N6065,N6066,N6067,N6068,N6069,N6070,N6071,N6072,N6073,N6074,N6075,N6076,N6077,
  N6078,N6079,N6080,N6081,N6082,N6083,N6084,N6085,N6086,N6087,N6088,N6089,N6090,
  N6091,N6092,N6093,N6094,N6095,N6096,N6097,N6098,N6099,N6100,N6101,N6102,N6103,N6104,
  N6105,N6106,N6107,N6108,N6109,N6110,N6111,N6112,N6113,N6114,N6115,N6116,N6117,
  N6118,N6119,N6120,N6121,N6122,N6123,N6124,N6125,N6126,N6127,N6128,N6129,N6130,
  N6131,N6132,N6133,N6134,N6135,N6136,N6137,N6138,N6139,N6140,N6141,N6142,N6143,N6144,
  N6145,N6146,N6147,N6148,N6149,N6150,N6151,N6152,N6153,N6154,N6155,N6156,N6157,
  N6158,N6159,N6160,N6161,N6162,N6163,N6164,N6165,N6166,N6167,N6168,N6169,N6170,
  N6171,N6172,N6173,N6174,N6175,N6176,N6177,N6178,N6179,N6180,N6181,N6182,N6183,N6184,
  N6185,N6186,N6187,N6188,N6189,N6190,N6191,N6192,N6193,N6194,N6195,N6196,N6197,
  N6198,N6199,N6200,N6201,N6202,N6203,N6204,N6205,N6206,N6207,N6208,N6209,N6210,
  N6211,N6212,N6213,N6214,N6215,N6216,N6217,N6218,N6219,N6220,N6221,N6222,N6223,N6224,
  N6225,N6226,N6227,N6228,N6229,N6230,N6231,N6232,N6233,N6234,N6235,N6236,N6237,
  N6238,N6239,N6240,N6241,N6242,N6243,N6244,N6245,N6246,N6247,N6248,N6249,N6250,
  N6251,N6252,N6253,N6254,N6255,N6256,N6257,N6258,N6259,N6260,N6261,N6262,N6263,N6264,
  N6265,N6266,N6267,N6268,N6269,N6270,N6271,N6272,N6273,N6274,N6275,N6276,N6277,
  N6278,N6279,N6280,N6281,N6282,N6283,N6284,N6285,N6286,N6287,N6288,N6289,N6290,
  N6291,N6292,N6293,N6294,N6295,N6296,N6297,N6298,N6299,N6300,N6301,N6302,N6303,N6304,
  N6305,N6306,N6307,N6308,N6309,N6310,N6311,N6312,N6313,N6314,N6315,N6316,N6317,
  N6318,N6319,N6320,N6321,N6322,N6323,N6324,N6325,N6326,N6327,N6328,N6329,N6330,
  N6331,N6332,N6333,N6334,N6335,N6336,N6337,N6338,N6339,N6340,N6341,N6342,N6343,N6344,
  N6345,N6346,N6347,N6348,N6349,N6350,N6351,N6352,N6353,N6354,N6355,N6356,N6357,
  N6358,N6359,N6360,N6361,N6362,N6363,N6364,N6365,N6366,N6367,N6368,N6369,N6370,
  N6371,N6372,N6373,N6374,N6375,N6376,N6377,N6378,N6379,N6380,N6381,N6382,N6383,N6384,
  N6385,N6386,N6387,N6388,N6389,N6390,N6391,N6392,N6393,N6394,N6395,N6396,N6397,
  N6398,N6399,N6400,N6401,N6402,N6403,N6404,N6405,N6406,N6407,N6408,N6409,N6410,
  N6411,N6412,N6413,N6414,N6415,N6416,N6417,N6418,N6419,N6420,N6421,N6422,N6423,N6424,
  N6425,N6426,N6427,N6428,N6429,N6430,N6431,N6432,N6433,N6434,N6435,N6436,N6437,
  N6438,N6439,N6440,N6441,N6442,N6443,N6444,N6445,N6446,N6447,N6448,N6449,N6450,
  N6451,N6452,N6453,N6454,N6455,N6456,N6457,N6458,N6459,N6460,N6461,N6462,N6463,N6464,
  N6465,N6466,N6467,N6468,N6469,N6470,N6471,N6472,N6473,N6474,N6475,N6476,N6477,
  N6478,N6479,N6480,N6481,N6482,N6483,N6484,N6485,N6486,N6487,N6488,N6489,N6490,
  N6491,N6492,N6493,N6494,N6495,N6496,N6497,N6498,N6499,N6500,N6501,N6502,N6503,N6504,
  N6505,N6506,N6507,N6508,N6509,N6510,N6511,N6512,N6513,N6514,N6515,N6516,N6517,
  N6518,N6519,N6520,N6521,N6522,N6523,N6524,N6525,N6526,N6527,N6528,N6529,N6530,
  N6531,N6532,N6533,N6534,N6535,N6536,N6537,N6538,N6539,N6540,N6541,N6542,N6543,N6544,
  N6545,N6546,N6547,N6548,N6549,N6550,N6551,N6552,N6553,N6554,N6555,N6556,N6557,
  N6558,N6559,N6560,N6561,N6562,N6563,N6564,N6565,N6566,N6567,N6568,N6569,N6570,
  N6571,N6572,N6573,N6574,N6575,N6576,N6577,N6578,N6579,N6580,N6581,N6582,N6583,N6584,
  N6585,N6586,N6587,N6588,N6589,N6590,N6591,N6592,N6593,N6594,N6595,N6596,N6597,
  N6598,N6599,N6600,N6601,N6602,N6603,N6604,N6605,N6606,N6607,N6608,N6609,N6610,
  N6611,N6612,N6613,N6614,N6615,N6616,N6617,N6618,N6619,N6620,N6621,N6622,N6623,N6624,
  N6625,N6626,N6627,N6628,N6629,N6630,N6631,N6632,N6633,N6634,N6635,N6636,N6637,
  N6638,N6639,N6640,N6641,N6642,N6643,N6644,N6645,N6646,N6647,N6648,N6649,N6650,
  N6651,N6652,N6653,N6654,N6655,N6656,N6657,N6658,N6659,N6660,N6661,N6662,N6663,N6664,
  N6665,N6666,N6667,N6668,N6669,N6670,N6671,N6672,N6673,N6674,N6675,N6676,N6677,
  N6678,N6679,N6680,N6681,N6682,N6683,N6684,N6685,N6686,N6687,N6688,N6689,N6690,
  N6691,N6692,N6693,N6694,N6695,N6696,N6697,N6698,N6699,N6700,N6701,N6702,N6703,N6704,
  N6705,N6706,N6707,N6708,N6709,N6710,N6711,N6712,N6713,N6714,N6715,N6716,N6717,
  N6718,N6719,N6720,N6721,N6722,N6723,N6724,N6725,N6726,N6727,N6728,N6729,N6730,
  N6731,N6732,N6733,N6734,N6735,N6736,N6737,N6738,N6739,N6740,N6741,N6742,N6743,N6744,
  N6745,N6746,N6747,N6748,N6749,N6750,N6751,N6752,N6753,N6754,N6755,N6756,N6757,
  N6758,N6759,N6760,N6761,N6762,N6763,N6764,N6765,N6766,N6767,N6768,N6769,N6770,
  N6771,N6772,N6773,N6774,N6775,N6776,N6777,N6778,N6779,N6780,N6781,N6782,N6783,N6784,
  N6785,N6786,N6787,N6788,N6789,N6790,N6791,N6792,N6793,N6794,N6795,N6796,N6797,
  N6798,N6799,N6800,N6801,N6802,N6803,N6804,N6805,N6806,N6807,N6808,N6809,N6810,
  N6811,N6812,N6813,N6814,N6815,N6816,N6817,N6818,N6819,N6820,N6821,N6822,N6823,N6824,
  N6825,N6826,N6827,N6828,N6829,N6830,N6831,N6832,N6833,N6834,N6835,N6836,N6837,
  N6838,N6839,N6840,N6841,N6842,N6843,N6844,N6845,N6846,N6847,N6848,N6849,N6850,
  N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6858,N6859,N6860,N6861,N6862,N6863,N6864,
  N6865,N6866,N6867,N6868,N6869,N6870,N6871,N6872,N6873,N6874,N6875,N6876,N6877,
  N6878,N6879,N6880,N6881,N6882,N6883,N6884,N6885,N6886,N6887,N6888,N6889,N6890,
  N6891,N6892,N6893,N6894,N6895,N6896,N6897,N6898,N6899,N6900,N6901,N6902,N6903,N6904,
  N6905,N6906,N6907,N6908,N6909,N6910,N6911,N6912,N6913,N6914,N6915,N6916,N6917,
  N6918,N6919,N6920,N6921,N6922,N6923,N6924,N6925,N6926,N6927,N6928,N6929,N6930,
  N6931,N6932,N6933,N6934,N6935,N6936,N6937,N6938,N6939,N6940,N6941,N6942,N6943,N6944,
  N6945,N6946,N6947,N6948,N6949,N6950,N6951,N6952,N6953,N6954,N6955,N6956,N6957,
  N6958,N6959,N6960,N6961,N6962,N6963,N6964,N6965,N6966,N6967,N6968,N6969,N6970,
  N6971,N6972,N6973,N6974,N6975,N6976,N6977,N6978,N6979,N6980,N6981,N6982,N6983,N6984,
  N6985,N6986,N6987,N6988,N6989,N6990,N6991,N6992,N6993,N6994,N6995,N6996,N6997,
  N6998,N6999,N7000,N7001,N7002,N7003,N7004,N7005,N7006,N7007,N7008,N7009,N7010,
  N7011,N7012,N7013,N7014,N7015,N7016,N7017,N7018,N7019,N7020,N7021,N7022,N7023,N7024,
  N7025,N7026,N7027,N7028,N7029,N7030,N7031,N7032,N7033,N7034,N7035,N7036,N7037,
  N7038,N7039,N7040,N7041,N7042,N7043,N7044,N7045,N7046,N7047,N7048,N7049,N7050,
  N7051,N7052,N7053,N7054,N7055,N7056,N7057,N7058,N7059,N7060,N7061,N7062,N7063,N7064,
  N7065,N7066,N7067,N7068,N7069,N7070,N7071,N7072,N7073,N7074,N7075,N7076,N7077,
  N7078,N7079,N7080,N7081,N7082,N7083,N7084,N7085,N7086,N7087,N7088,N7089,N7090,
  N7091,N7092,N7093,N7094,N7095,N7096,N7097,N7098,N7099,N7100,N7101,N7102,N7103,N7104,
  N7105,N7106,N7107,N7108,N7109,N7110,N7111,N7112,N7113,N7114,N7115,N7116,N7117,
  N7118,N7119,N7120,N7121,N7122,N7123,N7124,N7125,N7126,N7127,N7128,N7129,N7130,
  N7131,N7132,N7133,N7134,N7135,N7136,N7137,N7138,N7139,N7140,N7141,N7142,N7143,N7144,
  N7145,N7146,N7147,N7148,N7149,N7150,N7151,N7152,N7153,N7154,N7155,N7156,N7157,
  N7158,N7159,N7160,N7161,N7162,N7163,N7164,N7165,N7166,N7167,N7168,N7169,N7170,
  N7171,N7172,N7173,N7174,N7175,pe_o_6__6_,pe_o_6__5_,pe_o_6__4_,pe_o_6__3_,
  pe_o_6__2_,pe_o_6__1_,pe_o_6__0_,pe_o_5__6_,pe_o_5__5_,pe_o_5__4_,pe_o_5__3_,pe_o_5__2_,
  pe_o_5__1_,pe_o_5__0_,pe_o_4__6_,pe_o_4__5_,pe_o_4__4_,pe_o_4__3_,pe_o_4__2_,
  pe_o_4__1_,pe_o_4__0_,pe_o_3__6_,pe_o_3__5_,pe_o_3__4_,pe_o_3__3_,pe_o_3__2_,
  pe_o_3__1_,pe_o_3__0_,pe_o_2__6_,pe_o_2__5_,pe_o_2__4_,pe_o_2__3_,pe_o_2__2_,pe_o_2__1_,
  pe_o_2__0_,pe_o_1__6_,pe_o_1__5_,pe_o_1__4_,pe_o_1__3_,pe_o_1__2_,pe_o_1__1_,
  pe_o_1__0_,N7176,N7177,N7178,N7179,N7180,N7181,N7182,N7183,N7184,N7185,N7186,N7187,
  N7188,N7189,N7190,N7191,N7192,N7193,N7194,N7195,N7196,N7197,N7198,N7199,N7200,
  N7201,N7202,N7203,N7204,N7205,N7206,N7207,N7208,N7209,N7210,N7211,N7212,N7213,
  N7214,N7215,N7216,N7217,N7218,N7219,N7220,N7221,N7222,N7223,N7224,N7225,N7226,N7227,
  N7228,N7229,N7230,N7231,N7232,N7233,N7234,N7235,N7236,N7237,N7238,N7239,N7240,
  N7241,N7242,N7243,N7244,N7245,N7246,N7247,N7248,N7249,N7250,N7251,N7252,N7253,
  N7254,N7255,N7256,N7257,N7258,N7259,N7260,N7261,N7262,N7263,N7264,N7265,N7266,N7267,
  N7268,N7269,N7270,N7271,N7272,N7273,N7274,N7275,N7276,N7277,N7278,N7279,N7280,
  N7281,N7282,N7283,N7284,N7285,N7286,N7287,N7288,N7289,N7290,N7291,N7292,N7293,
  N7294,N7295,N7296,N7297,N7298,N7299,N7300,N7301,N7302,N7303,N7304,N7305,N7306,N7307,
  N7308,N7309,N7310,N7311,N7312,N7313,N7314,N7315,N7316,N7317,N7318,N7319,N7320,
  N7321,N7322,N7323,N7324,N7325,N7326,N7327,N7328,N7329,N7330,N7331,N7332,N7333,
  N7334,N7335,N7336,N7337,N7338,N7339,N7340,N7341,N7342,N7343,N7344,N7345,N7346,N7347,
  N7348,N7349,N7350,N7351,N7352,N7353,N7354,N7355,N7356,N7357,N7358,N7359,N7360,
  N7361,N7362,N7363,N7364,N7365,N7366,N7367,N7368,N7369,N7370,N7371,N7372,N7373,
  N7374,N7375,N7376,N7377,N7378,N7379,N7380,N7381,N7382,N7383,N7384,N7385,N7386,N7387,
  N7388,N7389,N7390,N7391,N7392,N7393,N7394,N7395,N7396,N7397,N7398,N7399,N7400,
  N7401,N7402,N7403,N7404,N7405,N7406,N7407,N7408,N7409,N7410,N7411,N7412,N7413,
  N7414,N7415,N7416,N7417,N7418,N7419,N7420,N7421,N7422,N7423,N7424,N7425,N7426,N7427,
  pe_i_6__126_,pe_i_6__125_,pe_i_6__124_,pe_i_6__123_,pe_i_6__122_,pe_i_6__121_,
  pe_i_6__120_,pe_i_6__119_,pe_i_6__118_,pe_i_6__117_,pe_i_6__116_,pe_i_6__115_,
  pe_i_6__114_,pe_i_6__113_,pe_i_6__112_,pe_i_6__111_,pe_i_6__110_,pe_i_6__109_,
  pe_i_6__108_,pe_i_6__107_,pe_i_6__106_,pe_i_6__105_,pe_i_6__104_,pe_i_6__103_,
  pe_i_6__102_,pe_i_6__101_,pe_i_6__100_,pe_i_6__99_,pe_i_6__98_,pe_i_6__97_,pe_i_6__96_,
  pe_i_6__95_,pe_i_6__94_,pe_i_6__93_,pe_i_6__92_,pe_i_6__91_,pe_i_6__90_,
  pe_i_6__89_,pe_i_6__88_,pe_i_6__87_,pe_i_6__86_,pe_i_6__85_,pe_i_6__84_,pe_i_6__83_,
  pe_i_6__82_,pe_i_6__81_,pe_i_6__80_,pe_i_6__79_,pe_i_6__78_,pe_i_6__77_,pe_i_6__76_,
  pe_i_6__75_,pe_i_6__74_,pe_i_6__73_,pe_i_6__72_,pe_i_6__71_,pe_i_6__70_,
  pe_i_6__69_,pe_i_6__68_,pe_i_6__67_,pe_i_6__66_,pe_i_6__65_,pe_i_6__64_,pe_i_6__63_,
  pe_i_6__62_,pe_i_6__61_,pe_i_6__60_,pe_i_6__59_,pe_i_6__58_,pe_i_6__57_,pe_i_6__56_,
  pe_i_6__55_,pe_i_6__54_,pe_i_6__53_,pe_i_6__52_,pe_i_6__51_,pe_i_6__50_,
  pe_i_6__49_,pe_i_6__48_,pe_i_6__47_,pe_i_6__46_,pe_i_6__45_,pe_i_6__44_,pe_i_6__43_,
  pe_i_6__42_,pe_i_6__41_,pe_i_6__40_,pe_i_6__39_,pe_i_6__38_,pe_i_6__37_,pe_i_6__36_,
  pe_i_6__35_,pe_i_6__34_,pe_i_6__33_,pe_i_6__32_,pe_i_6__31_,pe_i_6__30_,
  pe_i_6__29_,pe_i_6__28_,pe_i_6__27_,pe_i_6__26_,pe_i_6__25_,pe_i_6__24_,pe_i_6__23_,
  pe_i_6__22_,pe_i_6__21_,pe_i_6__20_,pe_i_6__19_,pe_i_6__18_,pe_i_6__17_,pe_i_6__16_,
  pe_i_6__15_,pe_i_6__14_,pe_i_6__13_,pe_i_6__12_,pe_i_6__11_,pe_i_6__10_,
  pe_i_6__9_,pe_i_6__8_,pe_i_6__7_,pe_i_6__6_,pe_i_6__5_,pe_i_6__4_,pe_i_6__3_,pe_i_6__2_,
  pe_i_6__1_,pe_i_6__0_,pe_i_5__126_,pe_i_5__125_,pe_i_5__124_,pe_i_5__123_,
  pe_i_5__122_,pe_i_5__121_,pe_i_5__120_,pe_i_5__119_,pe_i_5__118_,pe_i_5__117_,
  pe_i_5__116_,pe_i_5__115_,pe_i_5__114_,pe_i_5__113_,pe_i_5__112_,pe_i_5__111_,
  pe_i_5__110_,pe_i_5__109_,pe_i_5__108_,pe_i_5__107_,pe_i_5__106_,pe_i_5__105_,pe_i_5__104_,
  pe_i_5__103_,pe_i_5__102_,pe_i_5__101_,pe_i_5__100_,pe_i_5__99_,pe_i_5__98_,
  pe_i_5__97_,pe_i_5__96_,pe_i_5__95_,pe_i_5__94_,pe_i_5__93_,pe_i_5__92_,pe_i_5__91_,
  pe_i_5__90_,pe_i_5__89_,pe_i_5__88_,pe_i_5__87_,pe_i_5__86_,pe_i_5__85_,
  pe_i_5__84_,pe_i_5__83_,pe_i_5__82_,pe_i_5__81_,pe_i_5__80_,pe_i_5__79_,pe_i_5__78_,
  pe_i_5__77_,pe_i_5__76_,pe_i_5__75_,pe_i_5__74_,pe_i_5__73_,pe_i_5__72_,pe_i_5__71_,
  pe_i_5__70_,pe_i_5__69_,pe_i_5__68_,pe_i_5__67_,pe_i_5__66_,pe_i_5__65_,
  pe_i_5__64_,pe_i_5__63_,pe_i_5__62_,pe_i_5__61_,pe_i_5__60_,pe_i_5__59_,pe_i_5__58_,
  pe_i_5__57_,pe_i_5__56_,pe_i_5__55_,pe_i_5__54_,pe_i_5__53_,pe_i_5__52_,pe_i_5__51_,
  pe_i_5__50_,pe_i_5__49_,pe_i_5__48_,pe_i_5__47_,pe_i_5__46_,pe_i_5__45_,
  pe_i_5__44_,pe_i_5__43_,pe_i_5__42_,pe_i_5__41_,pe_i_5__40_,pe_i_5__39_,pe_i_5__38_,
  pe_i_5__37_,pe_i_5__36_,pe_i_5__35_,pe_i_5__34_,pe_i_5__33_,pe_i_5__32_,pe_i_5__31_,
  pe_i_5__30_,pe_i_5__29_,pe_i_5__28_,pe_i_5__27_,pe_i_5__26_,pe_i_5__25_,
  pe_i_5__24_,pe_i_5__23_,pe_i_5__22_,pe_i_5__21_,pe_i_5__20_,pe_i_5__19_,pe_i_5__18_,
  pe_i_5__17_,pe_i_5__16_,pe_i_5__15_,pe_i_5__14_,pe_i_5__13_,pe_i_5__12_,pe_i_5__11_,
  pe_i_5__10_,pe_i_5__9_,pe_i_5__8_,pe_i_5__7_,pe_i_5__6_,pe_i_5__5_,pe_i_5__4_,
  pe_i_5__3_,pe_i_5__2_,pe_i_5__1_,pe_i_5__0_,pe_i_4__126_,pe_i_4__125_,
  pe_i_4__124_,pe_i_4__123_,pe_i_4__122_,pe_i_4__121_,pe_i_4__120_,pe_i_4__119_,pe_i_4__118_,
  pe_i_4__117_,pe_i_4__116_,pe_i_4__115_,pe_i_4__114_,pe_i_4__113_,pe_i_4__112_,
  pe_i_4__111_,pe_i_4__110_,pe_i_4__109_,pe_i_4__108_,pe_i_4__107_,pe_i_4__106_,
  pe_i_4__105_,pe_i_4__104_,pe_i_4__103_,pe_i_4__102_,pe_i_4__101_,pe_i_4__100_,
  pe_i_4__99_,pe_i_4__98_,pe_i_4__97_,pe_i_4__96_,pe_i_4__95_,pe_i_4__94_,pe_i_4__93_,
  pe_i_4__92_,pe_i_4__91_,pe_i_4__90_,pe_i_4__89_,pe_i_4__88_,pe_i_4__87_,
  pe_i_4__86_,pe_i_4__85_,pe_i_4__84_,pe_i_4__83_,pe_i_4__82_,pe_i_4__81_,pe_i_4__80_,
  pe_i_4__79_,pe_i_4__78_,pe_i_4__77_,pe_i_4__76_,pe_i_4__75_,pe_i_4__74_,pe_i_4__73_,
  pe_i_4__72_,pe_i_4__71_,pe_i_4__70_,pe_i_4__69_,pe_i_4__68_,pe_i_4__67_,
  pe_i_4__66_,pe_i_4__65_,pe_i_4__64_,pe_i_4__63_,pe_i_4__62_,pe_i_4__61_,pe_i_4__60_,
  pe_i_4__59_,pe_i_4__58_,pe_i_4__57_,pe_i_4__56_,pe_i_4__55_,pe_i_4__54_,pe_i_4__53_,
  pe_i_4__52_,pe_i_4__51_,pe_i_4__50_,pe_i_4__49_,pe_i_4__48_,pe_i_4__47_,
  pe_i_4__46_,pe_i_4__45_,pe_i_4__44_,pe_i_4__43_,pe_i_4__42_,pe_i_4__41_,pe_i_4__40_,
  pe_i_4__39_,pe_i_4__38_,pe_i_4__37_,pe_i_4__36_,pe_i_4__35_,pe_i_4__34_,pe_i_4__33_,
  pe_i_4__32_,pe_i_4__31_,pe_i_4__30_,pe_i_4__29_,pe_i_4__28_,pe_i_4__27_,
  pe_i_4__26_,pe_i_4__25_,pe_i_4__24_,pe_i_4__23_,pe_i_4__22_,pe_i_4__21_,pe_i_4__20_,
  pe_i_4__19_,pe_i_4__18_,pe_i_4__17_,pe_i_4__16_,pe_i_4__15_,pe_i_4__14_,pe_i_4__13_,
  pe_i_4__12_,pe_i_4__11_,pe_i_4__10_,pe_i_4__9_,pe_i_4__8_,pe_i_4__7_,pe_i_4__6_,
  pe_i_4__5_,pe_i_4__4_,pe_i_4__3_,pe_i_4__2_,pe_i_4__1_,pe_i_4__0_,pe_i_3__126_,
  pe_i_3__125_,pe_i_3__124_,pe_i_3__123_,pe_i_3__122_,pe_i_3__121_,pe_i_3__120_,
  pe_i_3__119_,pe_i_3__118_,pe_i_3__117_,pe_i_3__116_,pe_i_3__115_,pe_i_3__114_,
  pe_i_3__113_,pe_i_3__112_,pe_i_3__111_,pe_i_3__110_,pe_i_3__109_,pe_i_3__108_,
  pe_i_3__107_,pe_i_3__106_,pe_i_3__105_,pe_i_3__104_,pe_i_3__103_,pe_i_3__102_,
  pe_i_3__101_,pe_i_3__100_,pe_i_3__99_,pe_i_3__98_,pe_i_3__97_,pe_i_3__96_,pe_i_3__95_,
  pe_i_3__94_,pe_i_3__93_,pe_i_3__92_,pe_i_3__91_,pe_i_3__90_,pe_i_3__89_,pe_i_3__88_,
  pe_i_3__87_,pe_i_3__86_,pe_i_3__85_,pe_i_3__84_,pe_i_3__83_,pe_i_3__82_,
  pe_i_3__81_,pe_i_3__80_,pe_i_3__79_,pe_i_3__78_,pe_i_3__77_,pe_i_3__76_,pe_i_3__75_,
  pe_i_3__74_,pe_i_3__73_,pe_i_3__72_,pe_i_3__71_,pe_i_3__70_,pe_i_3__69_,pe_i_3__68_,
  pe_i_3__67_,pe_i_3__66_,pe_i_3__65_,pe_i_3__64_,pe_i_3__63_,pe_i_3__62_,
  pe_i_3__61_,pe_i_3__60_,pe_i_3__59_,pe_i_3__58_,pe_i_3__57_,pe_i_3__56_,pe_i_3__55_,
  pe_i_3__54_,pe_i_3__53_,pe_i_3__52_,pe_i_3__51_,pe_i_3__50_,pe_i_3__49_,pe_i_3__48_,
  pe_i_3__47_,pe_i_3__46_,pe_i_3__45_,pe_i_3__44_,pe_i_3__43_,pe_i_3__42_,
  pe_i_3__41_,pe_i_3__40_,pe_i_3__39_,pe_i_3__38_,pe_i_3__37_,pe_i_3__36_,pe_i_3__35_,
  pe_i_3__34_,pe_i_3__33_,pe_i_3__32_,pe_i_3__31_,pe_i_3__30_,pe_i_3__29_,pe_i_3__28_,
  pe_i_3__27_,pe_i_3__26_,pe_i_3__25_,pe_i_3__24_,pe_i_3__23_,pe_i_3__22_,
  pe_i_3__21_,pe_i_3__20_,pe_i_3__19_,pe_i_3__18_,pe_i_3__17_,pe_i_3__16_,pe_i_3__15_,
  pe_i_3__14_,pe_i_3__13_,pe_i_3__12_,pe_i_3__11_,pe_i_3__10_,pe_i_3__9_,pe_i_3__8_,
  pe_i_3__7_,pe_i_3__6_,pe_i_3__5_,pe_i_3__4_,pe_i_3__3_,pe_i_3__2_,pe_i_3__1_,
  pe_i_3__0_,pe_i_2__126_,pe_i_2__125_,pe_i_2__124_,pe_i_2__123_,pe_i_2__122_,
  pe_i_2__121_,pe_i_2__120_,pe_i_2__119_,pe_i_2__118_,pe_i_2__117_,pe_i_2__116_,pe_i_2__115_,
  pe_i_2__114_,pe_i_2__113_,pe_i_2__112_,pe_i_2__111_,pe_i_2__110_,pe_i_2__109_,
  pe_i_2__108_,pe_i_2__107_,pe_i_2__106_,pe_i_2__105_,pe_i_2__104_,pe_i_2__103_,
  pe_i_2__102_,pe_i_2__101_,pe_i_2__100_,pe_i_2__99_,pe_i_2__98_,pe_i_2__97_,
  pe_i_2__96_,pe_i_2__95_,pe_i_2__94_,pe_i_2__93_,pe_i_2__92_,pe_i_2__91_,pe_i_2__90_,
  pe_i_2__89_,pe_i_2__88_,pe_i_2__87_,pe_i_2__86_,pe_i_2__85_,pe_i_2__84_,pe_i_2__83_,
  pe_i_2__82_,pe_i_2__81_,pe_i_2__80_,pe_i_2__79_,pe_i_2__78_,pe_i_2__77_,
  pe_i_2__76_,pe_i_2__75_,pe_i_2__74_,pe_i_2__73_,pe_i_2__72_,pe_i_2__71_,pe_i_2__70_,
  pe_i_2__69_,pe_i_2__68_,pe_i_2__67_,pe_i_2__66_,pe_i_2__65_,pe_i_2__64_,pe_i_2__63_,
  pe_i_2__62_,pe_i_2__61_,pe_i_2__60_,pe_i_2__59_,pe_i_2__58_,pe_i_2__57_,
  pe_i_2__56_,pe_i_2__55_,pe_i_2__54_,pe_i_2__53_,pe_i_2__52_,pe_i_2__51_,pe_i_2__50_,
  pe_i_2__49_,pe_i_2__48_,pe_i_2__47_,pe_i_2__46_,pe_i_2__45_,pe_i_2__44_,pe_i_2__43_,
  pe_i_2__42_,pe_i_2__41_,pe_i_2__40_,pe_i_2__39_,pe_i_2__38_,pe_i_2__37_,
  pe_i_2__36_,pe_i_2__35_,pe_i_2__34_,pe_i_2__33_,pe_i_2__32_,pe_i_2__31_,pe_i_2__30_,
  pe_i_2__29_,pe_i_2__28_,pe_i_2__27_,pe_i_2__26_,pe_i_2__25_,pe_i_2__24_,pe_i_2__23_,
  pe_i_2__22_,pe_i_2__21_,pe_i_2__20_,pe_i_2__19_,pe_i_2__18_,pe_i_2__17_,
  pe_i_2__16_,pe_i_2__15_,pe_i_2__14_,pe_i_2__13_,pe_i_2__12_,pe_i_2__11_,pe_i_2__10_,
  pe_i_2__9_,pe_i_2__8_,pe_i_2__7_,pe_i_2__6_,pe_i_2__5_,pe_i_2__4_,pe_i_2__3_,
  pe_i_2__2_,pe_i_2__1_,pe_i_2__0_,pe_i_1__126_,pe_i_1__125_,pe_i_1__124_,pe_i_1__123_,
  pe_i_1__122_,pe_i_1__121_,pe_i_1__120_,pe_i_1__119_,pe_i_1__118_,pe_i_1__117_,
  pe_i_1__116_,pe_i_1__115_,pe_i_1__114_,pe_i_1__113_,pe_i_1__112_,pe_i_1__111_,
  pe_i_1__110_,pe_i_1__109_,pe_i_1__108_,pe_i_1__107_,pe_i_1__106_,pe_i_1__105_,
  pe_i_1__104_,pe_i_1__103_,pe_i_1__102_,pe_i_1__101_,pe_i_1__100_,pe_i_1__99_,pe_i_1__98_,
  pe_i_1__97_,pe_i_1__96_,pe_i_1__95_,pe_i_1__94_,pe_i_1__93_,pe_i_1__92_,
  pe_i_1__91_,pe_i_1__90_,pe_i_1__89_,pe_i_1__88_,pe_i_1__87_,pe_i_1__86_,pe_i_1__85_,
  pe_i_1__84_,pe_i_1__83_,pe_i_1__82_,pe_i_1__81_,pe_i_1__80_,pe_i_1__79_,pe_i_1__78_,
  pe_i_1__77_,pe_i_1__76_,pe_i_1__75_,pe_i_1__74_,pe_i_1__73_,pe_i_1__72_,
  pe_i_1__71_,pe_i_1__70_,pe_i_1__69_,pe_i_1__68_,pe_i_1__67_,pe_i_1__66_,pe_i_1__65_,
  pe_i_1__64_,pe_i_1__63_,pe_i_1__62_,pe_i_1__61_,pe_i_1__60_,pe_i_1__59_,pe_i_1__58_,
  pe_i_1__57_,pe_i_1__56_,pe_i_1__55_,pe_i_1__54_,pe_i_1__53_,pe_i_1__52_,
  pe_i_1__51_,pe_i_1__50_,pe_i_1__49_,pe_i_1__48_,pe_i_1__47_,pe_i_1__46_,pe_i_1__45_,
  pe_i_1__44_,pe_i_1__43_,pe_i_1__42_,pe_i_1__41_,pe_i_1__40_,pe_i_1__39_,pe_i_1__38_,
  pe_i_1__37_,pe_i_1__36_,pe_i_1__35_,pe_i_1__34_,pe_i_1__33_,pe_i_1__32_,
  pe_i_1__31_,pe_i_1__30_,pe_i_1__29_,pe_i_1__28_,pe_i_1__27_,pe_i_1__26_,pe_i_1__25_,
  pe_i_1__24_,pe_i_1__23_,pe_i_1__22_,pe_i_1__21_,pe_i_1__20_,pe_i_1__19_,pe_i_1__18_,
  pe_i_1__17_,pe_i_1__16_,pe_i_1__15_,pe_i_1__14_,pe_i_1__13_,pe_i_1__12_,
  pe_i_1__11_,pe_i_1__10_,pe_i_1__9_,pe_i_1__8_,pe_i_1__7_,pe_i_1__6_,pe_i_1__5_,
  pe_i_1__4_,pe_i_1__3_,pe_i_1__2_,pe_i_1__1_,pe_i_1__0_,N7428,N7429,N7430,N7431,N7432,
  N7433,N7434,N7435,N7436,N7437,N7438,N7439,N7440,N7441,N7442,N7443,N7444,N7445,N7446,
  N7447,N7448,N7449,N7450,N7451,N7452,N7453,N7454,N7455,N7456,N7457,N7458,N7459,
  N7460,N7461,N7462,N7463,N7464,N7465,N7466,N7467,N7468,N7469,N7470,N7471,N7472,
  N7473,N7474,N7475,N7476,N7477,N7478,N7479,N7480,N7481,N7482,N7483,N7484,N7485,N7486,
  N7487,N7488,N7489,N7490,N7491,N7492,N7493,N7494,N7495,N7496,N7497,N7498,N7499,
  N7500,N7501,N7502,N7503,N7504,N7505,N7506,N7507,N7508,N7509,N7510,N7511,N7512,
  N7513,N7514,N7515,N7516,N7517,N7518,N7519,N7520,N7521,N7522,N7523,N7524,N7525,N7526,
  N7527,N7528,N7529,N7530,N7531,N7532,N7533,N7534,N7535,N7536,N7537,N7538,N7539,
  N7540,N7541,N7542,N7543,N7544,N7545,N7546,N7547,N7548,N7549,N7550,N7551,N7552,
  N7553,N7554,N7555,N7556,N7557,N7558,N7559,N7560,N7561,N7562,N7563,N7564,N7565,N7566,
  N7567,N7568,N7569,N7570,N7571,N7572,N7573,N7574,N7575,N7576,N7577,N7578,N7579,
  N7580,N7581,N7582,N7583,N7584,N7585,N7586,N7587,N7588,N7589,N7590,N7591,N7592,
  N7593,N7594,N7595,N7596,N7597,N7598,N7599,N7600,N7601,N7602,N7603,N7604,N7605,N7606,
  N7607,N7608,N7609,N7610,N7611,N7612,N7613,N7614,N7615,N7616,N7617,N7618,N7619,
  N7620,N7621,N7622,N7623,N7624,N7625,N7626,N7627,N7628,N7629,N7630,N7631,N7632,
  N7633,N7634,N7635,N7636,N7637,N7638,N7639,N7640,N7641,N7642,N7643,N7644,N7645,N7646,
  N7647,N7648,N7649,N7650,N7651,N7652,N7653,N7654,N7655,N7656,N7657,N7658,N7659,
  N7660,N7661,N7662,N7663,N7664,N7665,N7666,N7667,N7668,N7669,N7670,N7671,N7672,
  N7673,N7674,N7675,N7676,N7677,N7678,N7679,N7680,N7681,N7682,N7683,N7684,N7685,N7686,
  N7687,N7688,N7689,N7690,N7691,N7692,N7693,N7694,N7695,N7696,N7697,N7698,N7699,
  N7700,N7701,N7702,N7703,N7704,N7705,N7706,N7707,N7708,N7709,N7710,N7711,N7712,
  N7713,N7714,N7715,N7716,N7717,N7718,N7719,N7720,N7721,N7722,N7723,N7724,N7725,N7726,
  N7727,N7728,N7729,N7730,N7731,N7732,N7733,N7734,N7735,N7736,N7737,N7738,N7739,
  N7740,N7741,N7742,N7743,N7744,N7745,N7746,N7747,N7748,N7749,N7750,N7751,N7752,
  N7753,N7754,N7755,N7756,N7757,N7758,N7759,N7760,N7761,N7762,N7763,N7764,N7765,N7766,
  N7767,N7768,N7769,N7770,N7771,N7772,N7773,N7774,N7775,N7776,N7777,N7778,N7779,
  N7780,N7781,N7782,N7783,N7784,N7785,N7786,N7787,N7788,N7789,N7790,N7791,N7792,
  N7793,N7794,N7795,N7796,N7797,N7798,N7799,N7800,N7801,N7802,N7803,N7804,N7805,N7806,
  N7807,N7808,N7809,N7810,N7811,N7812,N7813,N7814,N7815,N7816,N7817,N7818,N7819,
  N7820,N7821,N7822,N7823,N7824,N7825,N7826,N7827,N7828,N7829,N7830,N7831,N7832,
  N7833,N7834,N7835,N7836,N7837,N7838,N7839,N7840,N7841,N7842,N7843,N7844,N7845,N7846,
  N7847,N7848,N7849,N7850,N7851,N7852,N7853,N7854,N7855,N7856,N7857,N7858,N7859,
  N7860,N7861,N7862,N7863,N7864,N7865,N7866,N7867,N7868,N7869,N7870,N7871,N7872,
  N7873,N7874,N7875,N7876,N7877,N7878,N7879,N7880,N7881,N7882,N7883,N7884,N7885,N7886,
  N7887,N7888,N7889,N7890,N7891,N7892,N7893,N7894,N7895,N7896,N7897,N7898,N7899,
  N7900,N7901,N7902,N7903,N7904,N7905,N7906,N7907,N7908,N7909,N7910,N7911,N7912,
  N7913,N7914,N7915,N7916,N7917,N7918,N7919,N7920,N7921,N7922,N7923,N7924,N7925,N7926,
  N7927,N7928,N7929,N7930,N7931,N7932,N7933,N7934,N7935,N7936,N7937,N7938,N7939,
  N7940,N7941,N7942,N7943,N7944,N7945,N7946,N7947,N7948,N7949,N7950,N7951,N7952,
  N7953,N7954,N7955,N7956,N7957,N7958,N7959,N7960,N7961,N7962,N7963,N7964,N7965,N7966,
  N7967,N7968,N7969,N7970,N7971,N7972,N7973,N7974,N7975,N7976,N7977,N7978,N7979,
  N7980,N7981,N7982,N7983,N7984,N7985,N7986,N7987,N7988,N7989,N7990,N7991,N7992,
  N7993,N7994,N7995,N7996,N7997,N7998,N7999,N8000,N8001,N8002,N8003,N8004,N8005,N8006,
  N8007,N8008,N8009,N8010,N8011,N8012,N8013,N8014,N8015,N8016,N8017,N8018,N8019,
  N8020,N8021,N8022,N8023,N8024,N8025,N8026,N8027,N8028,N8029,N8030,N8031,N8032,
  N8033,N8034,N8035,N8036,N8037,N8038,N8039,N8040,N8041,N8042,N8043,N8044,N8045,N8046,
  N8047,N8048,N8049,N8050,N8051,N8052,N8053,N8054,N8055,N8056,N8057,N8058,N8059,
  N8060,N8061,N8062,N8063,N8064,N8065,N8066,N8067,N8068,N8069,N8070,N8071,N8072,
  N8073,N8074,N8075,N8076,N8077,N8078,N8079,N8080,N8081,N8082,N8083,N8084,N8085,N8086,
  N8087,N8088,N8089,N8090,N8091,N8092,N8093,N8094,N8095,N8096,N8097,N8098,N8099,
  N8100,N8101,N8102,N8103,N8104,N8105,N8106,N8107,N8108,N8109,N8110,N8111,N8112,
  N8113,N8114,N8115,N8116,N8117,N8118,N8119,N8120,N8121,N8122,N8123,N8124,N8125,N8126,
  N8127,N8128,N8129,N8130,N8131,N8132,N8133,N8134,N8135,N8136,N8137,N8138,N8139,
  N8140,N8141,N8142,N8143,N8144,N8145,N8146,N8147,N8148,N8149,N8150,N8151,N8152,
  N8153,N8154,N8155,N8156,N8157,N8158,N8159,N8160,N8161,N8162,N8163,N8164,N8165,N8166,
  N8167,N8168,N8169,N8170,N8171,N8172,N8173,N8174,N8175,N8176,N8177,N8178,N8179,
  N8180,N8181,N8182,N8183,N8184,N8185,N8186,N8187,N8188,N8189,N8190,N8191,N8192,
  N8193,N8194,N8195,N8196,N8197,N8198,N8199,N8200,N8201,N8202,N8203,N8204,N8205,N8206,
  N8207,N8208,N8209,N8210,N8211,N8212,N8213,N8214,N8215,N8216,N8217,N8218,N8219,
  N8220,N8221,N8222,N8223,N8224,N8225,N8226,N8227,N8228,N8229,N8230,N8231,N8232,
  N8233,N8234,N8235,N8236,N8237,N8238,N8239,N8240,N8241,N8242,N8243,N8244,N8245,N8246,
  N8247,N8248,N8249,N8250,N8251,N8252,N8253,N8254,N8255,N8256,N8257,N8258,N8259,
  N8260,N8261,N8262,N8263,N8264,N8265,N8266,N8267,N8268,N8269,N8270,N8271,N8272,
  N8273,N8274,N8275,N8276,N8277,N8278,N8279,N8280,N8281,N8282,N8283,N8284,N8285,N8286,
  N8287,N8288,N8289,N8290,N8291,N8292,N8293,N8294,N8295,N8296,N8297,N8298,N8299,
  N8300,N8301,N8302,N8303,N8304,N8305,N8306,N8307,N8308,N8309,N8310,N8311,N8312,
  N8313,N8314,N8315,N8316,N8317,N8318,N8319,N8320,N8321,N8322,N8323,N8324,N8325,N8326,
  N8327,N8328,N8329,N8330,N8331,N8332,N8333,N8334,N8335,N8336,N8337,N8338,N8339,
  N8340,N8341,N8342,N8343,N8344,N8345,N8346,N8347,N8348,N8349,N8350,N8351,N8352,
  N8353,N8354,N8355,N8356,N8357,N8358,N8359,N8360,N8361,N8362,N8363,N8364,N8365,N8366,
  N8367,N8368,N8369,N8370,N8371,N8372,N8373,N8374,N8375,N8376,N8377,N8378,N8379,
  N8380,N8381,N8382,N8383,N8384,N8385,N8386,N8387,N8388,N8389,N8390,N8391,N8392,
  N8393,N8394,N8395,N8396,N8397,N8398,N8399,N8400,N8401,N8402,N8403,N8404,N8405,N8406,
  N8407,N8408,N8409,N8410,N8411,N8412,N8413,N8414,N8415,N8416,N8417,N8418,N8419,
  N8420,N8421,N8422,N8423,N8424,N8425,N8426,N8427,N8428,N8429,N8430,N8431,N8432,
  N8433,N8434,N8435,N8436,N8437,N8438,N8439,N8440,N8441,N8442,N8443,N8444,N8445,N8446,
  N8447,N8448,N8449,N8450,N8451,N8452,N8453,N8454,N8455,N8456,N8457,N8458,N8459,
  N8460,N8461,N8462,N8463,N8464,N8465,N8466,N8467,N8468,N8469,N8470,N8471,N8472,
  N8473,N8474,N8475,N8476,N8477,N8478,N8479,N8480,N8481,N8482,N8483,N8484,N8485,N8486,
  N8487,N8488,N8489,N8490,N8491,N8492,N8493,N8494,N8495,N8496,N8497,N8498,N8499,
  N8500,N8501,N8502,N8503,N8504,N8505,N8506,N8507,N8508,N8509,N8510,N8511,N8512,
  N8513,N8514,N8515,N8516,N8517,N8518,N8519,N8520,N8521,N8522,N8523,N8524,N8525,N8526,
  N8527,N8528,N8529,N8530,N8531,N8532,N8533,N8534,N8535,N8536,N8537,N8538,N8539,
  N8540,N8541,N8542,N8543,N8544,N8545,N8546,N8547,N8548,N8549,N8550,N8551,N8552,
  N8553,N8554,N8555,N8556,N8557,N8558,N8559,N8560,N8561,N8562,N8563,N8564,N8565,N8566,
  N8567,N8568,N8569,N8570,N8571,N8572,N8573,N8574,N8575,N8576,N8577,N8578,N8579,
  N8580,N8581,N8582,N8583,N8584,N8585,N8586,N8587,N8588,N8589,N8590,N8591,N8592,
  N8593,N8594,N8595,N8596,N8597,N8598,N8599,N8600,N8601,N8602,N8603,N8604,N8605,N8606,
  N8607,N8608,N8609,N8610,N8611,N8612,N8613,N8614,N8615,N8616,N8617,N8618,N8619,
  N8620,N8621,N8622,N8623,N8624,N8625,N8626,N8627,N8628,N8629,N8630,N8631,N8632,
  N8633,N8634,N8635,N8636,N8637,N8638,N8639,N8640,N8641,N8642,N8643,N8644,N8645,N8646,
  N8647,N8648,N8649,N8650,N8651,N8652,N8653,N8654,N8655,N8656,N8657,N8658,N8659,
  N8660,N8661,N8662,N8663,N8664,N8665,N8666,N8667,N8668,N8669,N8670,N8671,N8672,
  N8673,N8674,N8675,N8676,N8677,N8678,N8679,N8680,N8681,N8682,N8683,N8684,N8685,N8686,
  N8687,N8688,N8689,N8690,N8691,N8692,N8693,N8694,N8695,N8696,N8697,N8698,N8699,
  N8700,N8701,N8702,N8703,N8704,N8705,N8706,N8707,N8708,N8709,N8710,N8711,N8712,
  N8713,N8714,N8715,N8716,N8717,N8718,N8719,N8720,N8721,N8722,N8723,N8724,N8725,N8726,
  N8727,N8728,N8729,N8730,N8731,N8732,N8733,N8734,N8735,N8736,N8737,N8738,N8739,
  N8740,N8741,N8742,N8743,N8744,N8745,N8746,N8747,N8748,N8749,N8750,N8751,N8752,
  N8753,N8754,N8755,N8756,N8757,N8758,N8759,N8760,N8761,N8762,N8763,N8764,N8765,N8766,
  N8767,N8768,N8769,N8770,N8771,N8772,N8773,N8774,N8775,N8776,N8777,N8778,N8779,
  N8780,N8781,N8782,N8783,N8784,N8785,N8786,N8787,N8788,N8789,N8790,N8791,N8792,
  N8793,N8794,N8795,N8796,N8797,N8798,N8799,N8800,N8801,N8802,N8803,N8804,N8805,N8806,
  N8807,N8808,N8809,N8810,N8811,N8812,N8813,N8814,N8815,N8816,N8817,N8818,N8819,
  N8820,N8821,N8822,N8823,N8824,N8825,N8826,N8827,N8828,N8829,N8830,N8831,N8832,
  N8833,N8834,N8835,N8836,N8837,N8838,N8839,N8840,N8841,N8842,N8843,N8844,N8845,N8846,
  N8847,N8848,N8849,N8850,N8851,N8852,N8853,N8854,N8855,N8856,N8857,N8858,N8859,
  N8860,N8861,N8862,N8863,N8864,N8865,N8866,N8867,N8868,N8869,N8870,N8871,N8872,
  N8873,N8874,N8875,N8876,N8877,N8878,N8879,N8880,N8881,N8882,N8883,N8884,N8885,N8886,
  N8887;
  wire [126:1] mask;

  bsg_priority_encode
  rof2_1__fi3_pe
  (
    .i({ pe_i_1__126_, pe_i_1__125_, pe_i_1__124_, pe_i_1__123_, pe_i_1__122_, pe_i_1__121_, pe_i_1__120_, pe_i_1__119_, pe_i_1__118_, pe_i_1__117_, pe_i_1__116_, pe_i_1__115_, pe_i_1__114_, pe_i_1__113_, pe_i_1__112_, pe_i_1__111_, pe_i_1__110_, pe_i_1__109_, pe_i_1__108_, pe_i_1__107_, pe_i_1__106_, pe_i_1__105_, pe_i_1__104_, pe_i_1__103_, pe_i_1__102_, pe_i_1__101_, pe_i_1__100_, pe_i_1__99_, pe_i_1__98_, pe_i_1__97_, pe_i_1__96_, pe_i_1__95_, pe_i_1__94_, pe_i_1__93_, pe_i_1__92_, pe_i_1__91_, pe_i_1__90_, pe_i_1__89_, pe_i_1__88_, pe_i_1__87_, pe_i_1__86_, pe_i_1__85_, pe_i_1__84_, pe_i_1__83_, pe_i_1__82_, pe_i_1__81_, pe_i_1__80_, pe_i_1__79_, pe_i_1__78_, pe_i_1__77_, pe_i_1__76_, pe_i_1__75_, pe_i_1__74_, pe_i_1__73_, pe_i_1__72_, pe_i_1__71_, pe_i_1__70_, pe_i_1__69_, pe_i_1__68_, pe_i_1__67_, pe_i_1__66_, pe_i_1__65_, pe_i_1__64_, pe_i_1__63_, pe_i_1__62_, pe_i_1__61_, pe_i_1__60_, pe_i_1__59_, pe_i_1__58_, pe_i_1__57_, pe_i_1__56_, pe_i_1__55_, pe_i_1__54_, pe_i_1__53_, pe_i_1__52_, pe_i_1__51_, pe_i_1__50_, pe_i_1__49_, pe_i_1__48_, pe_i_1__47_, pe_i_1__46_, pe_i_1__45_, pe_i_1__44_, pe_i_1__43_, pe_i_1__42_, pe_i_1__41_, pe_i_1__40_, pe_i_1__39_, pe_i_1__38_, pe_i_1__37_, pe_i_1__36_, pe_i_1__35_, pe_i_1__34_, pe_i_1__33_, pe_i_1__32_, pe_i_1__31_, pe_i_1__30_, pe_i_1__29_, pe_i_1__28_, pe_i_1__27_, pe_i_1__26_, pe_i_1__25_, pe_i_1__24_, pe_i_1__23_, pe_i_1__22_, pe_i_1__21_, pe_i_1__20_, pe_i_1__19_, pe_i_1__18_, pe_i_1__17_, pe_i_1__16_, pe_i_1__15_, pe_i_1__14_, pe_i_1__13_, pe_i_1__12_, pe_i_1__11_, pe_i_1__10_, pe_i_1__9_, pe_i_1__8_, pe_i_1__7_, pe_i_1__6_, pe_i_1__5_, pe_i_1__4_, pe_i_1__3_, pe_i_1__2_, pe_i_1__1_, pe_i_1__0_ }),
    .addr_o({ pe_o_1__6_, pe_o_1__5_, pe_o_1__4_, pe_o_1__3_, pe_o_1__2_, pe_o_1__1_, pe_o_1__0_ })
  );

  assign { N7808, N7807, N7806, N7805, N7804, N7803, N7802, N7801, N7800, N7799, N7798, N7797, N7796, N7795, N7794, N7793, N7792, N7791, N7790, N7789, N7788, N7787, N7786, N7785, N7784, N7783, N7782, N7781, N7780, N7779, N7778, N7777, N7776, N7775, N7774, N7773, N7772, N7771, N7770, N7769, N7768, N7767, N7766, N7765, N7764, N7763, N7762, N7761, N7760, N7759, N7758, N7757, N7756, N7755, N7754, N7753, N7752, N7751, N7750, N7749, N7748, N7747, N7746, N7745, N7744, N7743, N7742, N7741, N7740, N7739, N7738, N7737, N7736, N7735, N7734, N7733, N7732, N7731, N7730, N7729, N7728, N7727, N7726, N7725, N7724, N7723, N7722, N7721, N7720, N7719, N7718, N7717, N7716, N7715, N7714, N7713, N7712, N7711, N7710, N7709, N7708, N7707, N7706, N7705, N7704, N7703, N7702, N7701, N7700, N7699, N7698, N7697, N7696, N7695, N7694, N7693, N7692, N7691, N7690, N7689, N7688, N7687, N7686, N7685, N7684, N7683, N7682 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << { pe_o_1__6_, pe_o_1__5_, pe_o_1__4_, pe_o_1__3_, pe_o_1__2_, pe_o_1__1_, pe_o_1__0_ };

  bsg_priority_encode
  rof2_2__fi3_pe
  (
    .i({ pe_i_2__126_, pe_i_2__125_, pe_i_2__124_, pe_i_2__123_, pe_i_2__122_, pe_i_2__121_, pe_i_2__120_, pe_i_2__119_, pe_i_2__118_, pe_i_2__117_, pe_i_2__116_, pe_i_2__115_, pe_i_2__114_, pe_i_2__113_, pe_i_2__112_, pe_i_2__111_, pe_i_2__110_, pe_i_2__109_, pe_i_2__108_, pe_i_2__107_, pe_i_2__106_, pe_i_2__105_, pe_i_2__104_, pe_i_2__103_, pe_i_2__102_, pe_i_2__101_, pe_i_2__100_, pe_i_2__99_, pe_i_2__98_, pe_i_2__97_, pe_i_2__96_, pe_i_2__95_, pe_i_2__94_, pe_i_2__93_, pe_i_2__92_, pe_i_2__91_, pe_i_2__90_, pe_i_2__89_, pe_i_2__88_, pe_i_2__87_, pe_i_2__86_, pe_i_2__85_, pe_i_2__84_, pe_i_2__83_, pe_i_2__82_, pe_i_2__81_, pe_i_2__80_, pe_i_2__79_, pe_i_2__78_, pe_i_2__77_, pe_i_2__76_, pe_i_2__75_, pe_i_2__74_, pe_i_2__73_, pe_i_2__72_, pe_i_2__71_, pe_i_2__70_, pe_i_2__69_, pe_i_2__68_, pe_i_2__67_, pe_i_2__66_, pe_i_2__65_, pe_i_2__64_, pe_i_2__63_, pe_i_2__62_, pe_i_2__61_, pe_i_2__60_, pe_i_2__59_, pe_i_2__58_, pe_i_2__57_, pe_i_2__56_, pe_i_2__55_, pe_i_2__54_, pe_i_2__53_, pe_i_2__52_, pe_i_2__51_, pe_i_2__50_, pe_i_2__49_, pe_i_2__48_, pe_i_2__47_, pe_i_2__46_, pe_i_2__45_, pe_i_2__44_, pe_i_2__43_, pe_i_2__42_, pe_i_2__41_, pe_i_2__40_, pe_i_2__39_, pe_i_2__38_, pe_i_2__37_, pe_i_2__36_, pe_i_2__35_, pe_i_2__34_, pe_i_2__33_, pe_i_2__32_, pe_i_2__31_, pe_i_2__30_, pe_i_2__29_, pe_i_2__28_, pe_i_2__27_, pe_i_2__26_, pe_i_2__25_, pe_i_2__24_, pe_i_2__23_, pe_i_2__22_, pe_i_2__21_, pe_i_2__20_, pe_i_2__19_, pe_i_2__18_, pe_i_2__17_, pe_i_2__16_, pe_i_2__15_, pe_i_2__14_, pe_i_2__13_, pe_i_2__12_, pe_i_2__11_, pe_i_2__10_, pe_i_2__9_, pe_i_2__8_, pe_i_2__7_, pe_i_2__6_, pe_i_2__5_, pe_i_2__4_, pe_i_2__3_, pe_i_2__2_, pe_i_2__1_, pe_i_2__0_ }),
    .addr_o({ pe_o_2__6_, pe_o_2__5_, pe_o_2__4_, pe_o_2__3_, pe_o_2__2_, pe_o_2__1_, pe_o_2__0_ })
  );

  assign { N8062, N8061, N8060, N8059, N8058, N8057, N8056, N8055, N8054, N8053, N8052, N8051, N8050, N8049, N8048, N8047, N8046, N8045, N8044, N8043, N8042, N8041, N8040, N8039, N8038, N8037, N8036, N8035, N8034, N8033, N8032, N8031, N8030, N8029, N8028, N8027, N8026, N8025, N8024, N8023, N8022, N8021, N8020, N8019, N8018, N8017, N8016, N8015, N8014, N8013, N8012, N8011, N8010, N8009, N8008, N8007, N8006, N8005, N8004, N8003, N8002, N8001, N8000, N7999, N7998, N7997, N7996, N7995, N7994, N7993, N7992, N7991, N7990, N7989, N7988, N7987, N7986, N7985, N7984, N7983, N7982, N7981, N7980, N7979, N7978, N7977, N7976, N7975, N7974, N7973, N7972, N7971, N7970, N7969, N7968, N7967, N7966, N7965, N7964, N7963, N7962, N7961, N7960, N7959, N7958, N7957, N7956, N7955, N7954, N7953, N7952, N7951, N7950, N7949, N7948, N7947, N7946, N7945, N7944, N7943, N7942, N7941, N7940, N7939, N7938, N7937, N7936 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << { pe_o_2__6_, pe_o_2__5_, pe_o_2__4_, pe_o_2__3_, pe_o_2__2_, pe_o_2__1_, pe_o_2__0_ };

  bsg_priority_encode
  rof2_3__fi3_pe
  (
    .i({ pe_i_3__126_, pe_i_3__125_, pe_i_3__124_, pe_i_3__123_, pe_i_3__122_, pe_i_3__121_, pe_i_3__120_, pe_i_3__119_, pe_i_3__118_, pe_i_3__117_, pe_i_3__116_, pe_i_3__115_, pe_i_3__114_, pe_i_3__113_, pe_i_3__112_, pe_i_3__111_, pe_i_3__110_, pe_i_3__109_, pe_i_3__108_, pe_i_3__107_, pe_i_3__106_, pe_i_3__105_, pe_i_3__104_, pe_i_3__103_, pe_i_3__102_, pe_i_3__101_, pe_i_3__100_, pe_i_3__99_, pe_i_3__98_, pe_i_3__97_, pe_i_3__96_, pe_i_3__95_, pe_i_3__94_, pe_i_3__93_, pe_i_3__92_, pe_i_3__91_, pe_i_3__90_, pe_i_3__89_, pe_i_3__88_, pe_i_3__87_, pe_i_3__86_, pe_i_3__85_, pe_i_3__84_, pe_i_3__83_, pe_i_3__82_, pe_i_3__81_, pe_i_3__80_, pe_i_3__79_, pe_i_3__78_, pe_i_3__77_, pe_i_3__76_, pe_i_3__75_, pe_i_3__74_, pe_i_3__73_, pe_i_3__72_, pe_i_3__71_, pe_i_3__70_, pe_i_3__69_, pe_i_3__68_, pe_i_3__67_, pe_i_3__66_, pe_i_3__65_, pe_i_3__64_, pe_i_3__63_, pe_i_3__62_, pe_i_3__61_, pe_i_3__60_, pe_i_3__59_, pe_i_3__58_, pe_i_3__57_, pe_i_3__56_, pe_i_3__55_, pe_i_3__54_, pe_i_3__53_, pe_i_3__52_, pe_i_3__51_, pe_i_3__50_, pe_i_3__49_, pe_i_3__48_, pe_i_3__47_, pe_i_3__46_, pe_i_3__45_, pe_i_3__44_, pe_i_3__43_, pe_i_3__42_, pe_i_3__41_, pe_i_3__40_, pe_i_3__39_, pe_i_3__38_, pe_i_3__37_, pe_i_3__36_, pe_i_3__35_, pe_i_3__34_, pe_i_3__33_, pe_i_3__32_, pe_i_3__31_, pe_i_3__30_, pe_i_3__29_, pe_i_3__28_, pe_i_3__27_, pe_i_3__26_, pe_i_3__25_, pe_i_3__24_, pe_i_3__23_, pe_i_3__22_, pe_i_3__21_, pe_i_3__20_, pe_i_3__19_, pe_i_3__18_, pe_i_3__17_, pe_i_3__16_, pe_i_3__15_, pe_i_3__14_, pe_i_3__13_, pe_i_3__12_, pe_i_3__11_, pe_i_3__10_, pe_i_3__9_, pe_i_3__8_, pe_i_3__7_, pe_i_3__6_, pe_i_3__5_, pe_i_3__4_, pe_i_3__3_, pe_i_3__2_, pe_i_3__1_, pe_i_3__0_ }),
    .addr_o({ pe_o_3__6_, pe_o_3__5_, pe_o_3__4_, pe_o_3__3_, pe_o_3__2_, pe_o_3__1_, pe_o_3__0_ })
  );

  assign { N8316, N8315, N8314, N8313, N8312, N8311, N8310, N8309, N8308, N8307, N8306, N8305, N8304, N8303, N8302, N8301, N8300, N8299, N8298, N8297, N8296, N8295, N8294, N8293, N8292, N8291, N8290, N8289, N8288, N8287, N8286, N8285, N8284, N8283, N8282, N8281, N8280, N8279, N8278, N8277, N8276, N8275, N8274, N8273, N8272, N8271, N8270, N8269, N8268, N8267, N8266, N8265, N8264, N8263, N8262, N8261, N8260, N8259, N8258, N8257, N8256, N8255, N8254, N8253, N8252, N8251, N8250, N8249, N8248, N8247, N8246, N8245, N8244, N8243, N8242, N8241, N8240, N8239, N8238, N8237, N8236, N8235, N8234, N8233, N8232, N8231, N8230, N8229, N8228, N8227, N8226, N8225, N8224, N8223, N8222, N8221, N8220, N8219, N8218, N8217, N8216, N8215, N8214, N8213, N8212, N8211, N8210, N8209, N8208, N8207, N8206, N8205, N8204, N8203, N8202, N8201, N8200, N8199, N8198, N8197, N8196, N8195, N8194, N8193, N8192, N8191, N8190 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << { pe_o_3__6_, pe_o_3__5_, pe_o_3__4_, pe_o_3__3_, pe_o_3__2_, pe_o_3__1_, pe_o_3__0_ };

  bsg_priority_encode
  rof2_4__fi3_pe
  (
    .i({ pe_i_4__126_, pe_i_4__125_, pe_i_4__124_, pe_i_4__123_, pe_i_4__122_, pe_i_4__121_, pe_i_4__120_, pe_i_4__119_, pe_i_4__118_, pe_i_4__117_, pe_i_4__116_, pe_i_4__115_, pe_i_4__114_, pe_i_4__113_, pe_i_4__112_, pe_i_4__111_, pe_i_4__110_, pe_i_4__109_, pe_i_4__108_, pe_i_4__107_, pe_i_4__106_, pe_i_4__105_, pe_i_4__104_, pe_i_4__103_, pe_i_4__102_, pe_i_4__101_, pe_i_4__100_, pe_i_4__99_, pe_i_4__98_, pe_i_4__97_, pe_i_4__96_, pe_i_4__95_, pe_i_4__94_, pe_i_4__93_, pe_i_4__92_, pe_i_4__91_, pe_i_4__90_, pe_i_4__89_, pe_i_4__88_, pe_i_4__87_, pe_i_4__86_, pe_i_4__85_, pe_i_4__84_, pe_i_4__83_, pe_i_4__82_, pe_i_4__81_, pe_i_4__80_, pe_i_4__79_, pe_i_4__78_, pe_i_4__77_, pe_i_4__76_, pe_i_4__75_, pe_i_4__74_, pe_i_4__73_, pe_i_4__72_, pe_i_4__71_, pe_i_4__70_, pe_i_4__69_, pe_i_4__68_, pe_i_4__67_, pe_i_4__66_, pe_i_4__65_, pe_i_4__64_, pe_i_4__63_, pe_i_4__62_, pe_i_4__61_, pe_i_4__60_, pe_i_4__59_, pe_i_4__58_, pe_i_4__57_, pe_i_4__56_, pe_i_4__55_, pe_i_4__54_, pe_i_4__53_, pe_i_4__52_, pe_i_4__51_, pe_i_4__50_, pe_i_4__49_, pe_i_4__48_, pe_i_4__47_, pe_i_4__46_, pe_i_4__45_, pe_i_4__44_, pe_i_4__43_, pe_i_4__42_, pe_i_4__41_, pe_i_4__40_, pe_i_4__39_, pe_i_4__38_, pe_i_4__37_, pe_i_4__36_, pe_i_4__35_, pe_i_4__34_, pe_i_4__33_, pe_i_4__32_, pe_i_4__31_, pe_i_4__30_, pe_i_4__29_, pe_i_4__28_, pe_i_4__27_, pe_i_4__26_, pe_i_4__25_, pe_i_4__24_, pe_i_4__23_, pe_i_4__22_, pe_i_4__21_, pe_i_4__20_, pe_i_4__19_, pe_i_4__18_, pe_i_4__17_, pe_i_4__16_, pe_i_4__15_, pe_i_4__14_, pe_i_4__13_, pe_i_4__12_, pe_i_4__11_, pe_i_4__10_, pe_i_4__9_, pe_i_4__8_, pe_i_4__7_, pe_i_4__6_, pe_i_4__5_, pe_i_4__4_, pe_i_4__3_, pe_i_4__2_, pe_i_4__1_, pe_i_4__0_ }),
    .addr_o({ pe_o_4__6_, pe_o_4__5_, pe_o_4__4_, pe_o_4__3_, pe_o_4__2_, pe_o_4__1_, pe_o_4__0_ })
  );

  assign { N8570, N8569, N8568, N8567, N8566, N8565, N8564, N8563, N8562, N8561, N8560, N8559, N8558, N8557, N8556, N8555, N8554, N8553, N8552, N8551, N8550, N8549, N8548, N8547, N8546, N8545, N8544, N8543, N8542, N8541, N8540, N8539, N8538, N8537, N8536, N8535, N8534, N8533, N8532, N8531, N8530, N8529, N8528, N8527, N8526, N8525, N8524, N8523, N8522, N8521, N8520, N8519, N8518, N8517, N8516, N8515, N8514, N8513, N8512, N8511, N8510, N8509, N8508, N8507, N8506, N8505, N8504, N8503, N8502, N8501, N8500, N8499, N8498, N8497, N8496, N8495, N8494, N8493, N8492, N8491, N8490, N8489, N8488, N8487, N8486, N8485, N8484, N8483, N8482, N8481, N8480, N8479, N8478, N8477, N8476, N8475, N8474, N8473, N8472, N8471, N8470, N8469, N8468, N8467, N8466, N8465, N8464, N8463, N8462, N8461, N8460, N8459, N8458, N8457, N8456, N8455, N8454, N8453, N8452, N8451, N8450, N8449, N8448, N8447, N8446, N8445, N8444 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << { pe_o_4__6_, pe_o_4__5_, pe_o_4__4_, pe_o_4__3_, pe_o_4__2_, pe_o_4__1_, pe_o_4__0_ };

  bsg_priority_encode
  rof2_5__fi3_pe
  (
    .i({ pe_i_5__126_, pe_i_5__125_, pe_i_5__124_, pe_i_5__123_, pe_i_5__122_, pe_i_5__121_, pe_i_5__120_, pe_i_5__119_, pe_i_5__118_, pe_i_5__117_, pe_i_5__116_, pe_i_5__115_, pe_i_5__114_, pe_i_5__113_, pe_i_5__112_, pe_i_5__111_, pe_i_5__110_, pe_i_5__109_, pe_i_5__108_, pe_i_5__107_, pe_i_5__106_, pe_i_5__105_, pe_i_5__104_, pe_i_5__103_, pe_i_5__102_, pe_i_5__101_, pe_i_5__100_, pe_i_5__99_, pe_i_5__98_, pe_i_5__97_, pe_i_5__96_, pe_i_5__95_, pe_i_5__94_, pe_i_5__93_, pe_i_5__92_, pe_i_5__91_, pe_i_5__90_, pe_i_5__89_, pe_i_5__88_, pe_i_5__87_, pe_i_5__86_, pe_i_5__85_, pe_i_5__84_, pe_i_5__83_, pe_i_5__82_, pe_i_5__81_, pe_i_5__80_, pe_i_5__79_, pe_i_5__78_, pe_i_5__77_, pe_i_5__76_, pe_i_5__75_, pe_i_5__74_, pe_i_5__73_, pe_i_5__72_, pe_i_5__71_, pe_i_5__70_, pe_i_5__69_, pe_i_5__68_, pe_i_5__67_, pe_i_5__66_, pe_i_5__65_, pe_i_5__64_, pe_i_5__63_, pe_i_5__62_, pe_i_5__61_, pe_i_5__60_, pe_i_5__59_, pe_i_5__58_, pe_i_5__57_, pe_i_5__56_, pe_i_5__55_, pe_i_5__54_, pe_i_5__53_, pe_i_5__52_, pe_i_5__51_, pe_i_5__50_, pe_i_5__49_, pe_i_5__48_, pe_i_5__47_, pe_i_5__46_, pe_i_5__45_, pe_i_5__44_, pe_i_5__43_, pe_i_5__42_, pe_i_5__41_, pe_i_5__40_, pe_i_5__39_, pe_i_5__38_, pe_i_5__37_, pe_i_5__36_, pe_i_5__35_, pe_i_5__34_, pe_i_5__33_, pe_i_5__32_, pe_i_5__31_, pe_i_5__30_, pe_i_5__29_, pe_i_5__28_, pe_i_5__27_, pe_i_5__26_, pe_i_5__25_, pe_i_5__24_, pe_i_5__23_, pe_i_5__22_, pe_i_5__21_, pe_i_5__20_, pe_i_5__19_, pe_i_5__18_, pe_i_5__17_, pe_i_5__16_, pe_i_5__15_, pe_i_5__14_, pe_i_5__13_, pe_i_5__12_, pe_i_5__11_, pe_i_5__10_, pe_i_5__9_, pe_i_5__8_, pe_i_5__7_, pe_i_5__6_, pe_i_5__5_, pe_i_5__4_, pe_i_5__3_, pe_i_5__2_, pe_i_5__1_, pe_i_5__0_ }),
    .addr_o({ pe_o_5__6_, pe_o_5__5_, pe_o_5__4_, pe_o_5__3_, pe_o_5__2_, pe_o_5__1_, pe_o_5__0_ })
  );

  assign { N8824, N8823, N8822, N8821, N8820, N8819, N8818, N8817, N8816, N8815, N8814, N8813, N8812, N8811, N8810, N8809, N8808, N8807, N8806, N8805, N8804, N8803, N8802, N8801, N8800, N8799, N8798, N8797, N8796, N8795, N8794, N8793, N8792, N8791, N8790, N8789, N8788, N8787, N8786, N8785, N8784, N8783, N8782, N8781, N8780, N8779, N8778, N8777, N8776, N8775, N8774, N8773, N8772, N8771, N8770, N8769, N8768, N8767, N8766, N8765, N8764, N8763, N8762, N8761, N8760, N8759, N8758, N8757, N8756, N8755, N8754, N8753, N8752, N8751, N8750, N8749, N8748, N8747, N8746, N8745, N8744, N8743, N8742, N8741, N8740, N8739, N8738, N8737, N8736, N8735, N8734, N8733, N8732, N8731, N8730, N8729, N8728, N8727, N8726, N8725, N8724, N8723, N8722, N8721, N8720, N8719, N8718, N8717, N8716, N8715, N8714, N8713, N8712, N8711, N8710, N8709, N8708, N8707, N8706, N8705, N8704, N8703, N8702, N8701, N8700, N8699, N8698 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << { pe_o_5__6_, pe_o_5__5_, pe_o_5__4_, pe_o_5__3_, pe_o_5__2_, pe_o_5__1_, pe_o_5__0_ };

  bsg_priority_encode
  rof2_6__fi3_pe
  (
    .i({ pe_i_6__126_, pe_i_6__125_, pe_i_6__124_, pe_i_6__123_, pe_i_6__122_, pe_i_6__121_, pe_i_6__120_, pe_i_6__119_, pe_i_6__118_, pe_i_6__117_, pe_i_6__116_, pe_i_6__115_, pe_i_6__114_, pe_i_6__113_, pe_i_6__112_, pe_i_6__111_, pe_i_6__110_, pe_i_6__109_, pe_i_6__108_, pe_i_6__107_, pe_i_6__106_, pe_i_6__105_, pe_i_6__104_, pe_i_6__103_, pe_i_6__102_, pe_i_6__101_, pe_i_6__100_, pe_i_6__99_, pe_i_6__98_, pe_i_6__97_, pe_i_6__96_, pe_i_6__95_, pe_i_6__94_, pe_i_6__93_, pe_i_6__92_, pe_i_6__91_, pe_i_6__90_, pe_i_6__89_, pe_i_6__88_, pe_i_6__87_, pe_i_6__86_, pe_i_6__85_, pe_i_6__84_, pe_i_6__83_, pe_i_6__82_, pe_i_6__81_, pe_i_6__80_, pe_i_6__79_, pe_i_6__78_, pe_i_6__77_, pe_i_6__76_, pe_i_6__75_, pe_i_6__74_, pe_i_6__73_, pe_i_6__72_, pe_i_6__71_, pe_i_6__70_, pe_i_6__69_, pe_i_6__68_, pe_i_6__67_, pe_i_6__66_, pe_i_6__65_, pe_i_6__64_, pe_i_6__63_, pe_i_6__62_, pe_i_6__61_, pe_i_6__60_, pe_i_6__59_, pe_i_6__58_, pe_i_6__57_, pe_i_6__56_, pe_i_6__55_, pe_i_6__54_, pe_i_6__53_, pe_i_6__52_, pe_i_6__51_, pe_i_6__50_, pe_i_6__49_, pe_i_6__48_, pe_i_6__47_, pe_i_6__46_, pe_i_6__45_, pe_i_6__44_, pe_i_6__43_, pe_i_6__42_, pe_i_6__41_, pe_i_6__40_, pe_i_6__39_, pe_i_6__38_, pe_i_6__37_, pe_i_6__36_, pe_i_6__35_, pe_i_6__34_, pe_i_6__33_, pe_i_6__32_, pe_i_6__31_, pe_i_6__30_, pe_i_6__29_, pe_i_6__28_, pe_i_6__27_, pe_i_6__26_, pe_i_6__25_, pe_i_6__24_, pe_i_6__23_, pe_i_6__22_, pe_i_6__21_, pe_i_6__20_, pe_i_6__19_, pe_i_6__18_, pe_i_6__17_, pe_i_6__16_, pe_i_6__15_, pe_i_6__14_, pe_i_6__13_, pe_i_6__12_, pe_i_6__11_, pe_i_6__10_, pe_i_6__9_, pe_i_6__8_, pe_i_6__7_, pe_i_6__6_, pe_i_6__5_, pe_i_6__4_, pe_i_6__3_, pe_i_6__2_, pe_i_6__1_, pe_i_6__0_ }),
    .addr_o({ pe_o_6__6_, pe_o_6__5_, pe_o_6__4_, pe_o_6__3_, pe_o_6__2_, pe_o_6__1_, pe_o_6__0_ })
  );

  assign N0 = N5 & N6;
  assign N1 = N0 & N7;
  assign N2 = N1 & N8;
  assign N3 = N2 & N9;
  assign N4 = N3 & N10;
  assign N7428 = N4 & N11;
  assign N5 = ~pe_o_1__6_;
  assign N6 = ~pe_o_1__5_;
  assign N7 = ~pe_o_1__4_;
  assign N8 = ~pe_o_1__3_;
  assign N9 = ~pe_o_1__2_;
  assign N10 = ~pe_o_1__0_;
  assign N11 = ~pe_o_1__1_;
  assign N12 = pe_o_1__6_ & N17;
  assign N13 = N12 & N18;
  assign N14 = N13 & N19;
  assign N15 = N14 & N20;
  assign N16 = N15 & N21;
  assign N7429 = N16 & N22;
  assign N17 = ~pe_o_1__5_;
  assign N18 = ~pe_o_1__4_;
  assign N19 = ~pe_o_1__3_;
  assign N20 = ~pe_o_1__2_;
  assign N21 = ~pe_o_1__0_;
  assign N22 = ~pe_o_1__1_;
  assign N23 = N28 & N29;
  assign N24 = N23 & N30;
  assign N25 = N24 & N31;
  assign N26 = N25 & N32;
  assign N27 = N26 & pe_o_1__0_;
  assign N7430 = N27 & N33;
  assign N28 = ~pe_o_1__6_;
  assign N29 = ~pe_o_1__5_;
  assign N30 = ~pe_o_1__4_;
  assign N31 = ~pe_o_1__3_;
  assign N32 = ~pe_o_1__2_;
  assign N33 = ~pe_o_1__1_;
  assign N34 = N39 & N40;
  assign N35 = N34 & N41;
  assign N36 = N35 & N42;
  assign N37 = N36 & N43;
  assign N38 = N37 & N44;
  assign N7432 = N38 & pe_o_1__1_;
  assign N39 = ~pe_o_1__6_;
  assign N40 = ~pe_o_1__5_;
  assign N41 = ~pe_o_1__4_;
  assign N42 = ~pe_o_1__3_;
  assign N43 = ~pe_o_1__2_;
  assign N44 = ~pe_o_1__0_;
  assign N45 = N50 & N51;
  assign N46 = N45 & N52;
  assign N47 = N46 & N53;
  assign N48 = N47 & N54;
  assign N49 = N48 & pe_o_1__0_;
  assign N7434 = N49 & pe_o_1__1_;
  assign N50 = ~pe_o_1__6_;
  assign N51 = ~pe_o_1__5_;
  assign N52 = ~pe_o_1__4_;
  assign N53 = ~pe_o_1__3_;
  assign N54 = ~pe_o_1__2_;
  assign N55 = N60 & N61;
  assign N56 = N55 & N62;
  assign N57 = N56 & N63;
  assign N58 = N57 & pe_o_1__2_;
  assign N59 = N58 & N64;
  assign N7436 = N59 & N65;
  assign N60 = ~pe_o_1__6_;
  assign N61 = ~pe_o_1__5_;
  assign N62 = ~pe_o_1__4_;
  assign N63 = ~pe_o_1__3_;
  assign N64 = ~pe_o_1__0_;
  assign N65 = ~pe_o_1__1_;
  assign N66 = N71 & N72;
  assign N67 = N66 & N73;
  assign N68 = N67 & N74;
  assign N69 = N68 & pe_o_1__2_;
  assign N70 = N69 & pe_o_1__0_;
  assign N7438 = N70 & N75;
  assign N71 = ~pe_o_1__6_;
  assign N72 = ~pe_o_1__5_;
  assign N73 = ~pe_o_1__4_;
  assign N74 = ~pe_o_1__3_;
  assign N75 = ~pe_o_1__1_;
  assign N76 = N81 & N82;
  assign N77 = N76 & N83;
  assign N78 = N77 & N84;
  assign N79 = N78 & pe_o_1__2_;
  assign N80 = N79 & N85;
  assign N7440 = N80 & pe_o_1__1_;
  assign N81 = ~pe_o_1__6_;
  assign N82 = ~pe_o_1__5_;
  assign N83 = ~pe_o_1__4_;
  assign N84 = ~pe_o_1__3_;
  assign N85 = ~pe_o_1__0_;
  assign N86 = N91 & N92;
  assign N87 = N86 & N93;
  assign N88 = N87 & N94;
  assign N89 = N88 & pe_o_1__2_;
  assign N90 = N89 & pe_o_1__0_;
  assign N7442 = N90 & pe_o_1__1_;
  assign N91 = ~pe_o_1__6_;
  assign N92 = ~pe_o_1__5_;
  assign N93 = ~pe_o_1__4_;
  assign N94 = ~pe_o_1__3_;
  assign N95 = N100 & N101;
  assign N96 = N95 & N102;
  assign N97 = N96 & pe_o_1__3_;
  assign N98 = N97 & N103;
  assign N99 = N98 & N104;
  assign N7444 = N99 & N105;
  assign N100 = ~pe_o_1__6_;
  assign N101 = ~pe_o_1__5_;
  assign N102 = ~pe_o_1__4_;
  assign N103 = ~pe_o_1__2_;
  assign N104 = ~pe_o_1__0_;
  assign N105 = ~pe_o_1__1_;
  assign N106 = N111 & N112;
  assign N107 = N106 & N113;
  assign N108 = N107 & pe_o_1__3_;
  assign N109 = N108 & N114;
  assign N110 = N109 & pe_o_1__0_;
  assign N7446 = N110 & N115;
  assign N111 = ~pe_o_1__6_;
  assign N112 = ~pe_o_1__5_;
  assign N113 = ~pe_o_1__4_;
  assign N114 = ~pe_o_1__2_;
  assign N115 = ~pe_o_1__1_;
  assign N116 = N121 & N122;
  assign N117 = N116 & N123;
  assign N118 = N117 & pe_o_1__3_;
  assign N119 = N118 & N124;
  assign N120 = N119 & N125;
  assign N7448 = N120 & pe_o_1__1_;
  assign N121 = ~pe_o_1__6_;
  assign N122 = ~pe_o_1__5_;
  assign N123 = ~pe_o_1__4_;
  assign N124 = ~pe_o_1__2_;
  assign N125 = ~pe_o_1__0_;
  assign N126 = N131 & N132;
  assign N127 = N126 & N133;
  assign N128 = N127 & pe_o_1__3_;
  assign N129 = N128 & N134;
  assign N130 = N129 & pe_o_1__0_;
  assign N7450 = N130 & pe_o_1__1_;
  assign N131 = ~pe_o_1__6_;
  assign N132 = ~pe_o_1__5_;
  assign N133 = ~pe_o_1__4_;
  assign N134 = ~pe_o_1__2_;
  assign N135 = N140 & N141;
  assign N136 = N135 & N142;
  assign N137 = N136 & pe_o_1__3_;
  assign N138 = N137 & pe_o_1__2_;
  assign N139 = N138 & N143;
  assign N7452 = N139 & N144;
  assign N140 = ~pe_o_1__6_;
  assign N141 = ~pe_o_1__5_;
  assign N142 = ~pe_o_1__4_;
  assign N143 = ~pe_o_1__0_;
  assign N144 = ~pe_o_1__1_;
  assign N145 = N150 & N151;
  assign N146 = N145 & N152;
  assign N147 = N146 & pe_o_1__3_;
  assign N148 = N147 & pe_o_1__2_;
  assign N149 = N148 & pe_o_1__0_;
  assign N7454 = N149 & N153;
  assign N150 = ~pe_o_1__6_;
  assign N151 = ~pe_o_1__5_;
  assign N152 = ~pe_o_1__4_;
  assign N153 = ~pe_o_1__1_;
  assign N154 = N159 & N160;
  assign N155 = N154 & N161;
  assign N156 = N155 & pe_o_1__3_;
  assign N157 = N156 & pe_o_1__2_;
  assign N158 = N157 & N162;
  assign N7456 = N158 & pe_o_1__1_;
  assign N159 = ~pe_o_1__6_;
  assign N160 = ~pe_o_1__5_;
  assign N161 = ~pe_o_1__4_;
  assign N162 = ~pe_o_1__0_;
  assign N163 = N168 & N169;
  assign N164 = N163 & N170;
  assign N165 = N164 & pe_o_1__3_;
  assign N166 = N165 & pe_o_1__2_;
  assign N167 = N166 & pe_o_1__0_;
  assign N7458 = N167 & pe_o_1__1_;
  assign N168 = ~pe_o_1__6_;
  assign N169 = ~pe_o_1__5_;
  assign N170 = ~pe_o_1__4_;
  assign N171 = N176 & N177;
  assign N172 = N171 & pe_o_1__4_;
  assign N173 = N172 & N178;
  assign N174 = N173 & N179;
  assign N175 = N174 & N180;
  assign N7460 = N175 & N181;
  assign N176 = ~pe_o_1__6_;
  assign N177 = ~pe_o_1__5_;
  assign N178 = ~pe_o_1__3_;
  assign N179 = ~pe_o_1__2_;
  assign N180 = ~pe_o_1__0_;
  assign N181 = ~pe_o_1__1_;
  assign N182 = N187 & N188;
  assign N183 = N182 & pe_o_1__4_;
  assign N184 = N183 & N189;
  assign N185 = N184 & N190;
  assign N186 = N185 & pe_o_1__0_;
  assign N7462 = N186 & N191;
  assign N187 = ~pe_o_1__6_;
  assign N188 = ~pe_o_1__5_;
  assign N189 = ~pe_o_1__3_;
  assign N190 = ~pe_o_1__2_;
  assign N191 = ~pe_o_1__1_;
  assign N192 = N197 & N198;
  assign N193 = N192 & pe_o_1__4_;
  assign N194 = N193 & N199;
  assign N195 = N194 & N200;
  assign N196 = N195 & N201;
  assign N7464 = N196 & pe_o_1__1_;
  assign N197 = ~pe_o_1__6_;
  assign N198 = ~pe_o_1__5_;
  assign N199 = ~pe_o_1__3_;
  assign N200 = ~pe_o_1__2_;
  assign N201 = ~pe_o_1__0_;
  assign N202 = N207 & N208;
  assign N203 = N202 & pe_o_1__4_;
  assign N204 = N203 & N209;
  assign N205 = N204 & N210;
  assign N206 = N205 & pe_o_1__0_;
  assign N7466 = N206 & pe_o_1__1_;
  assign N207 = ~pe_o_1__6_;
  assign N208 = ~pe_o_1__5_;
  assign N209 = ~pe_o_1__3_;
  assign N210 = ~pe_o_1__2_;
  assign N211 = N216 & N217;
  assign N212 = N211 & pe_o_1__4_;
  assign N213 = N212 & N218;
  assign N214 = N213 & pe_o_1__2_;
  assign N215 = N214 & N219;
  assign N7468 = N215 & N220;
  assign N216 = ~pe_o_1__6_;
  assign N217 = ~pe_o_1__5_;
  assign N218 = ~pe_o_1__3_;
  assign N219 = ~pe_o_1__0_;
  assign N220 = ~pe_o_1__1_;
  assign N221 = N226 & N227;
  assign N222 = N221 & pe_o_1__4_;
  assign N223 = N222 & N228;
  assign N224 = N223 & pe_o_1__2_;
  assign N225 = N224 & pe_o_1__0_;
  assign N7470 = N225 & N229;
  assign N226 = ~pe_o_1__6_;
  assign N227 = ~pe_o_1__5_;
  assign N228 = ~pe_o_1__3_;
  assign N229 = ~pe_o_1__1_;
  assign N230 = N235 & N236;
  assign N231 = N230 & pe_o_1__4_;
  assign N232 = N231 & N237;
  assign N233 = N232 & pe_o_1__2_;
  assign N234 = N233 & N238;
  assign N7472 = N234 & pe_o_1__1_;
  assign N235 = ~pe_o_1__6_;
  assign N236 = ~pe_o_1__5_;
  assign N237 = ~pe_o_1__3_;
  assign N238 = ~pe_o_1__0_;
  assign N239 = N244 & N245;
  assign N240 = N239 & pe_o_1__4_;
  assign N241 = N240 & N246;
  assign N242 = N241 & pe_o_1__2_;
  assign N243 = N242 & pe_o_1__0_;
  assign N7474 = N243 & pe_o_1__1_;
  assign N244 = ~pe_o_1__6_;
  assign N245 = ~pe_o_1__5_;
  assign N246 = ~pe_o_1__3_;
  assign N247 = N252 & N253;
  assign N248 = N247 & pe_o_1__4_;
  assign N249 = N248 & pe_o_1__3_;
  assign N250 = N249 & N254;
  assign N251 = N250 & N255;
  assign N7476 = N251 & N256;
  assign N252 = ~pe_o_1__6_;
  assign N253 = ~pe_o_1__5_;
  assign N254 = ~pe_o_1__2_;
  assign N255 = ~pe_o_1__0_;
  assign N256 = ~pe_o_1__1_;
  assign N257 = N262 & N263;
  assign N258 = N257 & pe_o_1__4_;
  assign N259 = N258 & pe_o_1__3_;
  assign N260 = N259 & N264;
  assign N261 = N260 & pe_o_1__0_;
  assign N7478 = N261 & N265;
  assign N262 = ~pe_o_1__6_;
  assign N263 = ~pe_o_1__5_;
  assign N264 = ~pe_o_1__2_;
  assign N265 = ~pe_o_1__1_;
  assign N266 = N271 & N272;
  assign N267 = N266 & pe_o_1__4_;
  assign N268 = N267 & pe_o_1__3_;
  assign N269 = N268 & N273;
  assign N270 = N269 & N274;
  assign N7480 = N270 & pe_o_1__1_;
  assign N271 = ~pe_o_1__6_;
  assign N272 = ~pe_o_1__5_;
  assign N273 = ~pe_o_1__2_;
  assign N274 = ~pe_o_1__0_;
  assign N275 = N280 & N281;
  assign N276 = N275 & pe_o_1__4_;
  assign N277 = N276 & pe_o_1__3_;
  assign N278 = N277 & N282;
  assign N279 = N278 & pe_o_1__0_;
  assign N7482 = N279 & pe_o_1__1_;
  assign N280 = ~pe_o_1__6_;
  assign N281 = ~pe_o_1__5_;
  assign N282 = ~pe_o_1__2_;
  assign N283 = N288 & N289;
  assign N284 = N283 & pe_o_1__4_;
  assign N285 = N284 & pe_o_1__3_;
  assign N286 = N285 & pe_o_1__2_;
  assign N287 = N286 & N290;
  assign N7484 = N287 & N291;
  assign N288 = ~pe_o_1__6_;
  assign N289 = ~pe_o_1__5_;
  assign N290 = ~pe_o_1__0_;
  assign N291 = ~pe_o_1__1_;
  assign N292 = N297 & N298;
  assign N293 = N292 & pe_o_1__4_;
  assign N294 = N293 & pe_o_1__3_;
  assign N295 = N294 & pe_o_1__2_;
  assign N296 = N295 & pe_o_1__0_;
  assign N7486 = N296 & N299;
  assign N297 = ~pe_o_1__6_;
  assign N298 = ~pe_o_1__5_;
  assign N299 = ~pe_o_1__1_;
  assign N300 = N305 & N306;
  assign N301 = N300 & pe_o_1__4_;
  assign N302 = N301 & pe_o_1__3_;
  assign N303 = N302 & pe_o_1__2_;
  assign N304 = N303 & N307;
  assign N7488 = N304 & pe_o_1__1_;
  assign N305 = ~pe_o_1__6_;
  assign N306 = ~pe_o_1__5_;
  assign N307 = ~pe_o_1__0_;
  assign N308 = N313 & N314;
  assign N309 = N308 & pe_o_1__4_;
  assign N310 = N309 & pe_o_1__3_;
  assign N311 = N310 & pe_o_1__2_;
  assign N312 = N311 & pe_o_1__0_;
  assign N7490 = N312 & pe_o_1__1_;
  assign N313 = ~pe_o_1__6_;
  assign N314 = ~pe_o_1__5_;
  assign N315 = N320 & pe_o_1__5_;
  assign N316 = N315 & N321;
  assign N317 = N316 & N322;
  assign N318 = N317 & N323;
  assign N319 = N318 & N324;
  assign N7492 = N319 & N325;
  assign N320 = ~pe_o_1__6_;
  assign N321 = ~pe_o_1__4_;
  assign N322 = ~pe_o_1__3_;
  assign N323 = ~pe_o_1__2_;
  assign N324 = ~pe_o_1__0_;
  assign N325 = ~pe_o_1__1_;
  assign N326 = N331 & pe_o_1__5_;
  assign N327 = N326 & N332;
  assign N328 = N327 & N333;
  assign N329 = N328 & N334;
  assign N330 = N329 & pe_o_1__0_;
  assign N7494 = N330 & N335;
  assign N331 = ~pe_o_1__6_;
  assign N332 = ~pe_o_1__4_;
  assign N333 = ~pe_o_1__3_;
  assign N334 = ~pe_o_1__2_;
  assign N335 = ~pe_o_1__1_;
  assign N336 = N341 & pe_o_1__5_;
  assign N337 = N336 & N342;
  assign N338 = N337 & N343;
  assign N339 = N338 & N344;
  assign N340 = N339 & N345;
  assign N7496 = N340 & pe_o_1__1_;
  assign N341 = ~pe_o_1__6_;
  assign N342 = ~pe_o_1__4_;
  assign N343 = ~pe_o_1__3_;
  assign N344 = ~pe_o_1__2_;
  assign N345 = ~pe_o_1__0_;
  assign N346 = N351 & pe_o_1__5_;
  assign N347 = N346 & N352;
  assign N348 = N347 & N353;
  assign N349 = N348 & N354;
  assign N350 = N349 & pe_o_1__0_;
  assign N7498 = N350 & pe_o_1__1_;
  assign N351 = ~pe_o_1__6_;
  assign N352 = ~pe_o_1__4_;
  assign N353 = ~pe_o_1__3_;
  assign N354 = ~pe_o_1__2_;
  assign N355 = N360 & pe_o_1__5_;
  assign N356 = N355 & N361;
  assign N357 = N356 & N362;
  assign N358 = N357 & pe_o_1__2_;
  assign N359 = N358 & N363;
  assign N7500 = N359 & N364;
  assign N360 = ~pe_o_1__6_;
  assign N361 = ~pe_o_1__4_;
  assign N362 = ~pe_o_1__3_;
  assign N363 = ~pe_o_1__0_;
  assign N364 = ~pe_o_1__1_;
  assign N365 = N370 & pe_o_1__5_;
  assign N366 = N365 & N371;
  assign N367 = N366 & N372;
  assign N368 = N367 & pe_o_1__2_;
  assign N369 = N368 & pe_o_1__0_;
  assign N7502 = N369 & N373;
  assign N370 = ~pe_o_1__6_;
  assign N371 = ~pe_o_1__4_;
  assign N372 = ~pe_o_1__3_;
  assign N373 = ~pe_o_1__1_;
  assign N374 = N379 & pe_o_1__5_;
  assign N375 = N374 & N380;
  assign N376 = N375 & N381;
  assign N377 = N376 & pe_o_1__2_;
  assign N378 = N377 & N382;
  assign N7504 = N378 & pe_o_1__1_;
  assign N379 = ~pe_o_1__6_;
  assign N380 = ~pe_o_1__4_;
  assign N381 = ~pe_o_1__3_;
  assign N382 = ~pe_o_1__0_;
  assign N383 = N388 & pe_o_1__5_;
  assign N384 = N383 & N389;
  assign N385 = N384 & N390;
  assign N386 = N385 & pe_o_1__2_;
  assign N387 = N386 & pe_o_1__0_;
  assign N7506 = N387 & pe_o_1__1_;
  assign N388 = ~pe_o_1__6_;
  assign N389 = ~pe_o_1__4_;
  assign N390 = ~pe_o_1__3_;
  assign N391 = N396 & pe_o_1__5_;
  assign N392 = N391 & N397;
  assign N393 = N392 & pe_o_1__3_;
  assign N394 = N393 & N398;
  assign N395 = N394 & N399;
  assign N7508 = N395 & N400;
  assign N396 = ~pe_o_1__6_;
  assign N397 = ~pe_o_1__4_;
  assign N398 = ~pe_o_1__2_;
  assign N399 = ~pe_o_1__0_;
  assign N400 = ~pe_o_1__1_;
  assign N401 = N406 & pe_o_1__5_;
  assign N402 = N401 & N407;
  assign N403 = N402 & pe_o_1__3_;
  assign N404 = N403 & N408;
  assign N405 = N404 & pe_o_1__0_;
  assign N7510 = N405 & N409;
  assign N406 = ~pe_o_1__6_;
  assign N407 = ~pe_o_1__4_;
  assign N408 = ~pe_o_1__2_;
  assign N409 = ~pe_o_1__1_;
  assign N410 = N415 & pe_o_1__5_;
  assign N411 = N410 & N416;
  assign N412 = N411 & pe_o_1__3_;
  assign N413 = N412 & N417;
  assign N414 = N413 & N418;
  assign N7512 = N414 & pe_o_1__1_;
  assign N415 = ~pe_o_1__6_;
  assign N416 = ~pe_o_1__4_;
  assign N417 = ~pe_o_1__2_;
  assign N418 = ~pe_o_1__0_;
  assign N419 = N424 & pe_o_1__5_;
  assign N420 = N419 & N425;
  assign N421 = N420 & pe_o_1__3_;
  assign N422 = N421 & N426;
  assign N423 = N422 & pe_o_1__0_;
  assign N7514 = N423 & pe_o_1__1_;
  assign N424 = ~pe_o_1__6_;
  assign N425 = ~pe_o_1__4_;
  assign N426 = ~pe_o_1__2_;
  assign N427 = N432 & pe_o_1__5_;
  assign N428 = N427 & N433;
  assign N429 = N428 & pe_o_1__3_;
  assign N430 = N429 & pe_o_1__2_;
  assign N431 = N430 & N434;
  assign N7516 = N431 & N435;
  assign N432 = ~pe_o_1__6_;
  assign N433 = ~pe_o_1__4_;
  assign N434 = ~pe_o_1__0_;
  assign N435 = ~pe_o_1__1_;
  assign N436 = N441 & pe_o_1__5_;
  assign N437 = N436 & N442;
  assign N438 = N437 & pe_o_1__3_;
  assign N439 = N438 & pe_o_1__2_;
  assign N440 = N439 & pe_o_1__0_;
  assign N7518 = N440 & N443;
  assign N441 = ~pe_o_1__6_;
  assign N442 = ~pe_o_1__4_;
  assign N443 = ~pe_o_1__1_;
  assign N444 = N449 & pe_o_1__5_;
  assign N445 = N444 & N450;
  assign N446 = N445 & pe_o_1__3_;
  assign N447 = N446 & pe_o_1__2_;
  assign N448 = N447 & N451;
  assign N7520 = N448 & pe_o_1__1_;
  assign N449 = ~pe_o_1__6_;
  assign N450 = ~pe_o_1__4_;
  assign N451 = ~pe_o_1__0_;
  assign N452 = N457 & pe_o_1__5_;
  assign N453 = N452 & N458;
  assign N454 = N453 & pe_o_1__3_;
  assign N455 = N454 & pe_o_1__2_;
  assign N456 = N455 & pe_o_1__0_;
  assign N7522 = N456 & pe_o_1__1_;
  assign N457 = ~pe_o_1__6_;
  assign N458 = ~pe_o_1__4_;
  assign N459 = N464 & pe_o_1__5_;
  assign N460 = N459 & pe_o_1__4_;
  assign N461 = N460 & N465;
  assign N462 = N461 & N466;
  assign N463 = N462 & N467;
  assign N7524 = N463 & N468;
  assign N464 = ~pe_o_1__6_;
  assign N465 = ~pe_o_1__3_;
  assign N466 = ~pe_o_1__2_;
  assign N467 = ~pe_o_1__0_;
  assign N468 = ~pe_o_1__1_;
  assign N469 = N474 & pe_o_1__5_;
  assign N470 = N469 & pe_o_1__4_;
  assign N471 = N470 & N475;
  assign N472 = N471 & N476;
  assign N473 = N472 & pe_o_1__0_;
  assign N7526 = N473 & N477;
  assign N474 = ~pe_o_1__6_;
  assign N475 = ~pe_o_1__3_;
  assign N476 = ~pe_o_1__2_;
  assign N477 = ~pe_o_1__1_;
  assign N478 = N483 & pe_o_1__5_;
  assign N479 = N478 & pe_o_1__4_;
  assign N480 = N479 & N484;
  assign N481 = N480 & N485;
  assign N482 = N481 & N486;
  assign N7528 = N482 & pe_o_1__1_;
  assign N483 = ~pe_o_1__6_;
  assign N484 = ~pe_o_1__3_;
  assign N485 = ~pe_o_1__2_;
  assign N486 = ~pe_o_1__0_;
  assign N487 = N492 & pe_o_1__5_;
  assign N488 = N487 & pe_o_1__4_;
  assign N489 = N488 & N493;
  assign N490 = N489 & N494;
  assign N491 = N490 & pe_o_1__0_;
  assign N7530 = N491 & pe_o_1__1_;
  assign N492 = ~pe_o_1__6_;
  assign N493 = ~pe_o_1__3_;
  assign N494 = ~pe_o_1__2_;
  assign N495 = N500 & pe_o_1__5_;
  assign N496 = N495 & pe_o_1__4_;
  assign N497 = N496 & N501;
  assign N498 = N497 & pe_o_1__2_;
  assign N499 = N498 & N502;
  assign N7532 = N499 & N503;
  assign N500 = ~pe_o_1__6_;
  assign N501 = ~pe_o_1__3_;
  assign N502 = ~pe_o_1__0_;
  assign N503 = ~pe_o_1__1_;
  assign N504 = N509 & pe_o_1__5_;
  assign N505 = N504 & pe_o_1__4_;
  assign N506 = N505 & N510;
  assign N507 = N506 & pe_o_1__2_;
  assign N508 = N507 & pe_o_1__0_;
  assign N7534 = N508 & N511;
  assign N509 = ~pe_o_1__6_;
  assign N510 = ~pe_o_1__3_;
  assign N511 = ~pe_o_1__1_;
  assign N512 = N517 & pe_o_1__5_;
  assign N513 = N512 & pe_o_1__4_;
  assign N514 = N513 & N518;
  assign N515 = N514 & pe_o_1__2_;
  assign N516 = N515 & N519;
  assign N7536 = N516 & pe_o_1__1_;
  assign N517 = ~pe_o_1__6_;
  assign N518 = ~pe_o_1__3_;
  assign N519 = ~pe_o_1__0_;
  assign N520 = N525 & pe_o_1__5_;
  assign N521 = N520 & pe_o_1__4_;
  assign N522 = N521 & N526;
  assign N523 = N522 & pe_o_1__2_;
  assign N524 = N523 & pe_o_1__0_;
  assign N7538 = N524 & pe_o_1__1_;
  assign N525 = ~pe_o_1__6_;
  assign N526 = ~pe_o_1__3_;
  assign N527 = N532 & pe_o_1__5_;
  assign N528 = N527 & pe_o_1__4_;
  assign N529 = N528 & pe_o_1__3_;
  assign N530 = N529 & N533;
  assign N531 = N530 & N534;
  assign N7540 = N531 & N535;
  assign N532 = ~pe_o_1__6_;
  assign N533 = ~pe_o_1__2_;
  assign N534 = ~pe_o_1__0_;
  assign N535 = ~pe_o_1__1_;
  assign N536 = N541 & pe_o_1__5_;
  assign N537 = N536 & pe_o_1__4_;
  assign N538 = N537 & pe_o_1__3_;
  assign N539 = N538 & N542;
  assign N540 = N539 & pe_o_1__0_;
  assign N7542 = N540 & N543;
  assign N541 = ~pe_o_1__6_;
  assign N542 = ~pe_o_1__2_;
  assign N543 = ~pe_o_1__1_;
  assign N544 = N549 & pe_o_1__5_;
  assign N545 = N544 & pe_o_1__4_;
  assign N546 = N545 & pe_o_1__3_;
  assign N547 = N546 & N550;
  assign N548 = N547 & N551;
  assign N7544 = N548 & pe_o_1__1_;
  assign N549 = ~pe_o_1__6_;
  assign N550 = ~pe_o_1__2_;
  assign N551 = ~pe_o_1__0_;
  assign N552 = N557 & pe_o_1__5_;
  assign N553 = N552 & pe_o_1__4_;
  assign N554 = N553 & pe_o_1__3_;
  assign N555 = N554 & N558;
  assign N556 = N555 & pe_o_1__0_;
  assign N7546 = N556 & pe_o_1__1_;
  assign N557 = ~pe_o_1__6_;
  assign N558 = ~pe_o_1__2_;
  assign N559 = N564 & pe_o_1__5_;
  assign N560 = N559 & pe_o_1__4_;
  assign N561 = N560 & pe_o_1__3_;
  assign N562 = N561 & pe_o_1__2_;
  assign N563 = N562 & N565;
  assign N7548 = N563 & N566;
  assign N564 = ~pe_o_1__6_;
  assign N565 = ~pe_o_1__0_;
  assign N566 = ~pe_o_1__1_;
  assign N567 = N572 & pe_o_1__5_;
  assign N568 = N567 & pe_o_1__4_;
  assign N569 = N568 & pe_o_1__3_;
  assign N570 = N569 & pe_o_1__2_;
  assign N571 = N570 & pe_o_1__0_;
  assign N7550 = N571 & N573;
  assign N572 = ~pe_o_1__6_;
  assign N573 = ~pe_o_1__1_;
  assign N574 = N579 & pe_o_1__5_;
  assign N575 = N574 & pe_o_1__4_;
  assign N576 = N575 & pe_o_1__3_;
  assign N577 = N576 & pe_o_1__2_;
  assign N578 = N577 & N580;
  assign N7552 = N578 & pe_o_1__1_;
  assign N579 = ~pe_o_1__6_;
  assign N580 = ~pe_o_1__0_;
  assign N581 = pe_o_1__5_ & pe_o_1__4_;
  assign N582 = N581 & pe_o_1__3_;
  assign N583 = N582 & pe_o_1__2_;
  assign N584 = N583 & pe_o_1__0_;
  assign N7554 = N584 & pe_o_1__1_;
  assign N585 = pe_o_1__6_ & N590;
  assign N586 = N585 & N591;
  assign N587 = N586 & N592;
  assign N588 = N587 & N593;
  assign N589 = N588 & pe_o_1__0_;
  assign N7431 = N589 & N594;
  assign N590 = ~pe_o_1__5_;
  assign N591 = ~pe_o_1__4_;
  assign N592 = ~pe_o_1__3_;
  assign N593 = ~pe_o_1__2_;
  assign N594 = ~pe_o_1__1_;
  assign N595 = pe_o_1__6_ & N600;
  assign N596 = N595 & N601;
  assign N597 = N596 & N602;
  assign N598 = N597 & N603;
  assign N599 = N598 & N604;
  assign N7433 = N599 & pe_o_1__1_;
  assign N600 = ~pe_o_1__5_;
  assign N601 = ~pe_o_1__4_;
  assign N602 = ~pe_o_1__3_;
  assign N603 = ~pe_o_1__2_;
  assign N604 = ~pe_o_1__0_;
  assign N605 = pe_o_1__6_ & N610;
  assign N606 = N605 & N611;
  assign N607 = N606 & N612;
  assign N608 = N607 & N613;
  assign N609 = N608 & pe_o_1__0_;
  assign N7435 = N609 & pe_o_1__1_;
  assign N610 = ~pe_o_1__5_;
  assign N611 = ~pe_o_1__4_;
  assign N612 = ~pe_o_1__3_;
  assign N613 = ~pe_o_1__2_;
  assign N614 = pe_o_1__6_ & N619;
  assign N615 = N614 & N620;
  assign N616 = N615 & N621;
  assign N617 = N616 & pe_o_1__2_;
  assign N618 = N617 & N622;
  assign N7437 = N618 & N623;
  assign N619 = ~pe_o_1__5_;
  assign N620 = ~pe_o_1__4_;
  assign N621 = ~pe_o_1__3_;
  assign N622 = ~pe_o_1__0_;
  assign N623 = ~pe_o_1__1_;
  assign N624 = pe_o_1__6_ & N629;
  assign N625 = N624 & N630;
  assign N626 = N625 & N631;
  assign N627 = N626 & pe_o_1__2_;
  assign N628 = N627 & pe_o_1__0_;
  assign N7439 = N628 & N632;
  assign N629 = ~pe_o_1__5_;
  assign N630 = ~pe_o_1__4_;
  assign N631 = ~pe_o_1__3_;
  assign N632 = ~pe_o_1__1_;
  assign N633 = pe_o_1__6_ & N638;
  assign N634 = N633 & N639;
  assign N635 = N634 & N640;
  assign N636 = N635 & pe_o_1__2_;
  assign N637 = N636 & N641;
  assign N7441 = N637 & pe_o_1__1_;
  assign N638 = ~pe_o_1__5_;
  assign N639 = ~pe_o_1__4_;
  assign N640 = ~pe_o_1__3_;
  assign N641 = ~pe_o_1__0_;
  assign N642 = pe_o_1__6_ & N647;
  assign N643 = N642 & N648;
  assign N644 = N643 & N649;
  assign N645 = N644 & pe_o_1__2_;
  assign N646 = N645 & pe_o_1__0_;
  assign N7443 = N646 & pe_o_1__1_;
  assign N647 = ~pe_o_1__5_;
  assign N648 = ~pe_o_1__4_;
  assign N649 = ~pe_o_1__3_;
  assign N650 = pe_o_1__6_ & N655;
  assign N651 = N650 & N656;
  assign N652 = N651 & pe_o_1__3_;
  assign N653 = N652 & N657;
  assign N654 = N653 & N658;
  assign N7445 = N654 & N659;
  assign N655 = ~pe_o_1__5_;
  assign N656 = ~pe_o_1__4_;
  assign N657 = ~pe_o_1__2_;
  assign N658 = ~pe_o_1__0_;
  assign N659 = ~pe_o_1__1_;
  assign N660 = pe_o_1__6_ & N665;
  assign N661 = N660 & N666;
  assign N662 = N661 & pe_o_1__3_;
  assign N663 = N662 & N667;
  assign N664 = N663 & pe_o_1__0_;
  assign N7447 = N664 & N668;
  assign N665 = ~pe_o_1__5_;
  assign N666 = ~pe_o_1__4_;
  assign N667 = ~pe_o_1__2_;
  assign N668 = ~pe_o_1__1_;
  assign N669 = pe_o_1__6_ & N674;
  assign N670 = N669 & N675;
  assign N671 = N670 & pe_o_1__3_;
  assign N672 = N671 & N676;
  assign N673 = N672 & N677;
  assign N7449 = N673 & pe_o_1__1_;
  assign N674 = ~pe_o_1__5_;
  assign N675 = ~pe_o_1__4_;
  assign N676 = ~pe_o_1__2_;
  assign N677 = ~pe_o_1__0_;
  assign N678 = pe_o_1__6_ & N683;
  assign N679 = N678 & N684;
  assign N680 = N679 & pe_o_1__3_;
  assign N681 = N680 & N685;
  assign N682 = N681 & pe_o_1__0_;
  assign N7451 = N682 & pe_o_1__1_;
  assign N683 = ~pe_o_1__5_;
  assign N684 = ~pe_o_1__4_;
  assign N685 = ~pe_o_1__2_;
  assign N686 = pe_o_1__6_ & N691;
  assign N687 = N686 & N692;
  assign N688 = N687 & pe_o_1__3_;
  assign N689 = N688 & pe_o_1__2_;
  assign N690 = N689 & N693;
  assign N7453 = N690 & N694;
  assign N691 = ~pe_o_1__5_;
  assign N692 = ~pe_o_1__4_;
  assign N693 = ~pe_o_1__0_;
  assign N694 = ~pe_o_1__1_;
  assign N695 = pe_o_1__6_ & N700;
  assign N696 = N695 & N701;
  assign N697 = N696 & pe_o_1__3_;
  assign N698 = N697 & pe_o_1__2_;
  assign N699 = N698 & pe_o_1__0_;
  assign N7455 = N699 & N702;
  assign N700 = ~pe_o_1__5_;
  assign N701 = ~pe_o_1__4_;
  assign N702 = ~pe_o_1__1_;
  assign N703 = pe_o_1__6_ & N708;
  assign N704 = N703 & N709;
  assign N705 = N704 & pe_o_1__3_;
  assign N706 = N705 & pe_o_1__2_;
  assign N707 = N706 & N710;
  assign N7457 = N707 & pe_o_1__1_;
  assign N708 = ~pe_o_1__5_;
  assign N709 = ~pe_o_1__4_;
  assign N710 = ~pe_o_1__0_;
  assign N711 = pe_o_1__6_ & N716;
  assign N712 = N711 & N717;
  assign N713 = N712 & pe_o_1__3_;
  assign N714 = N713 & pe_o_1__2_;
  assign N715 = N714 & pe_o_1__0_;
  assign N7459 = N715 & pe_o_1__1_;
  assign N716 = ~pe_o_1__5_;
  assign N717 = ~pe_o_1__4_;
  assign N718 = pe_o_1__6_ & N723;
  assign N719 = N718 & pe_o_1__4_;
  assign N720 = N719 & N724;
  assign N721 = N720 & N725;
  assign N722 = N721 & N726;
  assign N7461 = N722 & N727;
  assign N723 = ~pe_o_1__5_;
  assign N724 = ~pe_o_1__3_;
  assign N725 = ~pe_o_1__2_;
  assign N726 = ~pe_o_1__0_;
  assign N727 = ~pe_o_1__1_;
  assign N728 = pe_o_1__6_ & N733;
  assign N729 = N728 & pe_o_1__4_;
  assign N730 = N729 & N734;
  assign N731 = N730 & N735;
  assign N732 = N731 & pe_o_1__0_;
  assign N7463 = N732 & N736;
  assign N733 = ~pe_o_1__5_;
  assign N734 = ~pe_o_1__3_;
  assign N735 = ~pe_o_1__2_;
  assign N736 = ~pe_o_1__1_;
  assign N737 = pe_o_1__6_ & N742;
  assign N738 = N737 & pe_o_1__4_;
  assign N739 = N738 & N743;
  assign N740 = N739 & N744;
  assign N741 = N740 & N745;
  assign N7465 = N741 & pe_o_1__1_;
  assign N742 = ~pe_o_1__5_;
  assign N743 = ~pe_o_1__3_;
  assign N744 = ~pe_o_1__2_;
  assign N745 = ~pe_o_1__0_;
  assign N746 = pe_o_1__6_ & N751;
  assign N747 = N746 & pe_o_1__4_;
  assign N748 = N747 & N752;
  assign N749 = N748 & N753;
  assign N750 = N749 & pe_o_1__0_;
  assign N7467 = N750 & pe_o_1__1_;
  assign N751 = ~pe_o_1__5_;
  assign N752 = ~pe_o_1__3_;
  assign N753 = ~pe_o_1__2_;
  assign N754 = pe_o_1__6_ & N759;
  assign N755 = N754 & pe_o_1__4_;
  assign N756 = N755 & N760;
  assign N757 = N756 & pe_o_1__2_;
  assign N758 = N757 & N761;
  assign N7469 = N758 & N762;
  assign N759 = ~pe_o_1__5_;
  assign N760 = ~pe_o_1__3_;
  assign N761 = ~pe_o_1__0_;
  assign N762 = ~pe_o_1__1_;
  assign N763 = pe_o_1__6_ & N768;
  assign N764 = N763 & pe_o_1__4_;
  assign N765 = N764 & N769;
  assign N766 = N765 & pe_o_1__2_;
  assign N767 = N766 & pe_o_1__0_;
  assign N7471 = N767 & N770;
  assign N768 = ~pe_o_1__5_;
  assign N769 = ~pe_o_1__3_;
  assign N770 = ~pe_o_1__1_;
  assign N771 = pe_o_1__6_ & N776;
  assign N772 = N771 & pe_o_1__4_;
  assign N773 = N772 & N777;
  assign N774 = N773 & pe_o_1__2_;
  assign N775 = N774 & N778;
  assign N7473 = N775 & pe_o_1__1_;
  assign N776 = ~pe_o_1__5_;
  assign N777 = ~pe_o_1__3_;
  assign N778 = ~pe_o_1__0_;
  assign N779 = pe_o_1__6_ & N784;
  assign N780 = N779 & pe_o_1__4_;
  assign N781 = N780 & N785;
  assign N782 = N781 & pe_o_1__2_;
  assign N783 = N782 & pe_o_1__0_;
  assign N7475 = N783 & pe_o_1__1_;
  assign N784 = ~pe_o_1__5_;
  assign N785 = ~pe_o_1__3_;
  assign N786 = pe_o_1__6_ & N791;
  assign N787 = N786 & pe_o_1__4_;
  assign N788 = N787 & pe_o_1__3_;
  assign N789 = N788 & N792;
  assign N790 = N789 & N793;
  assign N7477 = N790 & N794;
  assign N791 = ~pe_o_1__5_;
  assign N792 = ~pe_o_1__2_;
  assign N793 = ~pe_o_1__0_;
  assign N794 = ~pe_o_1__1_;
  assign N795 = pe_o_1__6_ & N800;
  assign N796 = N795 & pe_o_1__4_;
  assign N797 = N796 & pe_o_1__3_;
  assign N798 = N797 & N801;
  assign N799 = N798 & pe_o_1__0_;
  assign N7479 = N799 & N802;
  assign N800 = ~pe_o_1__5_;
  assign N801 = ~pe_o_1__2_;
  assign N802 = ~pe_o_1__1_;
  assign N803 = pe_o_1__6_ & N808;
  assign N804 = N803 & pe_o_1__4_;
  assign N805 = N804 & pe_o_1__3_;
  assign N806 = N805 & N809;
  assign N807 = N806 & N810;
  assign N7481 = N807 & pe_o_1__1_;
  assign N808 = ~pe_o_1__5_;
  assign N809 = ~pe_o_1__2_;
  assign N810 = ~pe_o_1__0_;
  assign N811 = pe_o_1__6_ & N816;
  assign N812 = N811 & pe_o_1__4_;
  assign N813 = N812 & pe_o_1__3_;
  assign N814 = N813 & N817;
  assign N815 = N814 & pe_o_1__0_;
  assign N7483 = N815 & pe_o_1__1_;
  assign N816 = ~pe_o_1__5_;
  assign N817 = ~pe_o_1__2_;
  assign N818 = pe_o_1__6_ & N823;
  assign N819 = N818 & pe_o_1__4_;
  assign N820 = N819 & pe_o_1__3_;
  assign N821 = N820 & pe_o_1__2_;
  assign N822 = N821 & N824;
  assign N7485 = N822 & N825;
  assign N823 = ~pe_o_1__5_;
  assign N824 = ~pe_o_1__0_;
  assign N825 = ~pe_o_1__1_;
  assign N826 = pe_o_1__6_ & N831;
  assign N827 = N826 & pe_o_1__4_;
  assign N828 = N827 & pe_o_1__3_;
  assign N829 = N828 & pe_o_1__2_;
  assign N830 = N829 & pe_o_1__0_;
  assign N7487 = N830 & N832;
  assign N831 = ~pe_o_1__5_;
  assign N832 = ~pe_o_1__1_;
  assign N833 = pe_o_1__6_ & N838;
  assign N834 = N833 & pe_o_1__4_;
  assign N835 = N834 & pe_o_1__3_;
  assign N836 = N835 & pe_o_1__2_;
  assign N837 = N836 & N839;
  assign N7489 = N837 & pe_o_1__1_;
  assign N838 = ~pe_o_1__5_;
  assign N839 = ~pe_o_1__0_;
  assign N840 = pe_o_1__6_ & pe_o_1__4_;
  assign N841 = N840 & pe_o_1__3_;
  assign N842 = N841 & pe_o_1__2_;
  assign N843 = N842 & pe_o_1__0_;
  assign N7491 = N843 & pe_o_1__1_;
  assign N844 = pe_o_1__6_ & pe_o_1__5_;
  assign N845 = N844 & N849;
  assign N846 = N845 & N850;
  assign N847 = N846 & N851;
  assign N848 = N847 & N852;
  assign N7493 = N848 & N853;
  assign N849 = ~pe_o_1__4_;
  assign N850 = ~pe_o_1__3_;
  assign N851 = ~pe_o_1__2_;
  assign N852 = ~pe_o_1__0_;
  assign N853 = ~pe_o_1__1_;
  assign N854 = pe_o_1__6_ & pe_o_1__5_;
  assign N855 = N854 & N859;
  assign N856 = N855 & N860;
  assign N857 = N856 & N861;
  assign N858 = N857 & pe_o_1__0_;
  assign N7495 = N858 & N862;
  assign N859 = ~pe_o_1__4_;
  assign N860 = ~pe_o_1__3_;
  assign N861 = ~pe_o_1__2_;
  assign N862 = ~pe_o_1__1_;
  assign N863 = pe_o_1__6_ & pe_o_1__5_;
  assign N864 = N863 & N868;
  assign N865 = N864 & N869;
  assign N866 = N865 & N870;
  assign N867 = N866 & N871;
  assign N7497 = N867 & pe_o_1__1_;
  assign N868 = ~pe_o_1__4_;
  assign N869 = ~pe_o_1__3_;
  assign N870 = ~pe_o_1__2_;
  assign N871 = ~pe_o_1__0_;
  assign N872 = pe_o_1__6_ & pe_o_1__5_;
  assign N873 = N872 & N877;
  assign N874 = N873 & N878;
  assign N875 = N874 & N879;
  assign N876 = N875 & pe_o_1__0_;
  assign N7499 = N876 & pe_o_1__1_;
  assign N877 = ~pe_o_1__4_;
  assign N878 = ~pe_o_1__3_;
  assign N879 = ~pe_o_1__2_;
  assign N880 = pe_o_1__6_ & pe_o_1__5_;
  assign N881 = N880 & N885;
  assign N882 = N881 & N886;
  assign N883 = N882 & pe_o_1__2_;
  assign N884 = N883 & N887;
  assign N7501 = N884 & N888;
  assign N885 = ~pe_o_1__4_;
  assign N886 = ~pe_o_1__3_;
  assign N887 = ~pe_o_1__0_;
  assign N888 = ~pe_o_1__1_;
  assign N889 = pe_o_1__6_ & pe_o_1__5_;
  assign N890 = N889 & N894;
  assign N891 = N890 & N895;
  assign N892 = N891 & pe_o_1__2_;
  assign N893 = N892 & pe_o_1__0_;
  assign N7503 = N893 & N896;
  assign N894 = ~pe_o_1__4_;
  assign N895 = ~pe_o_1__3_;
  assign N896 = ~pe_o_1__1_;
  assign N897 = pe_o_1__6_ & pe_o_1__5_;
  assign N898 = N897 & N902;
  assign N899 = N898 & N903;
  assign N900 = N899 & pe_o_1__2_;
  assign N901 = N900 & N904;
  assign N7505 = N901 & pe_o_1__1_;
  assign N902 = ~pe_o_1__4_;
  assign N903 = ~pe_o_1__3_;
  assign N904 = ~pe_o_1__0_;
  assign N905 = pe_o_1__6_ & pe_o_1__5_;
  assign N906 = N905 & N910;
  assign N907 = N906 & N911;
  assign N908 = N907 & pe_o_1__2_;
  assign N909 = N908 & pe_o_1__0_;
  assign N7507 = N909 & pe_o_1__1_;
  assign N910 = ~pe_o_1__4_;
  assign N911 = ~pe_o_1__3_;
  assign N912 = pe_o_1__6_ & pe_o_1__5_;
  assign N913 = N912 & N917;
  assign N914 = N913 & pe_o_1__3_;
  assign N915 = N914 & N918;
  assign N916 = N915 & N919;
  assign N7509 = N916 & N920;
  assign N917 = ~pe_o_1__4_;
  assign N918 = ~pe_o_1__2_;
  assign N919 = ~pe_o_1__0_;
  assign N920 = ~pe_o_1__1_;
  assign N921 = pe_o_1__6_ & pe_o_1__5_;
  assign N922 = N921 & N926;
  assign N923 = N922 & pe_o_1__3_;
  assign N924 = N923 & N927;
  assign N925 = N924 & pe_o_1__0_;
  assign N7511 = N925 & N928;
  assign N926 = ~pe_o_1__4_;
  assign N927 = ~pe_o_1__2_;
  assign N928 = ~pe_o_1__1_;
  assign N929 = pe_o_1__6_ & pe_o_1__5_;
  assign N930 = N929 & N934;
  assign N931 = N930 & pe_o_1__3_;
  assign N932 = N931 & N935;
  assign N933 = N932 & N936;
  assign N7513 = N933 & pe_o_1__1_;
  assign N934 = ~pe_o_1__4_;
  assign N935 = ~pe_o_1__2_;
  assign N936 = ~pe_o_1__0_;
  assign N937 = pe_o_1__6_ & pe_o_1__5_;
  assign N938 = N937 & N942;
  assign N939 = N938 & pe_o_1__3_;
  assign N940 = N939 & N943;
  assign N941 = N940 & pe_o_1__0_;
  assign N7515 = N941 & pe_o_1__1_;
  assign N942 = ~pe_o_1__4_;
  assign N943 = ~pe_o_1__2_;
  assign N944 = pe_o_1__6_ & pe_o_1__5_;
  assign N945 = N944 & N949;
  assign N946 = N945 & pe_o_1__3_;
  assign N947 = N946 & pe_o_1__2_;
  assign N948 = N947 & N950;
  assign N7517 = N948 & N951;
  assign N949 = ~pe_o_1__4_;
  assign N950 = ~pe_o_1__0_;
  assign N951 = ~pe_o_1__1_;
  assign N952 = pe_o_1__6_ & pe_o_1__5_;
  assign N953 = N952 & N957;
  assign N954 = N953 & pe_o_1__3_;
  assign N955 = N954 & pe_o_1__2_;
  assign N956 = N955 & pe_o_1__0_;
  assign N7519 = N956 & N958;
  assign N957 = ~pe_o_1__4_;
  assign N958 = ~pe_o_1__1_;
  assign N959 = pe_o_1__6_ & pe_o_1__5_;
  assign N960 = N959 & N964;
  assign N961 = N960 & pe_o_1__3_;
  assign N962 = N961 & pe_o_1__2_;
  assign N963 = N962 & N965;
  assign N7521 = N963 & pe_o_1__1_;
  assign N964 = ~pe_o_1__4_;
  assign N965 = ~pe_o_1__0_;
  assign N966 = pe_o_1__6_ & pe_o_1__5_;
  assign N967 = N966 & pe_o_1__3_;
  assign N968 = N967 & pe_o_1__2_;
  assign N969 = N968 & pe_o_1__0_;
  assign N7523 = N969 & pe_o_1__1_;
  assign N970 = pe_o_1__6_ & pe_o_1__5_;
  assign N971 = N970 & pe_o_1__4_;
  assign N972 = N971 & N975;
  assign N973 = N972 & N976;
  assign N974 = N973 & N977;
  assign N7525 = N974 & N978;
  assign N975 = ~pe_o_1__3_;
  assign N976 = ~pe_o_1__2_;
  assign N977 = ~pe_o_1__0_;
  assign N978 = ~pe_o_1__1_;
  assign N979 = pe_o_1__6_ & pe_o_1__5_;
  assign N980 = N979 & pe_o_1__4_;
  assign N981 = N980 & N984;
  assign N982 = N981 & N985;
  assign N983 = N982 & pe_o_1__0_;
  assign N7527 = N983 & N986;
  assign N984 = ~pe_o_1__3_;
  assign N985 = ~pe_o_1__2_;
  assign N986 = ~pe_o_1__1_;
  assign N987 = pe_o_1__6_ & pe_o_1__5_;
  assign N988 = N987 & pe_o_1__4_;
  assign N989 = N988 & N992;
  assign N990 = N989 & N993;
  assign N991 = N990 & N994;
  assign N7529 = N991 & pe_o_1__1_;
  assign N992 = ~pe_o_1__3_;
  assign N993 = ~pe_o_1__2_;
  assign N994 = ~pe_o_1__0_;
  assign N995 = pe_o_1__6_ & pe_o_1__5_;
  assign N996 = N995 & pe_o_1__4_;
  assign N997 = N996 & N1000;
  assign N998 = N997 & N1001;
  assign N999 = N998 & pe_o_1__0_;
  assign N7531 = N999 & pe_o_1__1_;
  assign N1000 = ~pe_o_1__3_;
  assign N1001 = ~pe_o_1__2_;
  assign N1002 = pe_o_1__6_ & pe_o_1__5_;
  assign N1003 = N1002 & pe_o_1__4_;
  assign N1004 = N1003 & N1007;
  assign N1005 = N1004 & pe_o_1__2_;
  assign N1006 = N1005 & N1008;
  assign N7533 = N1006 & N1009;
  assign N1007 = ~pe_o_1__3_;
  assign N1008 = ~pe_o_1__0_;
  assign N1009 = ~pe_o_1__1_;
  assign N1010 = pe_o_1__6_ & pe_o_1__5_;
  assign N1011 = N1010 & pe_o_1__4_;
  assign N1012 = N1011 & N1015;
  assign N1013 = N1012 & pe_o_1__2_;
  assign N1014 = N1013 & pe_o_1__0_;
  assign N7535 = N1014 & N1016;
  assign N1015 = ~pe_o_1__3_;
  assign N1016 = ~pe_o_1__1_;
  assign N1017 = pe_o_1__6_ & pe_o_1__5_;
  assign N1018 = N1017 & pe_o_1__4_;
  assign N1019 = N1018 & N1022;
  assign N1020 = N1019 & pe_o_1__2_;
  assign N1021 = N1020 & N1023;
  assign N7537 = N1021 & pe_o_1__1_;
  assign N1022 = ~pe_o_1__3_;
  assign N1023 = ~pe_o_1__0_;
  assign N1024 = pe_o_1__6_ & pe_o_1__5_;
  assign N1025 = N1024 & pe_o_1__4_;
  assign N1026 = N1025 & pe_o_1__2_;
  assign N1027 = N1026 & pe_o_1__0_;
  assign N7539 = N1027 & pe_o_1__1_;
  assign N1028 = pe_o_1__6_ & pe_o_1__5_;
  assign N1029 = N1028 & pe_o_1__4_;
  assign N1030 = N1029 & pe_o_1__3_;
  assign N1031 = N1030 & N1033;
  assign N1032 = N1031 & N1034;
  assign N7541 = N1032 & N1035;
  assign N1033 = ~pe_o_1__2_;
  assign N1034 = ~pe_o_1__0_;
  assign N1035 = ~pe_o_1__1_;
  assign N1036 = pe_o_1__6_ & pe_o_1__5_;
  assign N1037 = N1036 & pe_o_1__4_;
  assign N1038 = N1037 & pe_o_1__3_;
  assign N1039 = N1038 & N1041;
  assign N1040 = N1039 & pe_o_1__0_;
  assign N7543 = N1040 & N1042;
  assign N1041 = ~pe_o_1__2_;
  assign N1042 = ~pe_o_1__1_;
  assign N1043 = pe_o_1__6_ & pe_o_1__5_;
  assign N1044 = N1043 & pe_o_1__4_;
  assign N1045 = N1044 & pe_o_1__3_;
  assign N1046 = N1045 & N1048;
  assign N1047 = N1046 & N1049;
  assign N7545 = N1047 & pe_o_1__1_;
  assign N1048 = ~pe_o_1__2_;
  assign N1049 = ~pe_o_1__0_;
  assign N1050 = pe_o_1__6_ & pe_o_1__5_;
  assign N1051 = N1050 & pe_o_1__4_;
  assign N1052 = N1051 & pe_o_1__3_;
  assign N1053 = N1052 & pe_o_1__0_;
  assign N7547 = N1053 & pe_o_1__1_;
  assign N1054 = pe_o_1__6_ & pe_o_1__5_;
  assign N1055 = N1054 & pe_o_1__4_;
  assign N1056 = N1055 & pe_o_1__3_;
  assign N1057 = N1056 & pe_o_1__2_;
  assign N1058 = N1057 & N1059;
  assign N7549 = N1058 & N1060;
  assign N1059 = ~pe_o_1__0_;
  assign N1060 = ~pe_o_1__1_;
  assign N1061 = pe_o_1__6_ & pe_o_1__5_;
  assign N1062 = N1061 & pe_o_1__4_;
  assign N1063 = N1062 & pe_o_1__3_;
  assign N1064 = N1063 & pe_o_1__2_;
  assign N7551 = N1064 & pe_o_1__0_;
  assign N1065 = pe_o_1__6_ & pe_o_1__5_;
  assign N1066 = N1065 & pe_o_1__4_;
  assign N1067 = N1066 & pe_o_1__3_;
  assign N1068 = N1067 & pe_o_1__2_;
  assign N7553 = N1068 & pe_o_1__1_;
  assign N1069 = N1074 & N1075;
  assign N1070 = N1069 & N1076;
  assign N1071 = N1070 & N1077;
  assign N1072 = N1071 & N1078;
  assign N1073 = N1072 & N1079;
  assign N7555 = N1073 & N1080;
  assign N1074 = ~pe_o_2__6_;
  assign N1075 = ~pe_o_2__5_;
  assign N1076 = ~pe_o_2__4_;
  assign N1077 = ~pe_o_2__3_;
  assign N1078 = ~pe_o_2__2_;
  assign N1079 = ~pe_o_2__0_;
  assign N1080 = ~pe_o_2__1_;
  assign N1081 = pe_o_2__6_ & N1086;
  assign N1082 = N1081 & N1087;
  assign N1083 = N1082 & N1088;
  assign N1084 = N1083 & N1089;
  assign N1085 = N1084 & N1090;
  assign N7556 = N1085 & N1091;
  assign N1086 = ~pe_o_2__5_;
  assign N1087 = ~pe_o_2__4_;
  assign N1088 = ~pe_o_2__3_;
  assign N1089 = ~pe_o_2__2_;
  assign N1090 = ~pe_o_2__0_;
  assign N1091 = ~pe_o_2__1_;
  assign N1092 = N1097 & N1098;
  assign N1093 = N1092 & N1099;
  assign N1094 = N1093 & N1100;
  assign N1095 = N1094 & N1101;
  assign N1096 = N1095 & pe_o_2__0_;
  assign N7557 = N1096 & N1102;
  assign N1097 = ~pe_o_2__6_;
  assign N1098 = ~pe_o_2__5_;
  assign N1099 = ~pe_o_2__4_;
  assign N1100 = ~pe_o_2__3_;
  assign N1101 = ~pe_o_2__2_;
  assign N1102 = ~pe_o_2__1_;
  assign N1103 = N1108 & N1109;
  assign N1104 = N1103 & N1110;
  assign N1105 = N1104 & N1111;
  assign N1106 = N1105 & N1112;
  assign N1107 = N1106 & N1113;
  assign N7559 = N1107 & pe_o_2__1_;
  assign N1108 = ~pe_o_2__6_;
  assign N1109 = ~pe_o_2__5_;
  assign N1110 = ~pe_o_2__4_;
  assign N1111 = ~pe_o_2__3_;
  assign N1112 = ~pe_o_2__2_;
  assign N1113 = ~pe_o_2__0_;
  assign N1114 = N1119 & N1120;
  assign N1115 = N1114 & N1121;
  assign N1116 = N1115 & N1122;
  assign N1117 = N1116 & N1123;
  assign N1118 = N1117 & pe_o_2__0_;
  assign N7561 = N1118 & pe_o_2__1_;
  assign N1119 = ~pe_o_2__6_;
  assign N1120 = ~pe_o_2__5_;
  assign N1121 = ~pe_o_2__4_;
  assign N1122 = ~pe_o_2__3_;
  assign N1123 = ~pe_o_2__2_;
  assign N1124 = N1129 & N1130;
  assign N1125 = N1124 & N1131;
  assign N1126 = N1125 & N1132;
  assign N1127 = N1126 & pe_o_2__2_;
  assign N1128 = N1127 & N1133;
  assign N7563 = N1128 & N1134;
  assign N1129 = ~pe_o_2__6_;
  assign N1130 = ~pe_o_2__5_;
  assign N1131 = ~pe_o_2__4_;
  assign N1132 = ~pe_o_2__3_;
  assign N1133 = ~pe_o_2__0_;
  assign N1134 = ~pe_o_2__1_;
  assign N1135 = N1140 & N1141;
  assign N1136 = N1135 & N1142;
  assign N1137 = N1136 & N1143;
  assign N1138 = N1137 & pe_o_2__2_;
  assign N1139 = N1138 & pe_o_2__0_;
  assign N7565 = N1139 & N1144;
  assign N1140 = ~pe_o_2__6_;
  assign N1141 = ~pe_o_2__5_;
  assign N1142 = ~pe_o_2__4_;
  assign N1143 = ~pe_o_2__3_;
  assign N1144 = ~pe_o_2__1_;
  assign N1145 = N1150 & N1151;
  assign N1146 = N1145 & N1152;
  assign N1147 = N1146 & N1153;
  assign N1148 = N1147 & pe_o_2__2_;
  assign N1149 = N1148 & N1154;
  assign N7567 = N1149 & pe_o_2__1_;
  assign N1150 = ~pe_o_2__6_;
  assign N1151 = ~pe_o_2__5_;
  assign N1152 = ~pe_o_2__4_;
  assign N1153 = ~pe_o_2__3_;
  assign N1154 = ~pe_o_2__0_;
  assign N1155 = N1160 & N1161;
  assign N1156 = N1155 & N1162;
  assign N1157 = N1156 & N1163;
  assign N1158 = N1157 & pe_o_2__2_;
  assign N1159 = N1158 & pe_o_2__0_;
  assign N7569 = N1159 & pe_o_2__1_;
  assign N1160 = ~pe_o_2__6_;
  assign N1161 = ~pe_o_2__5_;
  assign N1162 = ~pe_o_2__4_;
  assign N1163 = ~pe_o_2__3_;
  assign N1164 = N1169 & N1170;
  assign N1165 = N1164 & N1171;
  assign N1166 = N1165 & pe_o_2__3_;
  assign N1167 = N1166 & N1172;
  assign N1168 = N1167 & N1173;
  assign N7571 = N1168 & N1174;
  assign N1169 = ~pe_o_2__6_;
  assign N1170 = ~pe_o_2__5_;
  assign N1171 = ~pe_o_2__4_;
  assign N1172 = ~pe_o_2__2_;
  assign N1173 = ~pe_o_2__0_;
  assign N1174 = ~pe_o_2__1_;
  assign N1175 = N1180 & N1181;
  assign N1176 = N1175 & N1182;
  assign N1177 = N1176 & pe_o_2__3_;
  assign N1178 = N1177 & N1183;
  assign N1179 = N1178 & pe_o_2__0_;
  assign N7573 = N1179 & N1184;
  assign N1180 = ~pe_o_2__6_;
  assign N1181 = ~pe_o_2__5_;
  assign N1182 = ~pe_o_2__4_;
  assign N1183 = ~pe_o_2__2_;
  assign N1184 = ~pe_o_2__1_;
  assign N1185 = N1190 & N1191;
  assign N1186 = N1185 & N1192;
  assign N1187 = N1186 & pe_o_2__3_;
  assign N1188 = N1187 & N1193;
  assign N1189 = N1188 & N1194;
  assign N7575 = N1189 & pe_o_2__1_;
  assign N1190 = ~pe_o_2__6_;
  assign N1191 = ~pe_o_2__5_;
  assign N1192 = ~pe_o_2__4_;
  assign N1193 = ~pe_o_2__2_;
  assign N1194 = ~pe_o_2__0_;
  assign N1195 = N1200 & N1201;
  assign N1196 = N1195 & N1202;
  assign N1197 = N1196 & pe_o_2__3_;
  assign N1198 = N1197 & N1203;
  assign N1199 = N1198 & pe_o_2__0_;
  assign N7577 = N1199 & pe_o_2__1_;
  assign N1200 = ~pe_o_2__6_;
  assign N1201 = ~pe_o_2__5_;
  assign N1202 = ~pe_o_2__4_;
  assign N1203 = ~pe_o_2__2_;
  assign N1204 = N1209 & N1210;
  assign N1205 = N1204 & N1211;
  assign N1206 = N1205 & pe_o_2__3_;
  assign N1207 = N1206 & pe_o_2__2_;
  assign N1208 = N1207 & N1212;
  assign N7579 = N1208 & N1213;
  assign N1209 = ~pe_o_2__6_;
  assign N1210 = ~pe_o_2__5_;
  assign N1211 = ~pe_o_2__4_;
  assign N1212 = ~pe_o_2__0_;
  assign N1213 = ~pe_o_2__1_;
  assign N1214 = N1219 & N1220;
  assign N1215 = N1214 & N1221;
  assign N1216 = N1215 & pe_o_2__3_;
  assign N1217 = N1216 & pe_o_2__2_;
  assign N1218 = N1217 & pe_o_2__0_;
  assign N7581 = N1218 & N1222;
  assign N1219 = ~pe_o_2__6_;
  assign N1220 = ~pe_o_2__5_;
  assign N1221 = ~pe_o_2__4_;
  assign N1222 = ~pe_o_2__1_;
  assign N1223 = N1228 & N1229;
  assign N1224 = N1223 & N1230;
  assign N1225 = N1224 & pe_o_2__3_;
  assign N1226 = N1225 & pe_o_2__2_;
  assign N1227 = N1226 & N1231;
  assign N7583 = N1227 & pe_o_2__1_;
  assign N1228 = ~pe_o_2__6_;
  assign N1229 = ~pe_o_2__5_;
  assign N1230 = ~pe_o_2__4_;
  assign N1231 = ~pe_o_2__0_;
  assign N1232 = N1237 & N1238;
  assign N1233 = N1232 & N1239;
  assign N1234 = N1233 & pe_o_2__3_;
  assign N1235 = N1234 & pe_o_2__2_;
  assign N1236 = N1235 & pe_o_2__0_;
  assign N7585 = N1236 & pe_o_2__1_;
  assign N1237 = ~pe_o_2__6_;
  assign N1238 = ~pe_o_2__5_;
  assign N1239 = ~pe_o_2__4_;
  assign N1240 = N1245 & N1246;
  assign N1241 = N1240 & pe_o_2__4_;
  assign N1242 = N1241 & N1247;
  assign N1243 = N1242 & N1248;
  assign N1244 = N1243 & N1249;
  assign N7587 = N1244 & N1250;
  assign N1245 = ~pe_o_2__6_;
  assign N1246 = ~pe_o_2__5_;
  assign N1247 = ~pe_o_2__3_;
  assign N1248 = ~pe_o_2__2_;
  assign N1249 = ~pe_o_2__0_;
  assign N1250 = ~pe_o_2__1_;
  assign N1251 = N1256 & N1257;
  assign N1252 = N1251 & pe_o_2__4_;
  assign N1253 = N1252 & N1258;
  assign N1254 = N1253 & N1259;
  assign N1255 = N1254 & pe_o_2__0_;
  assign N7589 = N1255 & N1260;
  assign N1256 = ~pe_o_2__6_;
  assign N1257 = ~pe_o_2__5_;
  assign N1258 = ~pe_o_2__3_;
  assign N1259 = ~pe_o_2__2_;
  assign N1260 = ~pe_o_2__1_;
  assign N1261 = N1266 & N1267;
  assign N1262 = N1261 & pe_o_2__4_;
  assign N1263 = N1262 & N1268;
  assign N1264 = N1263 & N1269;
  assign N1265 = N1264 & N1270;
  assign N7591 = N1265 & pe_o_2__1_;
  assign N1266 = ~pe_o_2__6_;
  assign N1267 = ~pe_o_2__5_;
  assign N1268 = ~pe_o_2__3_;
  assign N1269 = ~pe_o_2__2_;
  assign N1270 = ~pe_o_2__0_;
  assign N1271 = N1276 & N1277;
  assign N1272 = N1271 & pe_o_2__4_;
  assign N1273 = N1272 & N1278;
  assign N1274 = N1273 & N1279;
  assign N1275 = N1274 & pe_o_2__0_;
  assign N7593 = N1275 & pe_o_2__1_;
  assign N1276 = ~pe_o_2__6_;
  assign N1277 = ~pe_o_2__5_;
  assign N1278 = ~pe_o_2__3_;
  assign N1279 = ~pe_o_2__2_;
  assign N1280 = N1285 & N1286;
  assign N1281 = N1280 & pe_o_2__4_;
  assign N1282 = N1281 & N1287;
  assign N1283 = N1282 & pe_o_2__2_;
  assign N1284 = N1283 & N1288;
  assign N7595 = N1284 & N1289;
  assign N1285 = ~pe_o_2__6_;
  assign N1286 = ~pe_o_2__5_;
  assign N1287 = ~pe_o_2__3_;
  assign N1288 = ~pe_o_2__0_;
  assign N1289 = ~pe_o_2__1_;
  assign N1290 = N1295 & N1296;
  assign N1291 = N1290 & pe_o_2__4_;
  assign N1292 = N1291 & N1297;
  assign N1293 = N1292 & pe_o_2__2_;
  assign N1294 = N1293 & pe_o_2__0_;
  assign N7597 = N1294 & N1298;
  assign N1295 = ~pe_o_2__6_;
  assign N1296 = ~pe_o_2__5_;
  assign N1297 = ~pe_o_2__3_;
  assign N1298 = ~pe_o_2__1_;
  assign N1299 = N1304 & N1305;
  assign N1300 = N1299 & pe_o_2__4_;
  assign N1301 = N1300 & N1306;
  assign N1302 = N1301 & pe_o_2__2_;
  assign N1303 = N1302 & N1307;
  assign N7599 = N1303 & pe_o_2__1_;
  assign N1304 = ~pe_o_2__6_;
  assign N1305 = ~pe_o_2__5_;
  assign N1306 = ~pe_o_2__3_;
  assign N1307 = ~pe_o_2__0_;
  assign N1308 = N1313 & N1314;
  assign N1309 = N1308 & pe_o_2__4_;
  assign N1310 = N1309 & N1315;
  assign N1311 = N1310 & pe_o_2__2_;
  assign N1312 = N1311 & pe_o_2__0_;
  assign N7601 = N1312 & pe_o_2__1_;
  assign N1313 = ~pe_o_2__6_;
  assign N1314 = ~pe_o_2__5_;
  assign N1315 = ~pe_o_2__3_;
  assign N1316 = N1321 & N1322;
  assign N1317 = N1316 & pe_o_2__4_;
  assign N1318 = N1317 & pe_o_2__3_;
  assign N1319 = N1318 & N1323;
  assign N1320 = N1319 & N1324;
  assign N7603 = N1320 & N1325;
  assign N1321 = ~pe_o_2__6_;
  assign N1322 = ~pe_o_2__5_;
  assign N1323 = ~pe_o_2__2_;
  assign N1324 = ~pe_o_2__0_;
  assign N1325 = ~pe_o_2__1_;
  assign N1326 = N1331 & N1332;
  assign N1327 = N1326 & pe_o_2__4_;
  assign N1328 = N1327 & pe_o_2__3_;
  assign N1329 = N1328 & N1333;
  assign N1330 = N1329 & pe_o_2__0_;
  assign N7605 = N1330 & N1334;
  assign N1331 = ~pe_o_2__6_;
  assign N1332 = ~pe_o_2__5_;
  assign N1333 = ~pe_o_2__2_;
  assign N1334 = ~pe_o_2__1_;
  assign N1335 = N1340 & N1341;
  assign N1336 = N1335 & pe_o_2__4_;
  assign N1337 = N1336 & pe_o_2__3_;
  assign N1338 = N1337 & N1342;
  assign N1339 = N1338 & N1343;
  assign N7607 = N1339 & pe_o_2__1_;
  assign N1340 = ~pe_o_2__6_;
  assign N1341 = ~pe_o_2__5_;
  assign N1342 = ~pe_o_2__2_;
  assign N1343 = ~pe_o_2__0_;
  assign N1344 = N1349 & N1350;
  assign N1345 = N1344 & pe_o_2__4_;
  assign N1346 = N1345 & pe_o_2__3_;
  assign N1347 = N1346 & N1351;
  assign N1348 = N1347 & pe_o_2__0_;
  assign N7609 = N1348 & pe_o_2__1_;
  assign N1349 = ~pe_o_2__6_;
  assign N1350 = ~pe_o_2__5_;
  assign N1351 = ~pe_o_2__2_;
  assign N1352 = N1357 & N1358;
  assign N1353 = N1352 & pe_o_2__4_;
  assign N1354 = N1353 & pe_o_2__3_;
  assign N1355 = N1354 & pe_o_2__2_;
  assign N1356 = N1355 & N1359;
  assign N7611 = N1356 & N1360;
  assign N1357 = ~pe_o_2__6_;
  assign N1358 = ~pe_o_2__5_;
  assign N1359 = ~pe_o_2__0_;
  assign N1360 = ~pe_o_2__1_;
  assign N1361 = N1366 & N1367;
  assign N1362 = N1361 & pe_o_2__4_;
  assign N1363 = N1362 & pe_o_2__3_;
  assign N1364 = N1363 & pe_o_2__2_;
  assign N1365 = N1364 & pe_o_2__0_;
  assign N7613 = N1365 & N1368;
  assign N1366 = ~pe_o_2__6_;
  assign N1367 = ~pe_o_2__5_;
  assign N1368 = ~pe_o_2__1_;
  assign N1369 = N1374 & N1375;
  assign N1370 = N1369 & pe_o_2__4_;
  assign N1371 = N1370 & pe_o_2__3_;
  assign N1372 = N1371 & pe_o_2__2_;
  assign N1373 = N1372 & N1376;
  assign N7615 = N1373 & pe_o_2__1_;
  assign N1374 = ~pe_o_2__6_;
  assign N1375 = ~pe_o_2__5_;
  assign N1376 = ~pe_o_2__0_;
  assign N1377 = N1382 & N1383;
  assign N1378 = N1377 & pe_o_2__4_;
  assign N1379 = N1378 & pe_o_2__3_;
  assign N1380 = N1379 & pe_o_2__2_;
  assign N1381 = N1380 & pe_o_2__0_;
  assign N7617 = N1381 & pe_o_2__1_;
  assign N1382 = ~pe_o_2__6_;
  assign N1383 = ~pe_o_2__5_;
  assign N1384 = N1389 & pe_o_2__5_;
  assign N1385 = N1384 & N1390;
  assign N1386 = N1385 & N1391;
  assign N1387 = N1386 & N1392;
  assign N1388 = N1387 & N1393;
  assign N7619 = N1388 & N1394;
  assign N1389 = ~pe_o_2__6_;
  assign N1390 = ~pe_o_2__4_;
  assign N1391 = ~pe_o_2__3_;
  assign N1392 = ~pe_o_2__2_;
  assign N1393 = ~pe_o_2__0_;
  assign N1394 = ~pe_o_2__1_;
  assign N1395 = N1400 & pe_o_2__5_;
  assign N1396 = N1395 & N1401;
  assign N1397 = N1396 & N1402;
  assign N1398 = N1397 & N1403;
  assign N1399 = N1398 & pe_o_2__0_;
  assign N7621 = N1399 & N1404;
  assign N1400 = ~pe_o_2__6_;
  assign N1401 = ~pe_o_2__4_;
  assign N1402 = ~pe_o_2__3_;
  assign N1403 = ~pe_o_2__2_;
  assign N1404 = ~pe_o_2__1_;
  assign N1405 = N1410 & pe_o_2__5_;
  assign N1406 = N1405 & N1411;
  assign N1407 = N1406 & N1412;
  assign N1408 = N1407 & N1413;
  assign N1409 = N1408 & N1414;
  assign N7623 = N1409 & pe_o_2__1_;
  assign N1410 = ~pe_o_2__6_;
  assign N1411 = ~pe_o_2__4_;
  assign N1412 = ~pe_o_2__3_;
  assign N1413 = ~pe_o_2__2_;
  assign N1414 = ~pe_o_2__0_;
  assign N1415 = N1420 & pe_o_2__5_;
  assign N1416 = N1415 & N1421;
  assign N1417 = N1416 & N1422;
  assign N1418 = N1417 & N1423;
  assign N1419 = N1418 & pe_o_2__0_;
  assign N7625 = N1419 & pe_o_2__1_;
  assign N1420 = ~pe_o_2__6_;
  assign N1421 = ~pe_o_2__4_;
  assign N1422 = ~pe_o_2__3_;
  assign N1423 = ~pe_o_2__2_;
  assign N1424 = N1429 & pe_o_2__5_;
  assign N1425 = N1424 & N1430;
  assign N1426 = N1425 & N1431;
  assign N1427 = N1426 & pe_o_2__2_;
  assign N1428 = N1427 & N1432;
  assign N7627 = N1428 & N1433;
  assign N1429 = ~pe_o_2__6_;
  assign N1430 = ~pe_o_2__4_;
  assign N1431 = ~pe_o_2__3_;
  assign N1432 = ~pe_o_2__0_;
  assign N1433 = ~pe_o_2__1_;
  assign N1434 = N1439 & pe_o_2__5_;
  assign N1435 = N1434 & N1440;
  assign N1436 = N1435 & N1441;
  assign N1437 = N1436 & pe_o_2__2_;
  assign N1438 = N1437 & pe_o_2__0_;
  assign N7629 = N1438 & N1442;
  assign N1439 = ~pe_o_2__6_;
  assign N1440 = ~pe_o_2__4_;
  assign N1441 = ~pe_o_2__3_;
  assign N1442 = ~pe_o_2__1_;
  assign N1443 = N1448 & pe_o_2__5_;
  assign N1444 = N1443 & N1449;
  assign N1445 = N1444 & N1450;
  assign N1446 = N1445 & pe_o_2__2_;
  assign N1447 = N1446 & N1451;
  assign N7631 = N1447 & pe_o_2__1_;
  assign N1448 = ~pe_o_2__6_;
  assign N1449 = ~pe_o_2__4_;
  assign N1450 = ~pe_o_2__3_;
  assign N1451 = ~pe_o_2__0_;
  assign N1452 = N1457 & pe_o_2__5_;
  assign N1453 = N1452 & N1458;
  assign N1454 = N1453 & N1459;
  assign N1455 = N1454 & pe_o_2__2_;
  assign N1456 = N1455 & pe_o_2__0_;
  assign N7633 = N1456 & pe_o_2__1_;
  assign N1457 = ~pe_o_2__6_;
  assign N1458 = ~pe_o_2__4_;
  assign N1459 = ~pe_o_2__3_;
  assign N1460 = N1465 & pe_o_2__5_;
  assign N1461 = N1460 & N1466;
  assign N1462 = N1461 & pe_o_2__3_;
  assign N1463 = N1462 & N1467;
  assign N1464 = N1463 & N1468;
  assign N7635 = N1464 & N1469;
  assign N1465 = ~pe_o_2__6_;
  assign N1466 = ~pe_o_2__4_;
  assign N1467 = ~pe_o_2__2_;
  assign N1468 = ~pe_o_2__0_;
  assign N1469 = ~pe_o_2__1_;
  assign N1470 = N1475 & pe_o_2__5_;
  assign N1471 = N1470 & N1476;
  assign N1472 = N1471 & pe_o_2__3_;
  assign N1473 = N1472 & N1477;
  assign N1474 = N1473 & pe_o_2__0_;
  assign N7637 = N1474 & N1478;
  assign N1475 = ~pe_o_2__6_;
  assign N1476 = ~pe_o_2__4_;
  assign N1477 = ~pe_o_2__2_;
  assign N1478 = ~pe_o_2__1_;
  assign N1479 = N1484 & pe_o_2__5_;
  assign N1480 = N1479 & N1485;
  assign N1481 = N1480 & pe_o_2__3_;
  assign N1482 = N1481 & N1486;
  assign N1483 = N1482 & N1487;
  assign N7639 = N1483 & pe_o_2__1_;
  assign N1484 = ~pe_o_2__6_;
  assign N1485 = ~pe_o_2__4_;
  assign N1486 = ~pe_o_2__2_;
  assign N1487 = ~pe_o_2__0_;
  assign N1488 = N1493 & pe_o_2__5_;
  assign N1489 = N1488 & N1494;
  assign N1490 = N1489 & pe_o_2__3_;
  assign N1491 = N1490 & N1495;
  assign N1492 = N1491 & pe_o_2__0_;
  assign N7641 = N1492 & pe_o_2__1_;
  assign N1493 = ~pe_o_2__6_;
  assign N1494 = ~pe_o_2__4_;
  assign N1495 = ~pe_o_2__2_;
  assign N1496 = N1501 & pe_o_2__5_;
  assign N1497 = N1496 & N1502;
  assign N1498 = N1497 & pe_o_2__3_;
  assign N1499 = N1498 & pe_o_2__2_;
  assign N1500 = N1499 & N1503;
  assign N7643 = N1500 & N1504;
  assign N1501 = ~pe_o_2__6_;
  assign N1502 = ~pe_o_2__4_;
  assign N1503 = ~pe_o_2__0_;
  assign N1504 = ~pe_o_2__1_;
  assign N1505 = N1510 & pe_o_2__5_;
  assign N1506 = N1505 & N1511;
  assign N1507 = N1506 & pe_o_2__3_;
  assign N1508 = N1507 & pe_o_2__2_;
  assign N1509 = N1508 & pe_o_2__0_;
  assign N7645 = N1509 & N1512;
  assign N1510 = ~pe_o_2__6_;
  assign N1511 = ~pe_o_2__4_;
  assign N1512 = ~pe_o_2__1_;
  assign N1513 = N1518 & pe_o_2__5_;
  assign N1514 = N1513 & N1519;
  assign N1515 = N1514 & pe_o_2__3_;
  assign N1516 = N1515 & pe_o_2__2_;
  assign N1517 = N1516 & N1520;
  assign N7647 = N1517 & pe_o_2__1_;
  assign N1518 = ~pe_o_2__6_;
  assign N1519 = ~pe_o_2__4_;
  assign N1520 = ~pe_o_2__0_;
  assign N1521 = N1526 & pe_o_2__5_;
  assign N1522 = N1521 & N1527;
  assign N1523 = N1522 & pe_o_2__3_;
  assign N1524 = N1523 & pe_o_2__2_;
  assign N1525 = N1524 & pe_o_2__0_;
  assign N7649 = N1525 & pe_o_2__1_;
  assign N1526 = ~pe_o_2__6_;
  assign N1527 = ~pe_o_2__4_;
  assign N1528 = N1533 & pe_o_2__5_;
  assign N1529 = N1528 & pe_o_2__4_;
  assign N1530 = N1529 & N1534;
  assign N1531 = N1530 & N1535;
  assign N1532 = N1531 & N1536;
  assign N7651 = N1532 & N1537;
  assign N1533 = ~pe_o_2__6_;
  assign N1534 = ~pe_o_2__3_;
  assign N1535 = ~pe_o_2__2_;
  assign N1536 = ~pe_o_2__0_;
  assign N1537 = ~pe_o_2__1_;
  assign N1538 = N1543 & pe_o_2__5_;
  assign N1539 = N1538 & pe_o_2__4_;
  assign N1540 = N1539 & N1544;
  assign N1541 = N1540 & N1545;
  assign N1542 = N1541 & pe_o_2__0_;
  assign N7653 = N1542 & N1546;
  assign N1543 = ~pe_o_2__6_;
  assign N1544 = ~pe_o_2__3_;
  assign N1545 = ~pe_o_2__2_;
  assign N1546 = ~pe_o_2__1_;
  assign N1547 = N1552 & pe_o_2__5_;
  assign N1548 = N1547 & pe_o_2__4_;
  assign N1549 = N1548 & N1553;
  assign N1550 = N1549 & N1554;
  assign N1551 = N1550 & N1555;
  assign N7655 = N1551 & pe_o_2__1_;
  assign N1552 = ~pe_o_2__6_;
  assign N1553 = ~pe_o_2__3_;
  assign N1554 = ~pe_o_2__2_;
  assign N1555 = ~pe_o_2__0_;
  assign N1556 = N1561 & pe_o_2__5_;
  assign N1557 = N1556 & pe_o_2__4_;
  assign N1558 = N1557 & N1562;
  assign N1559 = N1558 & N1563;
  assign N1560 = N1559 & pe_o_2__0_;
  assign N7657 = N1560 & pe_o_2__1_;
  assign N1561 = ~pe_o_2__6_;
  assign N1562 = ~pe_o_2__3_;
  assign N1563 = ~pe_o_2__2_;
  assign N1564 = N1569 & pe_o_2__5_;
  assign N1565 = N1564 & pe_o_2__4_;
  assign N1566 = N1565 & N1570;
  assign N1567 = N1566 & pe_o_2__2_;
  assign N1568 = N1567 & N1571;
  assign N7659 = N1568 & N1572;
  assign N1569 = ~pe_o_2__6_;
  assign N1570 = ~pe_o_2__3_;
  assign N1571 = ~pe_o_2__0_;
  assign N1572 = ~pe_o_2__1_;
  assign N1573 = N1578 & pe_o_2__5_;
  assign N1574 = N1573 & pe_o_2__4_;
  assign N1575 = N1574 & N1579;
  assign N1576 = N1575 & pe_o_2__2_;
  assign N1577 = N1576 & pe_o_2__0_;
  assign N7661 = N1577 & N1580;
  assign N1578 = ~pe_o_2__6_;
  assign N1579 = ~pe_o_2__3_;
  assign N1580 = ~pe_o_2__1_;
  assign N1581 = N1586 & pe_o_2__5_;
  assign N1582 = N1581 & pe_o_2__4_;
  assign N1583 = N1582 & N1587;
  assign N1584 = N1583 & pe_o_2__2_;
  assign N1585 = N1584 & N1588;
  assign N7663 = N1585 & pe_o_2__1_;
  assign N1586 = ~pe_o_2__6_;
  assign N1587 = ~pe_o_2__3_;
  assign N1588 = ~pe_o_2__0_;
  assign N1589 = N1594 & pe_o_2__5_;
  assign N1590 = N1589 & pe_o_2__4_;
  assign N1591 = N1590 & N1595;
  assign N1592 = N1591 & pe_o_2__2_;
  assign N1593 = N1592 & pe_o_2__0_;
  assign N7665 = N1593 & pe_o_2__1_;
  assign N1594 = ~pe_o_2__6_;
  assign N1595 = ~pe_o_2__3_;
  assign N1596 = N1601 & pe_o_2__5_;
  assign N1597 = N1596 & pe_o_2__4_;
  assign N1598 = N1597 & pe_o_2__3_;
  assign N1599 = N1598 & N1602;
  assign N1600 = N1599 & N1603;
  assign N7667 = N1600 & N1604;
  assign N1601 = ~pe_o_2__6_;
  assign N1602 = ~pe_o_2__2_;
  assign N1603 = ~pe_o_2__0_;
  assign N1604 = ~pe_o_2__1_;
  assign N1605 = N1610 & pe_o_2__5_;
  assign N1606 = N1605 & pe_o_2__4_;
  assign N1607 = N1606 & pe_o_2__3_;
  assign N1608 = N1607 & N1611;
  assign N1609 = N1608 & pe_o_2__0_;
  assign N7669 = N1609 & N1612;
  assign N1610 = ~pe_o_2__6_;
  assign N1611 = ~pe_o_2__2_;
  assign N1612 = ~pe_o_2__1_;
  assign N1613 = N1618 & pe_o_2__5_;
  assign N1614 = N1613 & pe_o_2__4_;
  assign N1615 = N1614 & pe_o_2__3_;
  assign N1616 = N1615 & N1619;
  assign N1617 = N1616 & N1620;
  assign N7671 = N1617 & pe_o_2__1_;
  assign N1618 = ~pe_o_2__6_;
  assign N1619 = ~pe_o_2__2_;
  assign N1620 = ~pe_o_2__0_;
  assign N1621 = N1626 & pe_o_2__5_;
  assign N1622 = N1621 & pe_o_2__4_;
  assign N1623 = N1622 & pe_o_2__3_;
  assign N1624 = N1623 & N1627;
  assign N1625 = N1624 & pe_o_2__0_;
  assign N7673 = N1625 & pe_o_2__1_;
  assign N1626 = ~pe_o_2__6_;
  assign N1627 = ~pe_o_2__2_;
  assign N1628 = N1633 & pe_o_2__5_;
  assign N1629 = N1628 & pe_o_2__4_;
  assign N1630 = N1629 & pe_o_2__3_;
  assign N1631 = N1630 & pe_o_2__2_;
  assign N1632 = N1631 & N1634;
  assign N7675 = N1632 & N1635;
  assign N1633 = ~pe_o_2__6_;
  assign N1634 = ~pe_o_2__0_;
  assign N1635 = ~pe_o_2__1_;
  assign N1636 = N1641 & pe_o_2__5_;
  assign N1637 = N1636 & pe_o_2__4_;
  assign N1638 = N1637 & pe_o_2__3_;
  assign N1639 = N1638 & pe_o_2__2_;
  assign N1640 = N1639 & pe_o_2__0_;
  assign N7677 = N1640 & N1642;
  assign N1641 = ~pe_o_2__6_;
  assign N1642 = ~pe_o_2__1_;
  assign N1643 = N1648 & pe_o_2__5_;
  assign N1644 = N1643 & pe_o_2__4_;
  assign N1645 = N1644 & pe_o_2__3_;
  assign N1646 = N1645 & pe_o_2__2_;
  assign N1647 = N1646 & N1649;
  assign N7679 = N1647 & pe_o_2__1_;
  assign N1648 = ~pe_o_2__6_;
  assign N1649 = ~pe_o_2__0_;
  assign N1650 = pe_o_2__5_ & pe_o_2__4_;
  assign N1651 = N1650 & pe_o_2__3_;
  assign N1652 = N1651 & pe_o_2__2_;
  assign N1653 = N1652 & pe_o_2__0_;
  assign N7681 = N1653 & pe_o_2__1_;
  assign N1654 = pe_o_2__6_ & N1659;
  assign N1655 = N1654 & N1660;
  assign N1656 = N1655 & N1661;
  assign N1657 = N1656 & N1662;
  assign N1658 = N1657 & pe_o_2__0_;
  assign N7558 = N1658 & N1663;
  assign N1659 = ~pe_o_2__5_;
  assign N1660 = ~pe_o_2__4_;
  assign N1661 = ~pe_o_2__3_;
  assign N1662 = ~pe_o_2__2_;
  assign N1663 = ~pe_o_2__1_;
  assign N1664 = pe_o_2__6_ & N1669;
  assign N1665 = N1664 & N1670;
  assign N1666 = N1665 & N1671;
  assign N1667 = N1666 & N1672;
  assign N1668 = N1667 & N1673;
  assign N7560 = N1668 & pe_o_2__1_;
  assign N1669 = ~pe_o_2__5_;
  assign N1670 = ~pe_o_2__4_;
  assign N1671 = ~pe_o_2__3_;
  assign N1672 = ~pe_o_2__2_;
  assign N1673 = ~pe_o_2__0_;
  assign N1674 = pe_o_2__6_ & N1679;
  assign N1675 = N1674 & N1680;
  assign N1676 = N1675 & N1681;
  assign N1677 = N1676 & N1682;
  assign N1678 = N1677 & pe_o_2__0_;
  assign N7562 = N1678 & pe_o_2__1_;
  assign N1679 = ~pe_o_2__5_;
  assign N1680 = ~pe_o_2__4_;
  assign N1681 = ~pe_o_2__3_;
  assign N1682 = ~pe_o_2__2_;
  assign N1683 = pe_o_2__6_ & N1688;
  assign N1684 = N1683 & N1689;
  assign N1685 = N1684 & N1690;
  assign N1686 = N1685 & pe_o_2__2_;
  assign N1687 = N1686 & N1691;
  assign N7564 = N1687 & N1692;
  assign N1688 = ~pe_o_2__5_;
  assign N1689 = ~pe_o_2__4_;
  assign N1690 = ~pe_o_2__3_;
  assign N1691 = ~pe_o_2__0_;
  assign N1692 = ~pe_o_2__1_;
  assign N1693 = pe_o_2__6_ & N1698;
  assign N1694 = N1693 & N1699;
  assign N1695 = N1694 & N1700;
  assign N1696 = N1695 & pe_o_2__2_;
  assign N1697 = N1696 & pe_o_2__0_;
  assign N7566 = N1697 & N1701;
  assign N1698 = ~pe_o_2__5_;
  assign N1699 = ~pe_o_2__4_;
  assign N1700 = ~pe_o_2__3_;
  assign N1701 = ~pe_o_2__1_;
  assign N1702 = pe_o_2__6_ & N1707;
  assign N1703 = N1702 & N1708;
  assign N1704 = N1703 & N1709;
  assign N1705 = N1704 & pe_o_2__2_;
  assign N1706 = N1705 & N1710;
  assign N7568 = N1706 & pe_o_2__1_;
  assign N1707 = ~pe_o_2__5_;
  assign N1708 = ~pe_o_2__4_;
  assign N1709 = ~pe_o_2__3_;
  assign N1710 = ~pe_o_2__0_;
  assign N1711 = pe_o_2__6_ & N1716;
  assign N1712 = N1711 & N1717;
  assign N1713 = N1712 & N1718;
  assign N1714 = N1713 & pe_o_2__2_;
  assign N1715 = N1714 & pe_o_2__0_;
  assign N7570 = N1715 & pe_o_2__1_;
  assign N1716 = ~pe_o_2__5_;
  assign N1717 = ~pe_o_2__4_;
  assign N1718 = ~pe_o_2__3_;
  assign N1719 = pe_o_2__6_ & N1724;
  assign N1720 = N1719 & N1725;
  assign N1721 = N1720 & pe_o_2__3_;
  assign N1722 = N1721 & N1726;
  assign N1723 = N1722 & N1727;
  assign N7572 = N1723 & N1728;
  assign N1724 = ~pe_o_2__5_;
  assign N1725 = ~pe_o_2__4_;
  assign N1726 = ~pe_o_2__2_;
  assign N1727 = ~pe_o_2__0_;
  assign N1728 = ~pe_o_2__1_;
  assign N1729 = pe_o_2__6_ & N1734;
  assign N1730 = N1729 & N1735;
  assign N1731 = N1730 & pe_o_2__3_;
  assign N1732 = N1731 & N1736;
  assign N1733 = N1732 & pe_o_2__0_;
  assign N7574 = N1733 & N1737;
  assign N1734 = ~pe_o_2__5_;
  assign N1735 = ~pe_o_2__4_;
  assign N1736 = ~pe_o_2__2_;
  assign N1737 = ~pe_o_2__1_;
  assign N1738 = pe_o_2__6_ & N1743;
  assign N1739 = N1738 & N1744;
  assign N1740 = N1739 & pe_o_2__3_;
  assign N1741 = N1740 & N1745;
  assign N1742 = N1741 & N1746;
  assign N7576 = N1742 & pe_o_2__1_;
  assign N1743 = ~pe_o_2__5_;
  assign N1744 = ~pe_o_2__4_;
  assign N1745 = ~pe_o_2__2_;
  assign N1746 = ~pe_o_2__0_;
  assign N1747 = pe_o_2__6_ & N1752;
  assign N1748 = N1747 & N1753;
  assign N1749 = N1748 & pe_o_2__3_;
  assign N1750 = N1749 & N1754;
  assign N1751 = N1750 & pe_o_2__0_;
  assign N7578 = N1751 & pe_o_2__1_;
  assign N1752 = ~pe_o_2__5_;
  assign N1753 = ~pe_o_2__4_;
  assign N1754 = ~pe_o_2__2_;
  assign N1755 = pe_o_2__6_ & N1760;
  assign N1756 = N1755 & N1761;
  assign N1757 = N1756 & pe_o_2__3_;
  assign N1758 = N1757 & pe_o_2__2_;
  assign N1759 = N1758 & N1762;
  assign N7580 = N1759 & N1763;
  assign N1760 = ~pe_o_2__5_;
  assign N1761 = ~pe_o_2__4_;
  assign N1762 = ~pe_o_2__0_;
  assign N1763 = ~pe_o_2__1_;
  assign N1764 = pe_o_2__6_ & N1769;
  assign N1765 = N1764 & N1770;
  assign N1766 = N1765 & pe_o_2__3_;
  assign N1767 = N1766 & pe_o_2__2_;
  assign N1768 = N1767 & pe_o_2__0_;
  assign N7582 = N1768 & N1771;
  assign N1769 = ~pe_o_2__5_;
  assign N1770 = ~pe_o_2__4_;
  assign N1771 = ~pe_o_2__1_;
  assign N1772 = pe_o_2__6_ & N1777;
  assign N1773 = N1772 & N1778;
  assign N1774 = N1773 & pe_o_2__3_;
  assign N1775 = N1774 & pe_o_2__2_;
  assign N1776 = N1775 & N1779;
  assign N7584 = N1776 & pe_o_2__1_;
  assign N1777 = ~pe_o_2__5_;
  assign N1778 = ~pe_o_2__4_;
  assign N1779 = ~pe_o_2__0_;
  assign N1780 = pe_o_2__6_ & N1785;
  assign N1781 = N1780 & N1786;
  assign N1782 = N1781 & pe_o_2__3_;
  assign N1783 = N1782 & pe_o_2__2_;
  assign N1784 = N1783 & pe_o_2__0_;
  assign N7586 = N1784 & pe_o_2__1_;
  assign N1785 = ~pe_o_2__5_;
  assign N1786 = ~pe_o_2__4_;
  assign N1787 = pe_o_2__6_ & N1792;
  assign N1788 = N1787 & pe_o_2__4_;
  assign N1789 = N1788 & N1793;
  assign N1790 = N1789 & N1794;
  assign N1791 = N1790 & N1795;
  assign N7588 = N1791 & N1796;
  assign N1792 = ~pe_o_2__5_;
  assign N1793 = ~pe_o_2__3_;
  assign N1794 = ~pe_o_2__2_;
  assign N1795 = ~pe_o_2__0_;
  assign N1796 = ~pe_o_2__1_;
  assign N1797 = pe_o_2__6_ & N1802;
  assign N1798 = N1797 & pe_o_2__4_;
  assign N1799 = N1798 & N1803;
  assign N1800 = N1799 & N1804;
  assign N1801 = N1800 & pe_o_2__0_;
  assign N7590 = N1801 & N1805;
  assign N1802 = ~pe_o_2__5_;
  assign N1803 = ~pe_o_2__3_;
  assign N1804 = ~pe_o_2__2_;
  assign N1805 = ~pe_o_2__1_;
  assign N1806 = pe_o_2__6_ & N1811;
  assign N1807 = N1806 & pe_o_2__4_;
  assign N1808 = N1807 & N1812;
  assign N1809 = N1808 & N1813;
  assign N1810 = N1809 & N1814;
  assign N7592 = N1810 & pe_o_2__1_;
  assign N1811 = ~pe_o_2__5_;
  assign N1812 = ~pe_o_2__3_;
  assign N1813 = ~pe_o_2__2_;
  assign N1814 = ~pe_o_2__0_;
  assign N1815 = pe_o_2__6_ & N1820;
  assign N1816 = N1815 & pe_o_2__4_;
  assign N1817 = N1816 & N1821;
  assign N1818 = N1817 & N1822;
  assign N1819 = N1818 & pe_o_2__0_;
  assign N7594 = N1819 & pe_o_2__1_;
  assign N1820 = ~pe_o_2__5_;
  assign N1821 = ~pe_o_2__3_;
  assign N1822 = ~pe_o_2__2_;
  assign N1823 = pe_o_2__6_ & N1828;
  assign N1824 = N1823 & pe_o_2__4_;
  assign N1825 = N1824 & N1829;
  assign N1826 = N1825 & pe_o_2__2_;
  assign N1827 = N1826 & N1830;
  assign N7596 = N1827 & N1831;
  assign N1828 = ~pe_o_2__5_;
  assign N1829 = ~pe_o_2__3_;
  assign N1830 = ~pe_o_2__0_;
  assign N1831 = ~pe_o_2__1_;
  assign N1832 = pe_o_2__6_ & N1837;
  assign N1833 = N1832 & pe_o_2__4_;
  assign N1834 = N1833 & N1838;
  assign N1835 = N1834 & pe_o_2__2_;
  assign N1836 = N1835 & pe_o_2__0_;
  assign N7598 = N1836 & N1839;
  assign N1837 = ~pe_o_2__5_;
  assign N1838 = ~pe_o_2__3_;
  assign N1839 = ~pe_o_2__1_;
  assign N1840 = pe_o_2__6_ & N1845;
  assign N1841 = N1840 & pe_o_2__4_;
  assign N1842 = N1841 & N1846;
  assign N1843 = N1842 & pe_o_2__2_;
  assign N1844 = N1843 & N1847;
  assign N7600 = N1844 & pe_o_2__1_;
  assign N1845 = ~pe_o_2__5_;
  assign N1846 = ~pe_o_2__3_;
  assign N1847 = ~pe_o_2__0_;
  assign N1848 = pe_o_2__6_ & N1853;
  assign N1849 = N1848 & pe_o_2__4_;
  assign N1850 = N1849 & N1854;
  assign N1851 = N1850 & pe_o_2__2_;
  assign N1852 = N1851 & pe_o_2__0_;
  assign N7602 = N1852 & pe_o_2__1_;
  assign N1853 = ~pe_o_2__5_;
  assign N1854 = ~pe_o_2__3_;
  assign N1855 = pe_o_2__6_ & N1860;
  assign N1856 = N1855 & pe_o_2__4_;
  assign N1857 = N1856 & pe_o_2__3_;
  assign N1858 = N1857 & N1861;
  assign N1859 = N1858 & N1862;
  assign N7604 = N1859 & N1863;
  assign N1860 = ~pe_o_2__5_;
  assign N1861 = ~pe_o_2__2_;
  assign N1862 = ~pe_o_2__0_;
  assign N1863 = ~pe_o_2__1_;
  assign N1864 = pe_o_2__6_ & N1869;
  assign N1865 = N1864 & pe_o_2__4_;
  assign N1866 = N1865 & pe_o_2__3_;
  assign N1867 = N1866 & N1870;
  assign N1868 = N1867 & pe_o_2__0_;
  assign N7606 = N1868 & N1871;
  assign N1869 = ~pe_o_2__5_;
  assign N1870 = ~pe_o_2__2_;
  assign N1871 = ~pe_o_2__1_;
  assign N1872 = pe_o_2__6_ & N1877;
  assign N1873 = N1872 & pe_o_2__4_;
  assign N1874 = N1873 & pe_o_2__3_;
  assign N1875 = N1874 & N1878;
  assign N1876 = N1875 & N1879;
  assign N7608 = N1876 & pe_o_2__1_;
  assign N1877 = ~pe_o_2__5_;
  assign N1878 = ~pe_o_2__2_;
  assign N1879 = ~pe_o_2__0_;
  assign N1880 = pe_o_2__6_ & N1885;
  assign N1881 = N1880 & pe_o_2__4_;
  assign N1882 = N1881 & pe_o_2__3_;
  assign N1883 = N1882 & N1886;
  assign N1884 = N1883 & pe_o_2__0_;
  assign N7610 = N1884 & pe_o_2__1_;
  assign N1885 = ~pe_o_2__5_;
  assign N1886 = ~pe_o_2__2_;
  assign N1887 = pe_o_2__6_ & N1892;
  assign N1888 = N1887 & pe_o_2__4_;
  assign N1889 = N1888 & pe_o_2__3_;
  assign N1890 = N1889 & pe_o_2__2_;
  assign N1891 = N1890 & N1893;
  assign N7612 = N1891 & N1894;
  assign N1892 = ~pe_o_2__5_;
  assign N1893 = ~pe_o_2__0_;
  assign N1894 = ~pe_o_2__1_;
  assign N1895 = pe_o_2__6_ & N1900;
  assign N1896 = N1895 & pe_o_2__4_;
  assign N1897 = N1896 & pe_o_2__3_;
  assign N1898 = N1897 & pe_o_2__2_;
  assign N1899 = N1898 & pe_o_2__0_;
  assign N7614 = N1899 & N1901;
  assign N1900 = ~pe_o_2__5_;
  assign N1901 = ~pe_o_2__1_;
  assign N1902 = pe_o_2__6_ & N1907;
  assign N1903 = N1902 & pe_o_2__4_;
  assign N1904 = N1903 & pe_o_2__3_;
  assign N1905 = N1904 & pe_o_2__2_;
  assign N1906 = N1905 & N1908;
  assign N7616 = N1906 & pe_o_2__1_;
  assign N1907 = ~pe_o_2__5_;
  assign N1908 = ~pe_o_2__0_;
  assign N1909 = pe_o_2__6_ & pe_o_2__4_;
  assign N1910 = N1909 & pe_o_2__3_;
  assign N1911 = N1910 & pe_o_2__2_;
  assign N1912 = N1911 & pe_o_2__0_;
  assign N7618 = N1912 & pe_o_2__1_;
  assign N1913 = pe_o_2__6_ & pe_o_2__5_;
  assign N1914 = N1913 & N1918;
  assign N1915 = N1914 & N1919;
  assign N1916 = N1915 & N1920;
  assign N1917 = N1916 & N1921;
  assign N7620 = N1917 & N1922;
  assign N1918 = ~pe_o_2__4_;
  assign N1919 = ~pe_o_2__3_;
  assign N1920 = ~pe_o_2__2_;
  assign N1921 = ~pe_o_2__0_;
  assign N1922 = ~pe_o_2__1_;
  assign N1923 = pe_o_2__6_ & pe_o_2__5_;
  assign N1924 = N1923 & N1928;
  assign N1925 = N1924 & N1929;
  assign N1926 = N1925 & N1930;
  assign N1927 = N1926 & pe_o_2__0_;
  assign N7622 = N1927 & N1931;
  assign N1928 = ~pe_o_2__4_;
  assign N1929 = ~pe_o_2__3_;
  assign N1930 = ~pe_o_2__2_;
  assign N1931 = ~pe_o_2__1_;
  assign N1932 = pe_o_2__6_ & pe_o_2__5_;
  assign N1933 = N1932 & N1937;
  assign N1934 = N1933 & N1938;
  assign N1935 = N1934 & N1939;
  assign N1936 = N1935 & N1940;
  assign N7624 = N1936 & pe_o_2__1_;
  assign N1937 = ~pe_o_2__4_;
  assign N1938 = ~pe_o_2__3_;
  assign N1939 = ~pe_o_2__2_;
  assign N1940 = ~pe_o_2__0_;
  assign N1941 = pe_o_2__6_ & pe_o_2__5_;
  assign N1942 = N1941 & N1946;
  assign N1943 = N1942 & N1947;
  assign N1944 = N1943 & N1948;
  assign N1945 = N1944 & pe_o_2__0_;
  assign N7626 = N1945 & pe_o_2__1_;
  assign N1946 = ~pe_o_2__4_;
  assign N1947 = ~pe_o_2__3_;
  assign N1948 = ~pe_o_2__2_;
  assign N1949 = pe_o_2__6_ & pe_o_2__5_;
  assign N1950 = N1949 & N1954;
  assign N1951 = N1950 & N1955;
  assign N1952 = N1951 & pe_o_2__2_;
  assign N1953 = N1952 & N1956;
  assign N7628 = N1953 & N1957;
  assign N1954 = ~pe_o_2__4_;
  assign N1955 = ~pe_o_2__3_;
  assign N1956 = ~pe_o_2__0_;
  assign N1957 = ~pe_o_2__1_;
  assign N1958 = pe_o_2__6_ & pe_o_2__5_;
  assign N1959 = N1958 & N1963;
  assign N1960 = N1959 & N1964;
  assign N1961 = N1960 & pe_o_2__2_;
  assign N1962 = N1961 & pe_o_2__0_;
  assign N7630 = N1962 & N1965;
  assign N1963 = ~pe_o_2__4_;
  assign N1964 = ~pe_o_2__3_;
  assign N1965 = ~pe_o_2__1_;
  assign N1966 = pe_o_2__6_ & pe_o_2__5_;
  assign N1967 = N1966 & N1971;
  assign N1968 = N1967 & N1972;
  assign N1969 = N1968 & pe_o_2__2_;
  assign N1970 = N1969 & N1973;
  assign N7632 = N1970 & pe_o_2__1_;
  assign N1971 = ~pe_o_2__4_;
  assign N1972 = ~pe_o_2__3_;
  assign N1973 = ~pe_o_2__0_;
  assign N1974 = pe_o_2__6_ & pe_o_2__5_;
  assign N1975 = N1974 & N1979;
  assign N1976 = N1975 & N1980;
  assign N1977 = N1976 & pe_o_2__2_;
  assign N1978 = N1977 & pe_o_2__0_;
  assign N7634 = N1978 & pe_o_2__1_;
  assign N1979 = ~pe_o_2__4_;
  assign N1980 = ~pe_o_2__3_;
  assign N1981 = pe_o_2__6_ & pe_o_2__5_;
  assign N1982 = N1981 & N1986;
  assign N1983 = N1982 & pe_o_2__3_;
  assign N1984 = N1983 & N1987;
  assign N1985 = N1984 & N1988;
  assign N7636 = N1985 & N1989;
  assign N1986 = ~pe_o_2__4_;
  assign N1987 = ~pe_o_2__2_;
  assign N1988 = ~pe_o_2__0_;
  assign N1989 = ~pe_o_2__1_;
  assign N1990 = pe_o_2__6_ & pe_o_2__5_;
  assign N1991 = N1990 & N1995;
  assign N1992 = N1991 & pe_o_2__3_;
  assign N1993 = N1992 & N1996;
  assign N1994 = N1993 & pe_o_2__0_;
  assign N7638 = N1994 & N1997;
  assign N1995 = ~pe_o_2__4_;
  assign N1996 = ~pe_o_2__2_;
  assign N1997 = ~pe_o_2__1_;
  assign N1998 = pe_o_2__6_ & pe_o_2__5_;
  assign N1999 = N1998 & N2003;
  assign N2000 = N1999 & pe_o_2__3_;
  assign N2001 = N2000 & N2004;
  assign N2002 = N2001 & N2005;
  assign N7640 = N2002 & pe_o_2__1_;
  assign N2003 = ~pe_o_2__4_;
  assign N2004 = ~pe_o_2__2_;
  assign N2005 = ~pe_o_2__0_;
  assign N2006 = pe_o_2__6_ & pe_o_2__5_;
  assign N2007 = N2006 & N2011;
  assign N2008 = N2007 & pe_o_2__3_;
  assign N2009 = N2008 & N2012;
  assign N2010 = N2009 & pe_o_2__0_;
  assign N7642 = N2010 & pe_o_2__1_;
  assign N2011 = ~pe_o_2__4_;
  assign N2012 = ~pe_o_2__2_;
  assign N2013 = pe_o_2__6_ & pe_o_2__5_;
  assign N2014 = N2013 & N2018;
  assign N2015 = N2014 & pe_o_2__3_;
  assign N2016 = N2015 & pe_o_2__2_;
  assign N2017 = N2016 & N2019;
  assign N7644 = N2017 & N2020;
  assign N2018 = ~pe_o_2__4_;
  assign N2019 = ~pe_o_2__0_;
  assign N2020 = ~pe_o_2__1_;
  assign N2021 = pe_o_2__6_ & pe_o_2__5_;
  assign N2022 = N2021 & N2026;
  assign N2023 = N2022 & pe_o_2__3_;
  assign N2024 = N2023 & pe_o_2__2_;
  assign N2025 = N2024 & pe_o_2__0_;
  assign N7646 = N2025 & N2027;
  assign N2026 = ~pe_o_2__4_;
  assign N2027 = ~pe_o_2__1_;
  assign N2028 = pe_o_2__6_ & pe_o_2__5_;
  assign N2029 = N2028 & N2033;
  assign N2030 = N2029 & pe_o_2__3_;
  assign N2031 = N2030 & pe_o_2__2_;
  assign N2032 = N2031 & N2034;
  assign N7648 = N2032 & pe_o_2__1_;
  assign N2033 = ~pe_o_2__4_;
  assign N2034 = ~pe_o_2__0_;
  assign N2035 = pe_o_2__6_ & pe_o_2__5_;
  assign N2036 = N2035 & pe_o_2__3_;
  assign N2037 = N2036 & pe_o_2__2_;
  assign N2038 = N2037 & pe_o_2__0_;
  assign N7650 = N2038 & pe_o_2__1_;
  assign N2039 = pe_o_2__6_ & pe_o_2__5_;
  assign N2040 = N2039 & pe_o_2__4_;
  assign N2041 = N2040 & N2044;
  assign N2042 = N2041 & N2045;
  assign N2043 = N2042 & N2046;
  assign N7652 = N2043 & N2047;
  assign N2044 = ~pe_o_2__3_;
  assign N2045 = ~pe_o_2__2_;
  assign N2046 = ~pe_o_2__0_;
  assign N2047 = ~pe_o_2__1_;
  assign N2048 = pe_o_2__6_ & pe_o_2__5_;
  assign N2049 = N2048 & pe_o_2__4_;
  assign N2050 = N2049 & N2053;
  assign N2051 = N2050 & N2054;
  assign N2052 = N2051 & pe_o_2__0_;
  assign N7654 = N2052 & N2055;
  assign N2053 = ~pe_o_2__3_;
  assign N2054 = ~pe_o_2__2_;
  assign N2055 = ~pe_o_2__1_;
  assign N2056 = pe_o_2__6_ & pe_o_2__5_;
  assign N2057 = N2056 & pe_o_2__4_;
  assign N2058 = N2057 & N2061;
  assign N2059 = N2058 & N2062;
  assign N2060 = N2059 & N2063;
  assign N7656 = N2060 & pe_o_2__1_;
  assign N2061 = ~pe_o_2__3_;
  assign N2062 = ~pe_o_2__2_;
  assign N2063 = ~pe_o_2__0_;
  assign N2064 = pe_o_2__6_ & pe_o_2__5_;
  assign N2065 = N2064 & pe_o_2__4_;
  assign N2066 = N2065 & N2069;
  assign N2067 = N2066 & N2070;
  assign N2068 = N2067 & pe_o_2__0_;
  assign N7658 = N2068 & pe_o_2__1_;
  assign N2069 = ~pe_o_2__3_;
  assign N2070 = ~pe_o_2__2_;
  assign N2071 = pe_o_2__6_ & pe_o_2__5_;
  assign N2072 = N2071 & pe_o_2__4_;
  assign N2073 = N2072 & N2076;
  assign N2074 = N2073 & pe_o_2__2_;
  assign N2075 = N2074 & N2077;
  assign N7660 = N2075 & N2078;
  assign N2076 = ~pe_o_2__3_;
  assign N2077 = ~pe_o_2__0_;
  assign N2078 = ~pe_o_2__1_;
  assign N2079 = pe_o_2__6_ & pe_o_2__5_;
  assign N2080 = N2079 & pe_o_2__4_;
  assign N2081 = N2080 & N2084;
  assign N2082 = N2081 & pe_o_2__2_;
  assign N2083 = N2082 & pe_o_2__0_;
  assign N7662 = N2083 & N2085;
  assign N2084 = ~pe_o_2__3_;
  assign N2085 = ~pe_o_2__1_;
  assign N2086 = pe_o_2__6_ & pe_o_2__5_;
  assign N2087 = N2086 & pe_o_2__4_;
  assign N2088 = N2087 & N2091;
  assign N2089 = N2088 & pe_o_2__2_;
  assign N2090 = N2089 & N2092;
  assign N7664 = N2090 & pe_o_2__1_;
  assign N2091 = ~pe_o_2__3_;
  assign N2092 = ~pe_o_2__0_;
  assign N2093 = pe_o_2__6_ & pe_o_2__5_;
  assign N2094 = N2093 & pe_o_2__4_;
  assign N2095 = N2094 & pe_o_2__2_;
  assign N2096 = N2095 & pe_o_2__0_;
  assign N7666 = N2096 & pe_o_2__1_;
  assign N2097 = pe_o_2__6_ & pe_o_2__5_;
  assign N2098 = N2097 & pe_o_2__4_;
  assign N2099 = N2098 & pe_o_2__3_;
  assign N2100 = N2099 & N2102;
  assign N2101 = N2100 & N2103;
  assign N7668 = N2101 & N2104;
  assign N2102 = ~pe_o_2__2_;
  assign N2103 = ~pe_o_2__0_;
  assign N2104 = ~pe_o_2__1_;
  assign N2105 = pe_o_2__6_ & pe_o_2__5_;
  assign N2106 = N2105 & pe_o_2__4_;
  assign N2107 = N2106 & pe_o_2__3_;
  assign N2108 = N2107 & N2110;
  assign N2109 = N2108 & pe_o_2__0_;
  assign N7670 = N2109 & N2111;
  assign N2110 = ~pe_o_2__2_;
  assign N2111 = ~pe_o_2__1_;
  assign N2112 = pe_o_2__6_ & pe_o_2__5_;
  assign N2113 = N2112 & pe_o_2__4_;
  assign N2114 = N2113 & pe_o_2__3_;
  assign N2115 = N2114 & N2117;
  assign N2116 = N2115 & N2118;
  assign N7672 = N2116 & pe_o_2__1_;
  assign N2117 = ~pe_o_2__2_;
  assign N2118 = ~pe_o_2__0_;
  assign N2119 = pe_o_2__6_ & pe_o_2__5_;
  assign N2120 = N2119 & pe_o_2__4_;
  assign N2121 = N2120 & pe_o_2__3_;
  assign N2122 = N2121 & pe_o_2__0_;
  assign N7674 = N2122 & pe_o_2__1_;
  assign N2123 = pe_o_2__6_ & pe_o_2__5_;
  assign N2124 = N2123 & pe_o_2__4_;
  assign N2125 = N2124 & pe_o_2__3_;
  assign N2126 = N2125 & pe_o_2__2_;
  assign N2127 = N2126 & N2128;
  assign N7676 = N2127 & N2129;
  assign N2128 = ~pe_o_2__0_;
  assign N2129 = ~pe_o_2__1_;
  assign N2130 = pe_o_2__6_ & pe_o_2__5_;
  assign N2131 = N2130 & pe_o_2__4_;
  assign N2132 = N2131 & pe_o_2__3_;
  assign N2133 = N2132 & pe_o_2__2_;
  assign N7678 = N2133 & pe_o_2__0_;
  assign N2134 = pe_o_2__6_ & pe_o_2__5_;
  assign N2135 = N2134 & pe_o_2__4_;
  assign N2136 = N2135 & pe_o_2__3_;
  assign N2137 = N2136 & pe_o_2__2_;
  assign N7680 = N2137 & pe_o_2__1_;
  assign N2138 = N2143 & N2144;
  assign N2139 = N2138 & N2145;
  assign N2140 = N2139 & N2146;
  assign N2141 = N2140 & N2147;
  assign N2142 = N2141 & N2148;
  assign N7809 = N2142 & N2149;
  assign N2143 = ~pe_o_3__6_;
  assign N2144 = ~pe_o_3__5_;
  assign N2145 = ~pe_o_3__4_;
  assign N2146 = ~pe_o_3__3_;
  assign N2147 = ~pe_o_3__2_;
  assign N2148 = ~pe_o_3__0_;
  assign N2149 = ~pe_o_3__1_;
  assign N2150 = pe_o_3__6_ & N2155;
  assign N2151 = N2150 & N2156;
  assign N2152 = N2151 & N2157;
  assign N2153 = N2152 & N2158;
  assign N2154 = N2153 & N2159;
  assign N7810 = N2154 & N2160;
  assign N2155 = ~pe_o_3__5_;
  assign N2156 = ~pe_o_3__4_;
  assign N2157 = ~pe_o_3__3_;
  assign N2158 = ~pe_o_3__2_;
  assign N2159 = ~pe_o_3__0_;
  assign N2160 = ~pe_o_3__1_;
  assign N2161 = N2166 & N2167;
  assign N2162 = N2161 & N2168;
  assign N2163 = N2162 & N2169;
  assign N2164 = N2163 & N2170;
  assign N2165 = N2164 & pe_o_3__0_;
  assign N7811 = N2165 & N2171;
  assign N2166 = ~pe_o_3__6_;
  assign N2167 = ~pe_o_3__5_;
  assign N2168 = ~pe_o_3__4_;
  assign N2169 = ~pe_o_3__3_;
  assign N2170 = ~pe_o_3__2_;
  assign N2171 = ~pe_o_3__1_;
  assign N2172 = N2177 & N2178;
  assign N2173 = N2172 & N2179;
  assign N2174 = N2173 & N2180;
  assign N2175 = N2174 & N2181;
  assign N2176 = N2175 & N2182;
  assign N7813 = N2176 & pe_o_3__1_;
  assign N2177 = ~pe_o_3__6_;
  assign N2178 = ~pe_o_3__5_;
  assign N2179 = ~pe_o_3__4_;
  assign N2180 = ~pe_o_3__3_;
  assign N2181 = ~pe_o_3__2_;
  assign N2182 = ~pe_o_3__0_;
  assign N2183 = N2188 & N2189;
  assign N2184 = N2183 & N2190;
  assign N2185 = N2184 & N2191;
  assign N2186 = N2185 & N2192;
  assign N2187 = N2186 & pe_o_3__0_;
  assign N7815 = N2187 & pe_o_3__1_;
  assign N2188 = ~pe_o_3__6_;
  assign N2189 = ~pe_o_3__5_;
  assign N2190 = ~pe_o_3__4_;
  assign N2191 = ~pe_o_3__3_;
  assign N2192 = ~pe_o_3__2_;
  assign N2193 = N2198 & N2199;
  assign N2194 = N2193 & N2200;
  assign N2195 = N2194 & N2201;
  assign N2196 = N2195 & pe_o_3__2_;
  assign N2197 = N2196 & N2202;
  assign N7817 = N2197 & N2203;
  assign N2198 = ~pe_o_3__6_;
  assign N2199 = ~pe_o_3__5_;
  assign N2200 = ~pe_o_3__4_;
  assign N2201 = ~pe_o_3__3_;
  assign N2202 = ~pe_o_3__0_;
  assign N2203 = ~pe_o_3__1_;
  assign N2204 = N2209 & N2210;
  assign N2205 = N2204 & N2211;
  assign N2206 = N2205 & N2212;
  assign N2207 = N2206 & pe_o_3__2_;
  assign N2208 = N2207 & pe_o_3__0_;
  assign N7819 = N2208 & N2213;
  assign N2209 = ~pe_o_3__6_;
  assign N2210 = ~pe_o_3__5_;
  assign N2211 = ~pe_o_3__4_;
  assign N2212 = ~pe_o_3__3_;
  assign N2213 = ~pe_o_3__1_;
  assign N2214 = N2219 & N2220;
  assign N2215 = N2214 & N2221;
  assign N2216 = N2215 & N2222;
  assign N2217 = N2216 & pe_o_3__2_;
  assign N2218 = N2217 & N2223;
  assign N7821 = N2218 & pe_o_3__1_;
  assign N2219 = ~pe_o_3__6_;
  assign N2220 = ~pe_o_3__5_;
  assign N2221 = ~pe_o_3__4_;
  assign N2222 = ~pe_o_3__3_;
  assign N2223 = ~pe_o_3__0_;
  assign N2224 = N2229 & N2230;
  assign N2225 = N2224 & N2231;
  assign N2226 = N2225 & N2232;
  assign N2227 = N2226 & pe_o_3__2_;
  assign N2228 = N2227 & pe_o_3__0_;
  assign N7823 = N2228 & pe_o_3__1_;
  assign N2229 = ~pe_o_3__6_;
  assign N2230 = ~pe_o_3__5_;
  assign N2231 = ~pe_o_3__4_;
  assign N2232 = ~pe_o_3__3_;
  assign N2233 = N2238 & N2239;
  assign N2234 = N2233 & N2240;
  assign N2235 = N2234 & pe_o_3__3_;
  assign N2236 = N2235 & N2241;
  assign N2237 = N2236 & N2242;
  assign N7825 = N2237 & N2243;
  assign N2238 = ~pe_o_3__6_;
  assign N2239 = ~pe_o_3__5_;
  assign N2240 = ~pe_o_3__4_;
  assign N2241 = ~pe_o_3__2_;
  assign N2242 = ~pe_o_3__0_;
  assign N2243 = ~pe_o_3__1_;
  assign N2244 = N2249 & N2250;
  assign N2245 = N2244 & N2251;
  assign N2246 = N2245 & pe_o_3__3_;
  assign N2247 = N2246 & N2252;
  assign N2248 = N2247 & pe_o_3__0_;
  assign N7827 = N2248 & N2253;
  assign N2249 = ~pe_o_3__6_;
  assign N2250 = ~pe_o_3__5_;
  assign N2251 = ~pe_o_3__4_;
  assign N2252 = ~pe_o_3__2_;
  assign N2253 = ~pe_o_3__1_;
  assign N2254 = N2259 & N2260;
  assign N2255 = N2254 & N2261;
  assign N2256 = N2255 & pe_o_3__3_;
  assign N2257 = N2256 & N2262;
  assign N2258 = N2257 & N2263;
  assign N7829 = N2258 & pe_o_3__1_;
  assign N2259 = ~pe_o_3__6_;
  assign N2260 = ~pe_o_3__5_;
  assign N2261 = ~pe_o_3__4_;
  assign N2262 = ~pe_o_3__2_;
  assign N2263 = ~pe_o_3__0_;
  assign N2264 = N2269 & N2270;
  assign N2265 = N2264 & N2271;
  assign N2266 = N2265 & pe_o_3__3_;
  assign N2267 = N2266 & N2272;
  assign N2268 = N2267 & pe_o_3__0_;
  assign N7831 = N2268 & pe_o_3__1_;
  assign N2269 = ~pe_o_3__6_;
  assign N2270 = ~pe_o_3__5_;
  assign N2271 = ~pe_o_3__4_;
  assign N2272 = ~pe_o_3__2_;
  assign N2273 = N2278 & N2279;
  assign N2274 = N2273 & N2280;
  assign N2275 = N2274 & pe_o_3__3_;
  assign N2276 = N2275 & pe_o_3__2_;
  assign N2277 = N2276 & N2281;
  assign N7833 = N2277 & N2282;
  assign N2278 = ~pe_o_3__6_;
  assign N2279 = ~pe_o_3__5_;
  assign N2280 = ~pe_o_3__4_;
  assign N2281 = ~pe_o_3__0_;
  assign N2282 = ~pe_o_3__1_;
  assign N2283 = N2288 & N2289;
  assign N2284 = N2283 & N2290;
  assign N2285 = N2284 & pe_o_3__3_;
  assign N2286 = N2285 & pe_o_3__2_;
  assign N2287 = N2286 & pe_o_3__0_;
  assign N7835 = N2287 & N2291;
  assign N2288 = ~pe_o_3__6_;
  assign N2289 = ~pe_o_3__5_;
  assign N2290 = ~pe_o_3__4_;
  assign N2291 = ~pe_o_3__1_;
  assign N2292 = N2297 & N2298;
  assign N2293 = N2292 & N2299;
  assign N2294 = N2293 & pe_o_3__3_;
  assign N2295 = N2294 & pe_o_3__2_;
  assign N2296 = N2295 & N2300;
  assign N7837 = N2296 & pe_o_3__1_;
  assign N2297 = ~pe_o_3__6_;
  assign N2298 = ~pe_o_3__5_;
  assign N2299 = ~pe_o_3__4_;
  assign N2300 = ~pe_o_3__0_;
  assign N2301 = N2306 & N2307;
  assign N2302 = N2301 & N2308;
  assign N2303 = N2302 & pe_o_3__3_;
  assign N2304 = N2303 & pe_o_3__2_;
  assign N2305 = N2304 & pe_o_3__0_;
  assign N7839 = N2305 & pe_o_3__1_;
  assign N2306 = ~pe_o_3__6_;
  assign N2307 = ~pe_o_3__5_;
  assign N2308 = ~pe_o_3__4_;
  assign N2309 = N2314 & N2315;
  assign N2310 = N2309 & pe_o_3__4_;
  assign N2311 = N2310 & N2316;
  assign N2312 = N2311 & N2317;
  assign N2313 = N2312 & N2318;
  assign N7841 = N2313 & N2319;
  assign N2314 = ~pe_o_3__6_;
  assign N2315 = ~pe_o_3__5_;
  assign N2316 = ~pe_o_3__3_;
  assign N2317 = ~pe_o_3__2_;
  assign N2318 = ~pe_o_3__0_;
  assign N2319 = ~pe_o_3__1_;
  assign N2320 = N2325 & N2326;
  assign N2321 = N2320 & pe_o_3__4_;
  assign N2322 = N2321 & N2327;
  assign N2323 = N2322 & N2328;
  assign N2324 = N2323 & pe_o_3__0_;
  assign N7843 = N2324 & N2329;
  assign N2325 = ~pe_o_3__6_;
  assign N2326 = ~pe_o_3__5_;
  assign N2327 = ~pe_o_3__3_;
  assign N2328 = ~pe_o_3__2_;
  assign N2329 = ~pe_o_3__1_;
  assign N2330 = N2335 & N2336;
  assign N2331 = N2330 & pe_o_3__4_;
  assign N2332 = N2331 & N2337;
  assign N2333 = N2332 & N2338;
  assign N2334 = N2333 & N2339;
  assign N7845 = N2334 & pe_o_3__1_;
  assign N2335 = ~pe_o_3__6_;
  assign N2336 = ~pe_o_3__5_;
  assign N2337 = ~pe_o_3__3_;
  assign N2338 = ~pe_o_3__2_;
  assign N2339 = ~pe_o_3__0_;
  assign N2340 = N2345 & N2346;
  assign N2341 = N2340 & pe_o_3__4_;
  assign N2342 = N2341 & N2347;
  assign N2343 = N2342 & N2348;
  assign N2344 = N2343 & pe_o_3__0_;
  assign N7847 = N2344 & pe_o_3__1_;
  assign N2345 = ~pe_o_3__6_;
  assign N2346 = ~pe_o_3__5_;
  assign N2347 = ~pe_o_3__3_;
  assign N2348 = ~pe_o_3__2_;
  assign N2349 = N2354 & N2355;
  assign N2350 = N2349 & pe_o_3__4_;
  assign N2351 = N2350 & N2356;
  assign N2352 = N2351 & pe_o_3__2_;
  assign N2353 = N2352 & N2357;
  assign N7849 = N2353 & N2358;
  assign N2354 = ~pe_o_3__6_;
  assign N2355 = ~pe_o_3__5_;
  assign N2356 = ~pe_o_3__3_;
  assign N2357 = ~pe_o_3__0_;
  assign N2358 = ~pe_o_3__1_;
  assign N2359 = N2364 & N2365;
  assign N2360 = N2359 & pe_o_3__4_;
  assign N2361 = N2360 & N2366;
  assign N2362 = N2361 & pe_o_3__2_;
  assign N2363 = N2362 & pe_o_3__0_;
  assign N7851 = N2363 & N2367;
  assign N2364 = ~pe_o_3__6_;
  assign N2365 = ~pe_o_3__5_;
  assign N2366 = ~pe_o_3__3_;
  assign N2367 = ~pe_o_3__1_;
  assign N2368 = N2373 & N2374;
  assign N2369 = N2368 & pe_o_3__4_;
  assign N2370 = N2369 & N2375;
  assign N2371 = N2370 & pe_o_3__2_;
  assign N2372 = N2371 & N2376;
  assign N7853 = N2372 & pe_o_3__1_;
  assign N2373 = ~pe_o_3__6_;
  assign N2374 = ~pe_o_3__5_;
  assign N2375 = ~pe_o_3__3_;
  assign N2376 = ~pe_o_3__0_;
  assign N2377 = N2382 & N2383;
  assign N2378 = N2377 & pe_o_3__4_;
  assign N2379 = N2378 & N2384;
  assign N2380 = N2379 & pe_o_3__2_;
  assign N2381 = N2380 & pe_o_3__0_;
  assign N7855 = N2381 & pe_o_3__1_;
  assign N2382 = ~pe_o_3__6_;
  assign N2383 = ~pe_o_3__5_;
  assign N2384 = ~pe_o_3__3_;
  assign N2385 = N2390 & N2391;
  assign N2386 = N2385 & pe_o_3__4_;
  assign N2387 = N2386 & pe_o_3__3_;
  assign N2388 = N2387 & N2392;
  assign N2389 = N2388 & N2393;
  assign N7857 = N2389 & N2394;
  assign N2390 = ~pe_o_3__6_;
  assign N2391 = ~pe_o_3__5_;
  assign N2392 = ~pe_o_3__2_;
  assign N2393 = ~pe_o_3__0_;
  assign N2394 = ~pe_o_3__1_;
  assign N2395 = N2400 & N2401;
  assign N2396 = N2395 & pe_o_3__4_;
  assign N2397 = N2396 & pe_o_3__3_;
  assign N2398 = N2397 & N2402;
  assign N2399 = N2398 & pe_o_3__0_;
  assign N7859 = N2399 & N2403;
  assign N2400 = ~pe_o_3__6_;
  assign N2401 = ~pe_o_3__5_;
  assign N2402 = ~pe_o_3__2_;
  assign N2403 = ~pe_o_3__1_;
  assign N2404 = N2409 & N2410;
  assign N2405 = N2404 & pe_o_3__4_;
  assign N2406 = N2405 & pe_o_3__3_;
  assign N2407 = N2406 & N2411;
  assign N2408 = N2407 & N2412;
  assign N7861 = N2408 & pe_o_3__1_;
  assign N2409 = ~pe_o_3__6_;
  assign N2410 = ~pe_o_3__5_;
  assign N2411 = ~pe_o_3__2_;
  assign N2412 = ~pe_o_3__0_;
  assign N2413 = N2418 & N2419;
  assign N2414 = N2413 & pe_o_3__4_;
  assign N2415 = N2414 & pe_o_3__3_;
  assign N2416 = N2415 & N2420;
  assign N2417 = N2416 & pe_o_3__0_;
  assign N7863 = N2417 & pe_o_3__1_;
  assign N2418 = ~pe_o_3__6_;
  assign N2419 = ~pe_o_3__5_;
  assign N2420 = ~pe_o_3__2_;
  assign N2421 = N2426 & N2427;
  assign N2422 = N2421 & pe_o_3__4_;
  assign N2423 = N2422 & pe_o_3__3_;
  assign N2424 = N2423 & pe_o_3__2_;
  assign N2425 = N2424 & N2428;
  assign N7865 = N2425 & N2429;
  assign N2426 = ~pe_o_3__6_;
  assign N2427 = ~pe_o_3__5_;
  assign N2428 = ~pe_o_3__0_;
  assign N2429 = ~pe_o_3__1_;
  assign N2430 = N2435 & N2436;
  assign N2431 = N2430 & pe_o_3__4_;
  assign N2432 = N2431 & pe_o_3__3_;
  assign N2433 = N2432 & pe_o_3__2_;
  assign N2434 = N2433 & pe_o_3__0_;
  assign N7867 = N2434 & N2437;
  assign N2435 = ~pe_o_3__6_;
  assign N2436 = ~pe_o_3__5_;
  assign N2437 = ~pe_o_3__1_;
  assign N2438 = N2443 & N2444;
  assign N2439 = N2438 & pe_o_3__4_;
  assign N2440 = N2439 & pe_o_3__3_;
  assign N2441 = N2440 & pe_o_3__2_;
  assign N2442 = N2441 & N2445;
  assign N7869 = N2442 & pe_o_3__1_;
  assign N2443 = ~pe_o_3__6_;
  assign N2444 = ~pe_o_3__5_;
  assign N2445 = ~pe_o_3__0_;
  assign N2446 = N2451 & N2452;
  assign N2447 = N2446 & pe_o_3__4_;
  assign N2448 = N2447 & pe_o_3__3_;
  assign N2449 = N2448 & pe_o_3__2_;
  assign N2450 = N2449 & pe_o_3__0_;
  assign N7871 = N2450 & pe_o_3__1_;
  assign N2451 = ~pe_o_3__6_;
  assign N2452 = ~pe_o_3__5_;
  assign N2453 = N2458 & pe_o_3__5_;
  assign N2454 = N2453 & N2459;
  assign N2455 = N2454 & N2460;
  assign N2456 = N2455 & N2461;
  assign N2457 = N2456 & N2462;
  assign N7873 = N2457 & N2463;
  assign N2458 = ~pe_o_3__6_;
  assign N2459 = ~pe_o_3__4_;
  assign N2460 = ~pe_o_3__3_;
  assign N2461 = ~pe_o_3__2_;
  assign N2462 = ~pe_o_3__0_;
  assign N2463 = ~pe_o_3__1_;
  assign N2464 = N2469 & pe_o_3__5_;
  assign N2465 = N2464 & N2470;
  assign N2466 = N2465 & N2471;
  assign N2467 = N2466 & N2472;
  assign N2468 = N2467 & pe_o_3__0_;
  assign N7875 = N2468 & N2473;
  assign N2469 = ~pe_o_3__6_;
  assign N2470 = ~pe_o_3__4_;
  assign N2471 = ~pe_o_3__3_;
  assign N2472 = ~pe_o_3__2_;
  assign N2473 = ~pe_o_3__1_;
  assign N2474 = N2479 & pe_o_3__5_;
  assign N2475 = N2474 & N2480;
  assign N2476 = N2475 & N2481;
  assign N2477 = N2476 & N2482;
  assign N2478 = N2477 & N2483;
  assign N7877 = N2478 & pe_o_3__1_;
  assign N2479 = ~pe_o_3__6_;
  assign N2480 = ~pe_o_3__4_;
  assign N2481 = ~pe_o_3__3_;
  assign N2482 = ~pe_o_3__2_;
  assign N2483 = ~pe_o_3__0_;
  assign N2484 = N2489 & pe_o_3__5_;
  assign N2485 = N2484 & N2490;
  assign N2486 = N2485 & N2491;
  assign N2487 = N2486 & N2492;
  assign N2488 = N2487 & pe_o_3__0_;
  assign N7879 = N2488 & pe_o_3__1_;
  assign N2489 = ~pe_o_3__6_;
  assign N2490 = ~pe_o_3__4_;
  assign N2491 = ~pe_o_3__3_;
  assign N2492 = ~pe_o_3__2_;
  assign N2493 = N2498 & pe_o_3__5_;
  assign N2494 = N2493 & N2499;
  assign N2495 = N2494 & N2500;
  assign N2496 = N2495 & pe_o_3__2_;
  assign N2497 = N2496 & N2501;
  assign N7881 = N2497 & N2502;
  assign N2498 = ~pe_o_3__6_;
  assign N2499 = ~pe_o_3__4_;
  assign N2500 = ~pe_o_3__3_;
  assign N2501 = ~pe_o_3__0_;
  assign N2502 = ~pe_o_3__1_;
  assign N2503 = N2508 & pe_o_3__5_;
  assign N2504 = N2503 & N2509;
  assign N2505 = N2504 & N2510;
  assign N2506 = N2505 & pe_o_3__2_;
  assign N2507 = N2506 & pe_o_3__0_;
  assign N7883 = N2507 & N2511;
  assign N2508 = ~pe_o_3__6_;
  assign N2509 = ~pe_o_3__4_;
  assign N2510 = ~pe_o_3__3_;
  assign N2511 = ~pe_o_3__1_;
  assign N2512 = N2517 & pe_o_3__5_;
  assign N2513 = N2512 & N2518;
  assign N2514 = N2513 & N2519;
  assign N2515 = N2514 & pe_o_3__2_;
  assign N2516 = N2515 & N2520;
  assign N7885 = N2516 & pe_o_3__1_;
  assign N2517 = ~pe_o_3__6_;
  assign N2518 = ~pe_o_3__4_;
  assign N2519 = ~pe_o_3__3_;
  assign N2520 = ~pe_o_3__0_;
  assign N2521 = N2526 & pe_o_3__5_;
  assign N2522 = N2521 & N2527;
  assign N2523 = N2522 & N2528;
  assign N2524 = N2523 & pe_o_3__2_;
  assign N2525 = N2524 & pe_o_3__0_;
  assign N7887 = N2525 & pe_o_3__1_;
  assign N2526 = ~pe_o_3__6_;
  assign N2527 = ~pe_o_3__4_;
  assign N2528 = ~pe_o_3__3_;
  assign N2529 = N2534 & pe_o_3__5_;
  assign N2530 = N2529 & N2535;
  assign N2531 = N2530 & pe_o_3__3_;
  assign N2532 = N2531 & N2536;
  assign N2533 = N2532 & N2537;
  assign N7889 = N2533 & N2538;
  assign N2534 = ~pe_o_3__6_;
  assign N2535 = ~pe_o_3__4_;
  assign N2536 = ~pe_o_3__2_;
  assign N2537 = ~pe_o_3__0_;
  assign N2538 = ~pe_o_3__1_;
  assign N2539 = N2544 & pe_o_3__5_;
  assign N2540 = N2539 & N2545;
  assign N2541 = N2540 & pe_o_3__3_;
  assign N2542 = N2541 & N2546;
  assign N2543 = N2542 & pe_o_3__0_;
  assign N7891 = N2543 & N2547;
  assign N2544 = ~pe_o_3__6_;
  assign N2545 = ~pe_o_3__4_;
  assign N2546 = ~pe_o_3__2_;
  assign N2547 = ~pe_o_3__1_;
  assign N2548 = N2553 & pe_o_3__5_;
  assign N2549 = N2548 & N2554;
  assign N2550 = N2549 & pe_o_3__3_;
  assign N2551 = N2550 & N2555;
  assign N2552 = N2551 & N2556;
  assign N7893 = N2552 & pe_o_3__1_;
  assign N2553 = ~pe_o_3__6_;
  assign N2554 = ~pe_o_3__4_;
  assign N2555 = ~pe_o_3__2_;
  assign N2556 = ~pe_o_3__0_;
  assign N2557 = N2562 & pe_o_3__5_;
  assign N2558 = N2557 & N2563;
  assign N2559 = N2558 & pe_o_3__3_;
  assign N2560 = N2559 & N2564;
  assign N2561 = N2560 & pe_o_3__0_;
  assign N7895 = N2561 & pe_o_3__1_;
  assign N2562 = ~pe_o_3__6_;
  assign N2563 = ~pe_o_3__4_;
  assign N2564 = ~pe_o_3__2_;
  assign N2565 = N2570 & pe_o_3__5_;
  assign N2566 = N2565 & N2571;
  assign N2567 = N2566 & pe_o_3__3_;
  assign N2568 = N2567 & pe_o_3__2_;
  assign N2569 = N2568 & N2572;
  assign N7897 = N2569 & N2573;
  assign N2570 = ~pe_o_3__6_;
  assign N2571 = ~pe_o_3__4_;
  assign N2572 = ~pe_o_3__0_;
  assign N2573 = ~pe_o_3__1_;
  assign N2574 = N2579 & pe_o_3__5_;
  assign N2575 = N2574 & N2580;
  assign N2576 = N2575 & pe_o_3__3_;
  assign N2577 = N2576 & pe_o_3__2_;
  assign N2578 = N2577 & pe_o_3__0_;
  assign N7899 = N2578 & N2581;
  assign N2579 = ~pe_o_3__6_;
  assign N2580 = ~pe_o_3__4_;
  assign N2581 = ~pe_o_3__1_;
  assign N2582 = N2587 & pe_o_3__5_;
  assign N2583 = N2582 & N2588;
  assign N2584 = N2583 & pe_o_3__3_;
  assign N2585 = N2584 & pe_o_3__2_;
  assign N2586 = N2585 & N2589;
  assign N7901 = N2586 & pe_o_3__1_;
  assign N2587 = ~pe_o_3__6_;
  assign N2588 = ~pe_o_3__4_;
  assign N2589 = ~pe_o_3__0_;
  assign N2590 = N2595 & pe_o_3__5_;
  assign N2591 = N2590 & N2596;
  assign N2592 = N2591 & pe_o_3__3_;
  assign N2593 = N2592 & pe_o_3__2_;
  assign N2594 = N2593 & pe_o_3__0_;
  assign N7903 = N2594 & pe_o_3__1_;
  assign N2595 = ~pe_o_3__6_;
  assign N2596 = ~pe_o_3__4_;
  assign N2597 = N2602 & pe_o_3__5_;
  assign N2598 = N2597 & pe_o_3__4_;
  assign N2599 = N2598 & N2603;
  assign N2600 = N2599 & N2604;
  assign N2601 = N2600 & N2605;
  assign N7905 = N2601 & N2606;
  assign N2602 = ~pe_o_3__6_;
  assign N2603 = ~pe_o_3__3_;
  assign N2604 = ~pe_o_3__2_;
  assign N2605 = ~pe_o_3__0_;
  assign N2606 = ~pe_o_3__1_;
  assign N2607 = N2612 & pe_o_3__5_;
  assign N2608 = N2607 & pe_o_3__4_;
  assign N2609 = N2608 & N2613;
  assign N2610 = N2609 & N2614;
  assign N2611 = N2610 & pe_o_3__0_;
  assign N7907 = N2611 & N2615;
  assign N2612 = ~pe_o_3__6_;
  assign N2613 = ~pe_o_3__3_;
  assign N2614 = ~pe_o_3__2_;
  assign N2615 = ~pe_o_3__1_;
  assign N2616 = N2621 & pe_o_3__5_;
  assign N2617 = N2616 & pe_o_3__4_;
  assign N2618 = N2617 & N2622;
  assign N2619 = N2618 & N2623;
  assign N2620 = N2619 & N2624;
  assign N7909 = N2620 & pe_o_3__1_;
  assign N2621 = ~pe_o_3__6_;
  assign N2622 = ~pe_o_3__3_;
  assign N2623 = ~pe_o_3__2_;
  assign N2624 = ~pe_o_3__0_;
  assign N2625 = N2630 & pe_o_3__5_;
  assign N2626 = N2625 & pe_o_3__4_;
  assign N2627 = N2626 & N2631;
  assign N2628 = N2627 & N2632;
  assign N2629 = N2628 & pe_o_3__0_;
  assign N7911 = N2629 & pe_o_3__1_;
  assign N2630 = ~pe_o_3__6_;
  assign N2631 = ~pe_o_3__3_;
  assign N2632 = ~pe_o_3__2_;
  assign N2633 = N2638 & pe_o_3__5_;
  assign N2634 = N2633 & pe_o_3__4_;
  assign N2635 = N2634 & N2639;
  assign N2636 = N2635 & pe_o_3__2_;
  assign N2637 = N2636 & N2640;
  assign N7913 = N2637 & N2641;
  assign N2638 = ~pe_o_3__6_;
  assign N2639 = ~pe_o_3__3_;
  assign N2640 = ~pe_o_3__0_;
  assign N2641 = ~pe_o_3__1_;
  assign N2642 = N2647 & pe_o_3__5_;
  assign N2643 = N2642 & pe_o_3__4_;
  assign N2644 = N2643 & N2648;
  assign N2645 = N2644 & pe_o_3__2_;
  assign N2646 = N2645 & pe_o_3__0_;
  assign N7915 = N2646 & N2649;
  assign N2647 = ~pe_o_3__6_;
  assign N2648 = ~pe_o_3__3_;
  assign N2649 = ~pe_o_3__1_;
  assign N2650 = N2655 & pe_o_3__5_;
  assign N2651 = N2650 & pe_o_3__4_;
  assign N2652 = N2651 & N2656;
  assign N2653 = N2652 & pe_o_3__2_;
  assign N2654 = N2653 & N2657;
  assign N7917 = N2654 & pe_o_3__1_;
  assign N2655 = ~pe_o_3__6_;
  assign N2656 = ~pe_o_3__3_;
  assign N2657 = ~pe_o_3__0_;
  assign N2658 = N2663 & pe_o_3__5_;
  assign N2659 = N2658 & pe_o_3__4_;
  assign N2660 = N2659 & N2664;
  assign N2661 = N2660 & pe_o_3__2_;
  assign N2662 = N2661 & pe_o_3__0_;
  assign N7919 = N2662 & pe_o_3__1_;
  assign N2663 = ~pe_o_3__6_;
  assign N2664 = ~pe_o_3__3_;
  assign N2665 = N2670 & pe_o_3__5_;
  assign N2666 = N2665 & pe_o_3__4_;
  assign N2667 = N2666 & pe_o_3__3_;
  assign N2668 = N2667 & N2671;
  assign N2669 = N2668 & N2672;
  assign N7921 = N2669 & N2673;
  assign N2670 = ~pe_o_3__6_;
  assign N2671 = ~pe_o_3__2_;
  assign N2672 = ~pe_o_3__0_;
  assign N2673 = ~pe_o_3__1_;
  assign N2674 = N2679 & pe_o_3__5_;
  assign N2675 = N2674 & pe_o_3__4_;
  assign N2676 = N2675 & pe_o_3__3_;
  assign N2677 = N2676 & N2680;
  assign N2678 = N2677 & pe_o_3__0_;
  assign N7923 = N2678 & N2681;
  assign N2679 = ~pe_o_3__6_;
  assign N2680 = ~pe_o_3__2_;
  assign N2681 = ~pe_o_3__1_;
  assign N2682 = N2687 & pe_o_3__5_;
  assign N2683 = N2682 & pe_o_3__4_;
  assign N2684 = N2683 & pe_o_3__3_;
  assign N2685 = N2684 & N2688;
  assign N2686 = N2685 & N2689;
  assign N7925 = N2686 & pe_o_3__1_;
  assign N2687 = ~pe_o_3__6_;
  assign N2688 = ~pe_o_3__2_;
  assign N2689 = ~pe_o_3__0_;
  assign N2690 = N2695 & pe_o_3__5_;
  assign N2691 = N2690 & pe_o_3__4_;
  assign N2692 = N2691 & pe_o_3__3_;
  assign N2693 = N2692 & N2696;
  assign N2694 = N2693 & pe_o_3__0_;
  assign N7927 = N2694 & pe_o_3__1_;
  assign N2695 = ~pe_o_3__6_;
  assign N2696 = ~pe_o_3__2_;
  assign N2697 = N2702 & pe_o_3__5_;
  assign N2698 = N2697 & pe_o_3__4_;
  assign N2699 = N2698 & pe_o_3__3_;
  assign N2700 = N2699 & pe_o_3__2_;
  assign N2701 = N2700 & N2703;
  assign N7929 = N2701 & N2704;
  assign N2702 = ~pe_o_3__6_;
  assign N2703 = ~pe_o_3__0_;
  assign N2704 = ~pe_o_3__1_;
  assign N2705 = N2710 & pe_o_3__5_;
  assign N2706 = N2705 & pe_o_3__4_;
  assign N2707 = N2706 & pe_o_3__3_;
  assign N2708 = N2707 & pe_o_3__2_;
  assign N2709 = N2708 & pe_o_3__0_;
  assign N7931 = N2709 & N2711;
  assign N2710 = ~pe_o_3__6_;
  assign N2711 = ~pe_o_3__1_;
  assign N2712 = N2717 & pe_o_3__5_;
  assign N2713 = N2712 & pe_o_3__4_;
  assign N2714 = N2713 & pe_o_3__3_;
  assign N2715 = N2714 & pe_o_3__2_;
  assign N2716 = N2715 & N2718;
  assign N7933 = N2716 & pe_o_3__1_;
  assign N2717 = ~pe_o_3__6_;
  assign N2718 = ~pe_o_3__0_;
  assign N2719 = pe_o_3__5_ & pe_o_3__4_;
  assign N2720 = N2719 & pe_o_3__3_;
  assign N2721 = N2720 & pe_o_3__2_;
  assign N2722 = N2721 & pe_o_3__0_;
  assign N7935 = N2722 & pe_o_3__1_;
  assign N2723 = pe_o_3__6_ & N2728;
  assign N2724 = N2723 & N2729;
  assign N2725 = N2724 & N2730;
  assign N2726 = N2725 & N2731;
  assign N2727 = N2726 & pe_o_3__0_;
  assign N7812 = N2727 & N2732;
  assign N2728 = ~pe_o_3__5_;
  assign N2729 = ~pe_o_3__4_;
  assign N2730 = ~pe_o_3__3_;
  assign N2731 = ~pe_o_3__2_;
  assign N2732 = ~pe_o_3__1_;
  assign N2733 = pe_o_3__6_ & N2738;
  assign N2734 = N2733 & N2739;
  assign N2735 = N2734 & N2740;
  assign N2736 = N2735 & N2741;
  assign N2737 = N2736 & N2742;
  assign N7814 = N2737 & pe_o_3__1_;
  assign N2738 = ~pe_o_3__5_;
  assign N2739 = ~pe_o_3__4_;
  assign N2740 = ~pe_o_3__3_;
  assign N2741 = ~pe_o_3__2_;
  assign N2742 = ~pe_o_3__0_;
  assign N2743 = pe_o_3__6_ & N2748;
  assign N2744 = N2743 & N2749;
  assign N2745 = N2744 & N2750;
  assign N2746 = N2745 & N2751;
  assign N2747 = N2746 & pe_o_3__0_;
  assign N7816 = N2747 & pe_o_3__1_;
  assign N2748 = ~pe_o_3__5_;
  assign N2749 = ~pe_o_3__4_;
  assign N2750 = ~pe_o_3__3_;
  assign N2751 = ~pe_o_3__2_;
  assign N2752 = pe_o_3__6_ & N2757;
  assign N2753 = N2752 & N2758;
  assign N2754 = N2753 & N2759;
  assign N2755 = N2754 & pe_o_3__2_;
  assign N2756 = N2755 & N2760;
  assign N7818 = N2756 & N2761;
  assign N2757 = ~pe_o_3__5_;
  assign N2758 = ~pe_o_3__4_;
  assign N2759 = ~pe_o_3__3_;
  assign N2760 = ~pe_o_3__0_;
  assign N2761 = ~pe_o_3__1_;
  assign N2762 = pe_o_3__6_ & N2767;
  assign N2763 = N2762 & N2768;
  assign N2764 = N2763 & N2769;
  assign N2765 = N2764 & pe_o_3__2_;
  assign N2766 = N2765 & pe_o_3__0_;
  assign N7820 = N2766 & N2770;
  assign N2767 = ~pe_o_3__5_;
  assign N2768 = ~pe_o_3__4_;
  assign N2769 = ~pe_o_3__3_;
  assign N2770 = ~pe_o_3__1_;
  assign N2771 = pe_o_3__6_ & N2776;
  assign N2772 = N2771 & N2777;
  assign N2773 = N2772 & N2778;
  assign N2774 = N2773 & pe_o_3__2_;
  assign N2775 = N2774 & N2779;
  assign N7822 = N2775 & pe_o_3__1_;
  assign N2776 = ~pe_o_3__5_;
  assign N2777 = ~pe_o_3__4_;
  assign N2778 = ~pe_o_3__3_;
  assign N2779 = ~pe_o_3__0_;
  assign N2780 = pe_o_3__6_ & N2785;
  assign N2781 = N2780 & N2786;
  assign N2782 = N2781 & N2787;
  assign N2783 = N2782 & pe_o_3__2_;
  assign N2784 = N2783 & pe_o_3__0_;
  assign N7824 = N2784 & pe_o_3__1_;
  assign N2785 = ~pe_o_3__5_;
  assign N2786 = ~pe_o_3__4_;
  assign N2787 = ~pe_o_3__3_;
  assign N2788 = pe_o_3__6_ & N2793;
  assign N2789 = N2788 & N2794;
  assign N2790 = N2789 & pe_o_3__3_;
  assign N2791 = N2790 & N2795;
  assign N2792 = N2791 & N2796;
  assign N7826 = N2792 & N2797;
  assign N2793 = ~pe_o_3__5_;
  assign N2794 = ~pe_o_3__4_;
  assign N2795 = ~pe_o_3__2_;
  assign N2796 = ~pe_o_3__0_;
  assign N2797 = ~pe_o_3__1_;
  assign N2798 = pe_o_3__6_ & N2803;
  assign N2799 = N2798 & N2804;
  assign N2800 = N2799 & pe_o_3__3_;
  assign N2801 = N2800 & N2805;
  assign N2802 = N2801 & pe_o_3__0_;
  assign N7828 = N2802 & N2806;
  assign N2803 = ~pe_o_3__5_;
  assign N2804 = ~pe_o_3__4_;
  assign N2805 = ~pe_o_3__2_;
  assign N2806 = ~pe_o_3__1_;
  assign N2807 = pe_o_3__6_ & N2812;
  assign N2808 = N2807 & N2813;
  assign N2809 = N2808 & pe_o_3__3_;
  assign N2810 = N2809 & N2814;
  assign N2811 = N2810 & N2815;
  assign N7830 = N2811 & pe_o_3__1_;
  assign N2812 = ~pe_o_3__5_;
  assign N2813 = ~pe_o_3__4_;
  assign N2814 = ~pe_o_3__2_;
  assign N2815 = ~pe_o_3__0_;
  assign N2816 = pe_o_3__6_ & N2821;
  assign N2817 = N2816 & N2822;
  assign N2818 = N2817 & pe_o_3__3_;
  assign N2819 = N2818 & N2823;
  assign N2820 = N2819 & pe_o_3__0_;
  assign N7832 = N2820 & pe_o_3__1_;
  assign N2821 = ~pe_o_3__5_;
  assign N2822 = ~pe_o_3__4_;
  assign N2823 = ~pe_o_3__2_;
  assign N2824 = pe_o_3__6_ & N2829;
  assign N2825 = N2824 & N2830;
  assign N2826 = N2825 & pe_o_3__3_;
  assign N2827 = N2826 & pe_o_3__2_;
  assign N2828 = N2827 & N2831;
  assign N7834 = N2828 & N2832;
  assign N2829 = ~pe_o_3__5_;
  assign N2830 = ~pe_o_3__4_;
  assign N2831 = ~pe_o_3__0_;
  assign N2832 = ~pe_o_3__1_;
  assign N2833 = pe_o_3__6_ & N2838;
  assign N2834 = N2833 & N2839;
  assign N2835 = N2834 & pe_o_3__3_;
  assign N2836 = N2835 & pe_o_3__2_;
  assign N2837 = N2836 & pe_o_3__0_;
  assign N7836 = N2837 & N2840;
  assign N2838 = ~pe_o_3__5_;
  assign N2839 = ~pe_o_3__4_;
  assign N2840 = ~pe_o_3__1_;
  assign N2841 = pe_o_3__6_ & N2846;
  assign N2842 = N2841 & N2847;
  assign N2843 = N2842 & pe_o_3__3_;
  assign N2844 = N2843 & pe_o_3__2_;
  assign N2845 = N2844 & N2848;
  assign N7838 = N2845 & pe_o_3__1_;
  assign N2846 = ~pe_o_3__5_;
  assign N2847 = ~pe_o_3__4_;
  assign N2848 = ~pe_o_3__0_;
  assign N2849 = pe_o_3__6_ & N2854;
  assign N2850 = N2849 & N2855;
  assign N2851 = N2850 & pe_o_3__3_;
  assign N2852 = N2851 & pe_o_3__2_;
  assign N2853 = N2852 & pe_o_3__0_;
  assign N7840 = N2853 & pe_o_3__1_;
  assign N2854 = ~pe_o_3__5_;
  assign N2855 = ~pe_o_3__4_;
  assign N2856 = pe_o_3__6_ & N2861;
  assign N2857 = N2856 & pe_o_3__4_;
  assign N2858 = N2857 & N2862;
  assign N2859 = N2858 & N2863;
  assign N2860 = N2859 & N2864;
  assign N7842 = N2860 & N2865;
  assign N2861 = ~pe_o_3__5_;
  assign N2862 = ~pe_o_3__3_;
  assign N2863 = ~pe_o_3__2_;
  assign N2864 = ~pe_o_3__0_;
  assign N2865 = ~pe_o_3__1_;
  assign N2866 = pe_o_3__6_ & N2871;
  assign N2867 = N2866 & pe_o_3__4_;
  assign N2868 = N2867 & N2872;
  assign N2869 = N2868 & N2873;
  assign N2870 = N2869 & pe_o_3__0_;
  assign N7844 = N2870 & N2874;
  assign N2871 = ~pe_o_3__5_;
  assign N2872 = ~pe_o_3__3_;
  assign N2873 = ~pe_o_3__2_;
  assign N2874 = ~pe_o_3__1_;
  assign N2875 = pe_o_3__6_ & N2880;
  assign N2876 = N2875 & pe_o_3__4_;
  assign N2877 = N2876 & N2881;
  assign N2878 = N2877 & N2882;
  assign N2879 = N2878 & N2883;
  assign N7846 = N2879 & pe_o_3__1_;
  assign N2880 = ~pe_o_3__5_;
  assign N2881 = ~pe_o_3__3_;
  assign N2882 = ~pe_o_3__2_;
  assign N2883 = ~pe_o_3__0_;
  assign N2884 = pe_o_3__6_ & N2889;
  assign N2885 = N2884 & pe_o_3__4_;
  assign N2886 = N2885 & N2890;
  assign N2887 = N2886 & N2891;
  assign N2888 = N2887 & pe_o_3__0_;
  assign N7848 = N2888 & pe_o_3__1_;
  assign N2889 = ~pe_o_3__5_;
  assign N2890 = ~pe_o_3__3_;
  assign N2891 = ~pe_o_3__2_;
  assign N2892 = pe_o_3__6_ & N2897;
  assign N2893 = N2892 & pe_o_3__4_;
  assign N2894 = N2893 & N2898;
  assign N2895 = N2894 & pe_o_3__2_;
  assign N2896 = N2895 & N2899;
  assign N7850 = N2896 & N2900;
  assign N2897 = ~pe_o_3__5_;
  assign N2898 = ~pe_o_3__3_;
  assign N2899 = ~pe_o_3__0_;
  assign N2900 = ~pe_o_3__1_;
  assign N2901 = pe_o_3__6_ & N2906;
  assign N2902 = N2901 & pe_o_3__4_;
  assign N2903 = N2902 & N2907;
  assign N2904 = N2903 & pe_o_3__2_;
  assign N2905 = N2904 & pe_o_3__0_;
  assign N7852 = N2905 & N2908;
  assign N2906 = ~pe_o_3__5_;
  assign N2907 = ~pe_o_3__3_;
  assign N2908 = ~pe_o_3__1_;
  assign N2909 = pe_o_3__6_ & N2914;
  assign N2910 = N2909 & pe_o_3__4_;
  assign N2911 = N2910 & N2915;
  assign N2912 = N2911 & pe_o_3__2_;
  assign N2913 = N2912 & N2916;
  assign N7854 = N2913 & pe_o_3__1_;
  assign N2914 = ~pe_o_3__5_;
  assign N2915 = ~pe_o_3__3_;
  assign N2916 = ~pe_o_3__0_;
  assign N2917 = pe_o_3__6_ & N2922;
  assign N2918 = N2917 & pe_o_3__4_;
  assign N2919 = N2918 & N2923;
  assign N2920 = N2919 & pe_o_3__2_;
  assign N2921 = N2920 & pe_o_3__0_;
  assign N7856 = N2921 & pe_o_3__1_;
  assign N2922 = ~pe_o_3__5_;
  assign N2923 = ~pe_o_3__3_;
  assign N2924 = pe_o_3__6_ & N2929;
  assign N2925 = N2924 & pe_o_3__4_;
  assign N2926 = N2925 & pe_o_3__3_;
  assign N2927 = N2926 & N2930;
  assign N2928 = N2927 & N2931;
  assign N7858 = N2928 & N2932;
  assign N2929 = ~pe_o_3__5_;
  assign N2930 = ~pe_o_3__2_;
  assign N2931 = ~pe_o_3__0_;
  assign N2932 = ~pe_o_3__1_;
  assign N2933 = pe_o_3__6_ & N2938;
  assign N2934 = N2933 & pe_o_3__4_;
  assign N2935 = N2934 & pe_o_3__3_;
  assign N2936 = N2935 & N2939;
  assign N2937 = N2936 & pe_o_3__0_;
  assign N7860 = N2937 & N2940;
  assign N2938 = ~pe_o_3__5_;
  assign N2939 = ~pe_o_3__2_;
  assign N2940 = ~pe_o_3__1_;
  assign N2941 = pe_o_3__6_ & N2946;
  assign N2942 = N2941 & pe_o_3__4_;
  assign N2943 = N2942 & pe_o_3__3_;
  assign N2944 = N2943 & N2947;
  assign N2945 = N2944 & N2948;
  assign N7862 = N2945 & pe_o_3__1_;
  assign N2946 = ~pe_o_3__5_;
  assign N2947 = ~pe_o_3__2_;
  assign N2948 = ~pe_o_3__0_;
  assign N2949 = pe_o_3__6_ & N2954;
  assign N2950 = N2949 & pe_o_3__4_;
  assign N2951 = N2950 & pe_o_3__3_;
  assign N2952 = N2951 & N2955;
  assign N2953 = N2952 & pe_o_3__0_;
  assign N7864 = N2953 & pe_o_3__1_;
  assign N2954 = ~pe_o_3__5_;
  assign N2955 = ~pe_o_3__2_;
  assign N2956 = pe_o_3__6_ & N2961;
  assign N2957 = N2956 & pe_o_3__4_;
  assign N2958 = N2957 & pe_o_3__3_;
  assign N2959 = N2958 & pe_o_3__2_;
  assign N2960 = N2959 & N2962;
  assign N7866 = N2960 & N2963;
  assign N2961 = ~pe_o_3__5_;
  assign N2962 = ~pe_o_3__0_;
  assign N2963 = ~pe_o_3__1_;
  assign N2964 = pe_o_3__6_ & N2969;
  assign N2965 = N2964 & pe_o_3__4_;
  assign N2966 = N2965 & pe_o_3__3_;
  assign N2967 = N2966 & pe_o_3__2_;
  assign N2968 = N2967 & pe_o_3__0_;
  assign N7868 = N2968 & N2970;
  assign N2969 = ~pe_o_3__5_;
  assign N2970 = ~pe_o_3__1_;
  assign N2971 = pe_o_3__6_ & N2976;
  assign N2972 = N2971 & pe_o_3__4_;
  assign N2973 = N2972 & pe_o_3__3_;
  assign N2974 = N2973 & pe_o_3__2_;
  assign N2975 = N2974 & N2977;
  assign N7870 = N2975 & pe_o_3__1_;
  assign N2976 = ~pe_o_3__5_;
  assign N2977 = ~pe_o_3__0_;
  assign N2978 = pe_o_3__6_ & pe_o_3__4_;
  assign N2979 = N2978 & pe_o_3__3_;
  assign N2980 = N2979 & pe_o_3__2_;
  assign N2981 = N2980 & pe_o_3__0_;
  assign N7872 = N2981 & pe_o_3__1_;
  assign N2982 = pe_o_3__6_ & pe_o_3__5_;
  assign N2983 = N2982 & N2987;
  assign N2984 = N2983 & N2988;
  assign N2985 = N2984 & N2989;
  assign N2986 = N2985 & N2990;
  assign N7874 = N2986 & N2991;
  assign N2987 = ~pe_o_3__4_;
  assign N2988 = ~pe_o_3__3_;
  assign N2989 = ~pe_o_3__2_;
  assign N2990 = ~pe_o_3__0_;
  assign N2991 = ~pe_o_3__1_;
  assign N2992 = pe_o_3__6_ & pe_o_3__5_;
  assign N2993 = N2992 & N2997;
  assign N2994 = N2993 & N2998;
  assign N2995 = N2994 & N2999;
  assign N2996 = N2995 & pe_o_3__0_;
  assign N7876 = N2996 & N3000;
  assign N2997 = ~pe_o_3__4_;
  assign N2998 = ~pe_o_3__3_;
  assign N2999 = ~pe_o_3__2_;
  assign N3000 = ~pe_o_3__1_;
  assign N3001 = pe_o_3__6_ & pe_o_3__5_;
  assign N3002 = N3001 & N3006;
  assign N3003 = N3002 & N3007;
  assign N3004 = N3003 & N3008;
  assign N3005 = N3004 & N3009;
  assign N7878 = N3005 & pe_o_3__1_;
  assign N3006 = ~pe_o_3__4_;
  assign N3007 = ~pe_o_3__3_;
  assign N3008 = ~pe_o_3__2_;
  assign N3009 = ~pe_o_3__0_;
  assign N3010 = pe_o_3__6_ & pe_o_3__5_;
  assign N3011 = N3010 & N3015;
  assign N3012 = N3011 & N3016;
  assign N3013 = N3012 & N3017;
  assign N3014 = N3013 & pe_o_3__0_;
  assign N7880 = N3014 & pe_o_3__1_;
  assign N3015 = ~pe_o_3__4_;
  assign N3016 = ~pe_o_3__3_;
  assign N3017 = ~pe_o_3__2_;
  assign N3018 = pe_o_3__6_ & pe_o_3__5_;
  assign N3019 = N3018 & N3023;
  assign N3020 = N3019 & N3024;
  assign N3021 = N3020 & pe_o_3__2_;
  assign N3022 = N3021 & N3025;
  assign N7882 = N3022 & N3026;
  assign N3023 = ~pe_o_3__4_;
  assign N3024 = ~pe_o_3__3_;
  assign N3025 = ~pe_o_3__0_;
  assign N3026 = ~pe_o_3__1_;
  assign N3027 = pe_o_3__6_ & pe_o_3__5_;
  assign N3028 = N3027 & N3032;
  assign N3029 = N3028 & N3033;
  assign N3030 = N3029 & pe_o_3__2_;
  assign N3031 = N3030 & pe_o_3__0_;
  assign N7884 = N3031 & N3034;
  assign N3032 = ~pe_o_3__4_;
  assign N3033 = ~pe_o_3__3_;
  assign N3034 = ~pe_o_3__1_;
  assign N3035 = pe_o_3__6_ & pe_o_3__5_;
  assign N3036 = N3035 & N3040;
  assign N3037 = N3036 & N3041;
  assign N3038 = N3037 & pe_o_3__2_;
  assign N3039 = N3038 & N3042;
  assign N7886 = N3039 & pe_o_3__1_;
  assign N3040 = ~pe_o_3__4_;
  assign N3041 = ~pe_o_3__3_;
  assign N3042 = ~pe_o_3__0_;
  assign N3043 = pe_o_3__6_ & pe_o_3__5_;
  assign N3044 = N3043 & N3048;
  assign N3045 = N3044 & N3049;
  assign N3046 = N3045 & pe_o_3__2_;
  assign N3047 = N3046 & pe_o_3__0_;
  assign N7888 = N3047 & pe_o_3__1_;
  assign N3048 = ~pe_o_3__4_;
  assign N3049 = ~pe_o_3__3_;
  assign N3050 = pe_o_3__6_ & pe_o_3__5_;
  assign N3051 = N3050 & N3055;
  assign N3052 = N3051 & pe_o_3__3_;
  assign N3053 = N3052 & N3056;
  assign N3054 = N3053 & N3057;
  assign N7890 = N3054 & N3058;
  assign N3055 = ~pe_o_3__4_;
  assign N3056 = ~pe_o_3__2_;
  assign N3057 = ~pe_o_3__0_;
  assign N3058 = ~pe_o_3__1_;
  assign N3059 = pe_o_3__6_ & pe_o_3__5_;
  assign N3060 = N3059 & N3064;
  assign N3061 = N3060 & pe_o_3__3_;
  assign N3062 = N3061 & N3065;
  assign N3063 = N3062 & pe_o_3__0_;
  assign N7892 = N3063 & N3066;
  assign N3064 = ~pe_o_3__4_;
  assign N3065 = ~pe_o_3__2_;
  assign N3066 = ~pe_o_3__1_;
  assign N3067 = pe_o_3__6_ & pe_o_3__5_;
  assign N3068 = N3067 & N3072;
  assign N3069 = N3068 & pe_o_3__3_;
  assign N3070 = N3069 & N3073;
  assign N3071 = N3070 & N3074;
  assign N7894 = N3071 & pe_o_3__1_;
  assign N3072 = ~pe_o_3__4_;
  assign N3073 = ~pe_o_3__2_;
  assign N3074 = ~pe_o_3__0_;
  assign N3075 = pe_o_3__6_ & pe_o_3__5_;
  assign N3076 = N3075 & N3080;
  assign N3077 = N3076 & pe_o_3__3_;
  assign N3078 = N3077 & N3081;
  assign N3079 = N3078 & pe_o_3__0_;
  assign N7896 = N3079 & pe_o_3__1_;
  assign N3080 = ~pe_o_3__4_;
  assign N3081 = ~pe_o_3__2_;
  assign N3082 = pe_o_3__6_ & pe_o_3__5_;
  assign N3083 = N3082 & N3087;
  assign N3084 = N3083 & pe_o_3__3_;
  assign N3085 = N3084 & pe_o_3__2_;
  assign N3086 = N3085 & N3088;
  assign N7898 = N3086 & N3089;
  assign N3087 = ~pe_o_3__4_;
  assign N3088 = ~pe_o_3__0_;
  assign N3089 = ~pe_o_3__1_;
  assign N3090 = pe_o_3__6_ & pe_o_3__5_;
  assign N3091 = N3090 & N3095;
  assign N3092 = N3091 & pe_o_3__3_;
  assign N3093 = N3092 & pe_o_3__2_;
  assign N3094 = N3093 & pe_o_3__0_;
  assign N7900 = N3094 & N3096;
  assign N3095 = ~pe_o_3__4_;
  assign N3096 = ~pe_o_3__1_;
  assign N3097 = pe_o_3__6_ & pe_o_3__5_;
  assign N3098 = N3097 & N3102;
  assign N3099 = N3098 & pe_o_3__3_;
  assign N3100 = N3099 & pe_o_3__2_;
  assign N3101 = N3100 & N3103;
  assign N7902 = N3101 & pe_o_3__1_;
  assign N3102 = ~pe_o_3__4_;
  assign N3103 = ~pe_o_3__0_;
  assign N3104 = pe_o_3__6_ & pe_o_3__5_;
  assign N3105 = N3104 & pe_o_3__3_;
  assign N3106 = N3105 & pe_o_3__2_;
  assign N3107 = N3106 & pe_o_3__0_;
  assign N7904 = N3107 & pe_o_3__1_;
  assign N3108 = pe_o_3__6_ & pe_o_3__5_;
  assign N3109 = N3108 & pe_o_3__4_;
  assign N3110 = N3109 & N3113;
  assign N3111 = N3110 & N3114;
  assign N3112 = N3111 & N3115;
  assign N7906 = N3112 & N3116;
  assign N3113 = ~pe_o_3__3_;
  assign N3114 = ~pe_o_3__2_;
  assign N3115 = ~pe_o_3__0_;
  assign N3116 = ~pe_o_3__1_;
  assign N3117 = pe_o_3__6_ & pe_o_3__5_;
  assign N3118 = N3117 & pe_o_3__4_;
  assign N3119 = N3118 & N3122;
  assign N3120 = N3119 & N3123;
  assign N3121 = N3120 & pe_o_3__0_;
  assign N7908 = N3121 & N3124;
  assign N3122 = ~pe_o_3__3_;
  assign N3123 = ~pe_o_3__2_;
  assign N3124 = ~pe_o_3__1_;
  assign N3125 = pe_o_3__6_ & pe_o_3__5_;
  assign N3126 = N3125 & pe_o_3__4_;
  assign N3127 = N3126 & N3130;
  assign N3128 = N3127 & N3131;
  assign N3129 = N3128 & N3132;
  assign N7910 = N3129 & pe_o_3__1_;
  assign N3130 = ~pe_o_3__3_;
  assign N3131 = ~pe_o_3__2_;
  assign N3132 = ~pe_o_3__0_;
  assign N3133 = pe_o_3__6_ & pe_o_3__5_;
  assign N3134 = N3133 & pe_o_3__4_;
  assign N3135 = N3134 & N3138;
  assign N3136 = N3135 & N3139;
  assign N3137 = N3136 & pe_o_3__0_;
  assign N7912 = N3137 & pe_o_3__1_;
  assign N3138 = ~pe_o_3__3_;
  assign N3139 = ~pe_o_3__2_;
  assign N3140 = pe_o_3__6_ & pe_o_3__5_;
  assign N3141 = N3140 & pe_o_3__4_;
  assign N3142 = N3141 & N3145;
  assign N3143 = N3142 & pe_o_3__2_;
  assign N3144 = N3143 & N3146;
  assign N7914 = N3144 & N3147;
  assign N3145 = ~pe_o_3__3_;
  assign N3146 = ~pe_o_3__0_;
  assign N3147 = ~pe_o_3__1_;
  assign N3148 = pe_o_3__6_ & pe_o_3__5_;
  assign N3149 = N3148 & pe_o_3__4_;
  assign N3150 = N3149 & N3153;
  assign N3151 = N3150 & pe_o_3__2_;
  assign N3152 = N3151 & pe_o_3__0_;
  assign N7916 = N3152 & N3154;
  assign N3153 = ~pe_o_3__3_;
  assign N3154 = ~pe_o_3__1_;
  assign N3155 = pe_o_3__6_ & pe_o_3__5_;
  assign N3156 = N3155 & pe_o_3__4_;
  assign N3157 = N3156 & N3160;
  assign N3158 = N3157 & pe_o_3__2_;
  assign N3159 = N3158 & N3161;
  assign N7918 = N3159 & pe_o_3__1_;
  assign N3160 = ~pe_o_3__3_;
  assign N3161 = ~pe_o_3__0_;
  assign N3162 = pe_o_3__6_ & pe_o_3__5_;
  assign N3163 = N3162 & pe_o_3__4_;
  assign N3164 = N3163 & pe_o_3__2_;
  assign N3165 = N3164 & pe_o_3__0_;
  assign N7920 = N3165 & pe_o_3__1_;
  assign N3166 = pe_o_3__6_ & pe_o_3__5_;
  assign N3167 = N3166 & pe_o_3__4_;
  assign N3168 = N3167 & pe_o_3__3_;
  assign N3169 = N3168 & N3171;
  assign N3170 = N3169 & N3172;
  assign N7922 = N3170 & N3173;
  assign N3171 = ~pe_o_3__2_;
  assign N3172 = ~pe_o_3__0_;
  assign N3173 = ~pe_o_3__1_;
  assign N3174 = pe_o_3__6_ & pe_o_3__5_;
  assign N3175 = N3174 & pe_o_3__4_;
  assign N3176 = N3175 & pe_o_3__3_;
  assign N3177 = N3176 & N3179;
  assign N3178 = N3177 & pe_o_3__0_;
  assign N7924 = N3178 & N3180;
  assign N3179 = ~pe_o_3__2_;
  assign N3180 = ~pe_o_3__1_;
  assign N3181 = pe_o_3__6_ & pe_o_3__5_;
  assign N3182 = N3181 & pe_o_3__4_;
  assign N3183 = N3182 & pe_o_3__3_;
  assign N3184 = N3183 & N3186;
  assign N3185 = N3184 & N3187;
  assign N7926 = N3185 & pe_o_3__1_;
  assign N3186 = ~pe_o_3__2_;
  assign N3187 = ~pe_o_3__0_;
  assign N3188 = pe_o_3__6_ & pe_o_3__5_;
  assign N3189 = N3188 & pe_o_3__4_;
  assign N3190 = N3189 & pe_o_3__3_;
  assign N3191 = N3190 & pe_o_3__0_;
  assign N7928 = N3191 & pe_o_3__1_;
  assign N3192 = pe_o_3__6_ & pe_o_3__5_;
  assign N3193 = N3192 & pe_o_3__4_;
  assign N3194 = N3193 & pe_o_3__3_;
  assign N3195 = N3194 & pe_o_3__2_;
  assign N3196 = N3195 & N3197;
  assign N7930 = N3196 & N3198;
  assign N3197 = ~pe_o_3__0_;
  assign N3198 = ~pe_o_3__1_;
  assign N3199 = pe_o_3__6_ & pe_o_3__5_;
  assign N3200 = N3199 & pe_o_3__4_;
  assign N3201 = N3200 & pe_o_3__3_;
  assign N3202 = N3201 & pe_o_3__2_;
  assign N7932 = N3202 & pe_o_3__0_;
  assign N3203 = pe_o_3__6_ & pe_o_3__5_;
  assign N3204 = N3203 & pe_o_3__4_;
  assign N3205 = N3204 & pe_o_3__3_;
  assign N3206 = N3205 & pe_o_3__2_;
  assign N7934 = N3206 & pe_o_3__1_;
  assign N3207 = N3212 & N3213;
  assign N3208 = N3207 & N3214;
  assign N3209 = N3208 & N3215;
  assign N3210 = N3209 & N3216;
  assign N3211 = N3210 & N3217;
  assign N8063 = N3211 & N3218;
  assign N3212 = ~pe_o_4__6_;
  assign N3213 = ~pe_o_4__5_;
  assign N3214 = ~pe_o_4__4_;
  assign N3215 = ~pe_o_4__3_;
  assign N3216 = ~pe_o_4__2_;
  assign N3217 = ~pe_o_4__0_;
  assign N3218 = ~pe_o_4__1_;
  assign N3219 = pe_o_4__6_ & N3224;
  assign N3220 = N3219 & N3225;
  assign N3221 = N3220 & N3226;
  assign N3222 = N3221 & N3227;
  assign N3223 = N3222 & N3228;
  assign N8064 = N3223 & N3229;
  assign N3224 = ~pe_o_4__5_;
  assign N3225 = ~pe_o_4__4_;
  assign N3226 = ~pe_o_4__3_;
  assign N3227 = ~pe_o_4__2_;
  assign N3228 = ~pe_o_4__0_;
  assign N3229 = ~pe_o_4__1_;
  assign N3230 = N3235 & N3236;
  assign N3231 = N3230 & N3237;
  assign N3232 = N3231 & N3238;
  assign N3233 = N3232 & N3239;
  assign N3234 = N3233 & pe_o_4__0_;
  assign N8065 = N3234 & N3240;
  assign N3235 = ~pe_o_4__6_;
  assign N3236 = ~pe_o_4__5_;
  assign N3237 = ~pe_o_4__4_;
  assign N3238 = ~pe_o_4__3_;
  assign N3239 = ~pe_o_4__2_;
  assign N3240 = ~pe_o_4__1_;
  assign N3241 = N3246 & N3247;
  assign N3242 = N3241 & N3248;
  assign N3243 = N3242 & N3249;
  assign N3244 = N3243 & N3250;
  assign N3245 = N3244 & N3251;
  assign N8067 = N3245 & pe_o_4__1_;
  assign N3246 = ~pe_o_4__6_;
  assign N3247 = ~pe_o_4__5_;
  assign N3248 = ~pe_o_4__4_;
  assign N3249 = ~pe_o_4__3_;
  assign N3250 = ~pe_o_4__2_;
  assign N3251 = ~pe_o_4__0_;
  assign N3252 = N3257 & N3258;
  assign N3253 = N3252 & N3259;
  assign N3254 = N3253 & N3260;
  assign N3255 = N3254 & N3261;
  assign N3256 = N3255 & pe_o_4__0_;
  assign N8069 = N3256 & pe_o_4__1_;
  assign N3257 = ~pe_o_4__6_;
  assign N3258 = ~pe_o_4__5_;
  assign N3259 = ~pe_o_4__4_;
  assign N3260 = ~pe_o_4__3_;
  assign N3261 = ~pe_o_4__2_;
  assign N3262 = N3267 & N3268;
  assign N3263 = N3262 & N3269;
  assign N3264 = N3263 & N3270;
  assign N3265 = N3264 & pe_o_4__2_;
  assign N3266 = N3265 & N3271;
  assign N8071 = N3266 & N3272;
  assign N3267 = ~pe_o_4__6_;
  assign N3268 = ~pe_o_4__5_;
  assign N3269 = ~pe_o_4__4_;
  assign N3270 = ~pe_o_4__3_;
  assign N3271 = ~pe_o_4__0_;
  assign N3272 = ~pe_o_4__1_;
  assign N3273 = N3278 & N3279;
  assign N3274 = N3273 & N3280;
  assign N3275 = N3274 & N3281;
  assign N3276 = N3275 & pe_o_4__2_;
  assign N3277 = N3276 & pe_o_4__0_;
  assign N8073 = N3277 & N3282;
  assign N3278 = ~pe_o_4__6_;
  assign N3279 = ~pe_o_4__5_;
  assign N3280 = ~pe_o_4__4_;
  assign N3281 = ~pe_o_4__3_;
  assign N3282 = ~pe_o_4__1_;
  assign N3283 = N3288 & N3289;
  assign N3284 = N3283 & N3290;
  assign N3285 = N3284 & N3291;
  assign N3286 = N3285 & pe_o_4__2_;
  assign N3287 = N3286 & N3292;
  assign N8075 = N3287 & pe_o_4__1_;
  assign N3288 = ~pe_o_4__6_;
  assign N3289 = ~pe_o_4__5_;
  assign N3290 = ~pe_o_4__4_;
  assign N3291 = ~pe_o_4__3_;
  assign N3292 = ~pe_o_4__0_;
  assign N3293 = N3298 & N3299;
  assign N3294 = N3293 & N3300;
  assign N3295 = N3294 & N3301;
  assign N3296 = N3295 & pe_o_4__2_;
  assign N3297 = N3296 & pe_o_4__0_;
  assign N8077 = N3297 & pe_o_4__1_;
  assign N3298 = ~pe_o_4__6_;
  assign N3299 = ~pe_o_4__5_;
  assign N3300 = ~pe_o_4__4_;
  assign N3301 = ~pe_o_4__3_;
  assign N3302 = N3307 & N3308;
  assign N3303 = N3302 & N3309;
  assign N3304 = N3303 & pe_o_4__3_;
  assign N3305 = N3304 & N3310;
  assign N3306 = N3305 & N3311;
  assign N8079 = N3306 & N3312;
  assign N3307 = ~pe_o_4__6_;
  assign N3308 = ~pe_o_4__5_;
  assign N3309 = ~pe_o_4__4_;
  assign N3310 = ~pe_o_4__2_;
  assign N3311 = ~pe_o_4__0_;
  assign N3312 = ~pe_o_4__1_;
  assign N3313 = N3318 & N3319;
  assign N3314 = N3313 & N3320;
  assign N3315 = N3314 & pe_o_4__3_;
  assign N3316 = N3315 & N3321;
  assign N3317 = N3316 & pe_o_4__0_;
  assign N8081 = N3317 & N3322;
  assign N3318 = ~pe_o_4__6_;
  assign N3319 = ~pe_o_4__5_;
  assign N3320 = ~pe_o_4__4_;
  assign N3321 = ~pe_o_4__2_;
  assign N3322 = ~pe_o_4__1_;
  assign N3323 = N3328 & N3329;
  assign N3324 = N3323 & N3330;
  assign N3325 = N3324 & pe_o_4__3_;
  assign N3326 = N3325 & N3331;
  assign N3327 = N3326 & N3332;
  assign N8083 = N3327 & pe_o_4__1_;
  assign N3328 = ~pe_o_4__6_;
  assign N3329 = ~pe_o_4__5_;
  assign N3330 = ~pe_o_4__4_;
  assign N3331 = ~pe_o_4__2_;
  assign N3332 = ~pe_o_4__0_;
  assign N3333 = N3338 & N3339;
  assign N3334 = N3333 & N3340;
  assign N3335 = N3334 & pe_o_4__3_;
  assign N3336 = N3335 & N3341;
  assign N3337 = N3336 & pe_o_4__0_;
  assign N8085 = N3337 & pe_o_4__1_;
  assign N3338 = ~pe_o_4__6_;
  assign N3339 = ~pe_o_4__5_;
  assign N3340 = ~pe_o_4__4_;
  assign N3341 = ~pe_o_4__2_;
  assign N3342 = N3347 & N3348;
  assign N3343 = N3342 & N3349;
  assign N3344 = N3343 & pe_o_4__3_;
  assign N3345 = N3344 & pe_o_4__2_;
  assign N3346 = N3345 & N3350;
  assign N8087 = N3346 & N3351;
  assign N3347 = ~pe_o_4__6_;
  assign N3348 = ~pe_o_4__5_;
  assign N3349 = ~pe_o_4__4_;
  assign N3350 = ~pe_o_4__0_;
  assign N3351 = ~pe_o_4__1_;
  assign N3352 = N3357 & N3358;
  assign N3353 = N3352 & N3359;
  assign N3354 = N3353 & pe_o_4__3_;
  assign N3355 = N3354 & pe_o_4__2_;
  assign N3356 = N3355 & pe_o_4__0_;
  assign N8089 = N3356 & N3360;
  assign N3357 = ~pe_o_4__6_;
  assign N3358 = ~pe_o_4__5_;
  assign N3359 = ~pe_o_4__4_;
  assign N3360 = ~pe_o_4__1_;
  assign N3361 = N3366 & N3367;
  assign N3362 = N3361 & N3368;
  assign N3363 = N3362 & pe_o_4__3_;
  assign N3364 = N3363 & pe_o_4__2_;
  assign N3365 = N3364 & N3369;
  assign N8091 = N3365 & pe_o_4__1_;
  assign N3366 = ~pe_o_4__6_;
  assign N3367 = ~pe_o_4__5_;
  assign N3368 = ~pe_o_4__4_;
  assign N3369 = ~pe_o_4__0_;
  assign N3370 = N3375 & N3376;
  assign N3371 = N3370 & N3377;
  assign N3372 = N3371 & pe_o_4__3_;
  assign N3373 = N3372 & pe_o_4__2_;
  assign N3374 = N3373 & pe_o_4__0_;
  assign N8093 = N3374 & pe_o_4__1_;
  assign N3375 = ~pe_o_4__6_;
  assign N3376 = ~pe_o_4__5_;
  assign N3377 = ~pe_o_4__4_;
  assign N3378 = N3383 & N3384;
  assign N3379 = N3378 & pe_o_4__4_;
  assign N3380 = N3379 & N3385;
  assign N3381 = N3380 & N3386;
  assign N3382 = N3381 & N3387;
  assign N8095 = N3382 & N3388;
  assign N3383 = ~pe_o_4__6_;
  assign N3384 = ~pe_o_4__5_;
  assign N3385 = ~pe_o_4__3_;
  assign N3386 = ~pe_o_4__2_;
  assign N3387 = ~pe_o_4__0_;
  assign N3388 = ~pe_o_4__1_;
  assign N3389 = N3394 & N3395;
  assign N3390 = N3389 & pe_o_4__4_;
  assign N3391 = N3390 & N3396;
  assign N3392 = N3391 & N3397;
  assign N3393 = N3392 & pe_o_4__0_;
  assign N8097 = N3393 & N3398;
  assign N3394 = ~pe_o_4__6_;
  assign N3395 = ~pe_o_4__5_;
  assign N3396 = ~pe_o_4__3_;
  assign N3397 = ~pe_o_4__2_;
  assign N3398 = ~pe_o_4__1_;
  assign N3399 = N3404 & N3405;
  assign N3400 = N3399 & pe_o_4__4_;
  assign N3401 = N3400 & N3406;
  assign N3402 = N3401 & N3407;
  assign N3403 = N3402 & N3408;
  assign N8099 = N3403 & pe_o_4__1_;
  assign N3404 = ~pe_o_4__6_;
  assign N3405 = ~pe_o_4__5_;
  assign N3406 = ~pe_o_4__3_;
  assign N3407 = ~pe_o_4__2_;
  assign N3408 = ~pe_o_4__0_;
  assign N3409 = N3414 & N3415;
  assign N3410 = N3409 & pe_o_4__4_;
  assign N3411 = N3410 & N3416;
  assign N3412 = N3411 & N3417;
  assign N3413 = N3412 & pe_o_4__0_;
  assign N8101 = N3413 & pe_o_4__1_;
  assign N3414 = ~pe_o_4__6_;
  assign N3415 = ~pe_o_4__5_;
  assign N3416 = ~pe_o_4__3_;
  assign N3417 = ~pe_o_4__2_;
  assign N3418 = N3423 & N3424;
  assign N3419 = N3418 & pe_o_4__4_;
  assign N3420 = N3419 & N3425;
  assign N3421 = N3420 & pe_o_4__2_;
  assign N3422 = N3421 & N3426;
  assign N8103 = N3422 & N3427;
  assign N3423 = ~pe_o_4__6_;
  assign N3424 = ~pe_o_4__5_;
  assign N3425 = ~pe_o_4__3_;
  assign N3426 = ~pe_o_4__0_;
  assign N3427 = ~pe_o_4__1_;
  assign N3428 = N3433 & N3434;
  assign N3429 = N3428 & pe_o_4__4_;
  assign N3430 = N3429 & N3435;
  assign N3431 = N3430 & pe_o_4__2_;
  assign N3432 = N3431 & pe_o_4__0_;
  assign N8105 = N3432 & N3436;
  assign N3433 = ~pe_o_4__6_;
  assign N3434 = ~pe_o_4__5_;
  assign N3435 = ~pe_o_4__3_;
  assign N3436 = ~pe_o_4__1_;
  assign N3437 = N3442 & N3443;
  assign N3438 = N3437 & pe_o_4__4_;
  assign N3439 = N3438 & N3444;
  assign N3440 = N3439 & pe_o_4__2_;
  assign N3441 = N3440 & N3445;
  assign N8107 = N3441 & pe_o_4__1_;
  assign N3442 = ~pe_o_4__6_;
  assign N3443 = ~pe_o_4__5_;
  assign N3444 = ~pe_o_4__3_;
  assign N3445 = ~pe_o_4__0_;
  assign N3446 = N3451 & N3452;
  assign N3447 = N3446 & pe_o_4__4_;
  assign N3448 = N3447 & N3453;
  assign N3449 = N3448 & pe_o_4__2_;
  assign N3450 = N3449 & pe_o_4__0_;
  assign N8109 = N3450 & pe_o_4__1_;
  assign N3451 = ~pe_o_4__6_;
  assign N3452 = ~pe_o_4__5_;
  assign N3453 = ~pe_o_4__3_;
  assign N3454 = N3459 & N3460;
  assign N3455 = N3454 & pe_o_4__4_;
  assign N3456 = N3455 & pe_o_4__3_;
  assign N3457 = N3456 & N3461;
  assign N3458 = N3457 & N3462;
  assign N8111 = N3458 & N3463;
  assign N3459 = ~pe_o_4__6_;
  assign N3460 = ~pe_o_4__5_;
  assign N3461 = ~pe_o_4__2_;
  assign N3462 = ~pe_o_4__0_;
  assign N3463 = ~pe_o_4__1_;
  assign N3464 = N3469 & N3470;
  assign N3465 = N3464 & pe_o_4__4_;
  assign N3466 = N3465 & pe_o_4__3_;
  assign N3467 = N3466 & N3471;
  assign N3468 = N3467 & pe_o_4__0_;
  assign N8113 = N3468 & N3472;
  assign N3469 = ~pe_o_4__6_;
  assign N3470 = ~pe_o_4__5_;
  assign N3471 = ~pe_o_4__2_;
  assign N3472 = ~pe_o_4__1_;
  assign N3473 = N3478 & N3479;
  assign N3474 = N3473 & pe_o_4__4_;
  assign N3475 = N3474 & pe_o_4__3_;
  assign N3476 = N3475 & N3480;
  assign N3477 = N3476 & N3481;
  assign N8115 = N3477 & pe_o_4__1_;
  assign N3478 = ~pe_o_4__6_;
  assign N3479 = ~pe_o_4__5_;
  assign N3480 = ~pe_o_4__2_;
  assign N3481 = ~pe_o_4__0_;
  assign N3482 = N3487 & N3488;
  assign N3483 = N3482 & pe_o_4__4_;
  assign N3484 = N3483 & pe_o_4__3_;
  assign N3485 = N3484 & N3489;
  assign N3486 = N3485 & pe_o_4__0_;
  assign N8117 = N3486 & pe_o_4__1_;
  assign N3487 = ~pe_o_4__6_;
  assign N3488 = ~pe_o_4__5_;
  assign N3489 = ~pe_o_4__2_;
  assign N3490 = N3495 & N3496;
  assign N3491 = N3490 & pe_o_4__4_;
  assign N3492 = N3491 & pe_o_4__3_;
  assign N3493 = N3492 & pe_o_4__2_;
  assign N3494 = N3493 & N3497;
  assign N8119 = N3494 & N3498;
  assign N3495 = ~pe_o_4__6_;
  assign N3496 = ~pe_o_4__5_;
  assign N3497 = ~pe_o_4__0_;
  assign N3498 = ~pe_o_4__1_;
  assign N3499 = N3504 & N3505;
  assign N3500 = N3499 & pe_o_4__4_;
  assign N3501 = N3500 & pe_o_4__3_;
  assign N3502 = N3501 & pe_o_4__2_;
  assign N3503 = N3502 & pe_o_4__0_;
  assign N8121 = N3503 & N3506;
  assign N3504 = ~pe_o_4__6_;
  assign N3505 = ~pe_o_4__5_;
  assign N3506 = ~pe_o_4__1_;
  assign N3507 = N3512 & N3513;
  assign N3508 = N3507 & pe_o_4__4_;
  assign N3509 = N3508 & pe_o_4__3_;
  assign N3510 = N3509 & pe_o_4__2_;
  assign N3511 = N3510 & N3514;
  assign N8123 = N3511 & pe_o_4__1_;
  assign N3512 = ~pe_o_4__6_;
  assign N3513 = ~pe_o_4__5_;
  assign N3514 = ~pe_o_4__0_;
  assign N3515 = N3520 & N3521;
  assign N3516 = N3515 & pe_o_4__4_;
  assign N3517 = N3516 & pe_o_4__3_;
  assign N3518 = N3517 & pe_o_4__2_;
  assign N3519 = N3518 & pe_o_4__0_;
  assign N8125 = N3519 & pe_o_4__1_;
  assign N3520 = ~pe_o_4__6_;
  assign N3521 = ~pe_o_4__5_;
  assign N3522 = N3527 & pe_o_4__5_;
  assign N3523 = N3522 & N3528;
  assign N3524 = N3523 & N3529;
  assign N3525 = N3524 & N3530;
  assign N3526 = N3525 & N3531;
  assign N8127 = N3526 & N3532;
  assign N3527 = ~pe_o_4__6_;
  assign N3528 = ~pe_o_4__4_;
  assign N3529 = ~pe_o_4__3_;
  assign N3530 = ~pe_o_4__2_;
  assign N3531 = ~pe_o_4__0_;
  assign N3532 = ~pe_o_4__1_;
  assign N3533 = N3538 & pe_o_4__5_;
  assign N3534 = N3533 & N3539;
  assign N3535 = N3534 & N3540;
  assign N3536 = N3535 & N3541;
  assign N3537 = N3536 & pe_o_4__0_;
  assign N8129 = N3537 & N3542;
  assign N3538 = ~pe_o_4__6_;
  assign N3539 = ~pe_o_4__4_;
  assign N3540 = ~pe_o_4__3_;
  assign N3541 = ~pe_o_4__2_;
  assign N3542 = ~pe_o_4__1_;
  assign N3543 = N3548 & pe_o_4__5_;
  assign N3544 = N3543 & N3549;
  assign N3545 = N3544 & N3550;
  assign N3546 = N3545 & N3551;
  assign N3547 = N3546 & N3552;
  assign N8131 = N3547 & pe_o_4__1_;
  assign N3548 = ~pe_o_4__6_;
  assign N3549 = ~pe_o_4__4_;
  assign N3550 = ~pe_o_4__3_;
  assign N3551 = ~pe_o_4__2_;
  assign N3552 = ~pe_o_4__0_;
  assign N3553 = N3558 & pe_o_4__5_;
  assign N3554 = N3553 & N3559;
  assign N3555 = N3554 & N3560;
  assign N3556 = N3555 & N3561;
  assign N3557 = N3556 & pe_o_4__0_;
  assign N8133 = N3557 & pe_o_4__1_;
  assign N3558 = ~pe_o_4__6_;
  assign N3559 = ~pe_o_4__4_;
  assign N3560 = ~pe_o_4__3_;
  assign N3561 = ~pe_o_4__2_;
  assign N3562 = N3567 & pe_o_4__5_;
  assign N3563 = N3562 & N3568;
  assign N3564 = N3563 & N3569;
  assign N3565 = N3564 & pe_o_4__2_;
  assign N3566 = N3565 & N3570;
  assign N8135 = N3566 & N3571;
  assign N3567 = ~pe_o_4__6_;
  assign N3568 = ~pe_o_4__4_;
  assign N3569 = ~pe_o_4__3_;
  assign N3570 = ~pe_o_4__0_;
  assign N3571 = ~pe_o_4__1_;
  assign N3572 = N3577 & pe_o_4__5_;
  assign N3573 = N3572 & N3578;
  assign N3574 = N3573 & N3579;
  assign N3575 = N3574 & pe_o_4__2_;
  assign N3576 = N3575 & pe_o_4__0_;
  assign N8137 = N3576 & N3580;
  assign N3577 = ~pe_o_4__6_;
  assign N3578 = ~pe_o_4__4_;
  assign N3579 = ~pe_o_4__3_;
  assign N3580 = ~pe_o_4__1_;
  assign N3581 = N3586 & pe_o_4__5_;
  assign N3582 = N3581 & N3587;
  assign N3583 = N3582 & N3588;
  assign N3584 = N3583 & pe_o_4__2_;
  assign N3585 = N3584 & N3589;
  assign N8139 = N3585 & pe_o_4__1_;
  assign N3586 = ~pe_o_4__6_;
  assign N3587 = ~pe_o_4__4_;
  assign N3588 = ~pe_o_4__3_;
  assign N3589 = ~pe_o_4__0_;
  assign N3590 = N3595 & pe_o_4__5_;
  assign N3591 = N3590 & N3596;
  assign N3592 = N3591 & N3597;
  assign N3593 = N3592 & pe_o_4__2_;
  assign N3594 = N3593 & pe_o_4__0_;
  assign N8141 = N3594 & pe_o_4__1_;
  assign N3595 = ~pe_o_4__6_;
  assign N3596 = ~pe_o_4__4_;
  assign N3597 = ~pe_o_4__3_;
  assign N3598 = N3603 & pe_o_4__5_;
  assign N3599 = N3598 & N3604;
  assign N3600 = N3599 & pe_o_4__3_;
  assign N3601 = N3600 & N3605;
  assign N3602 = N3601 & N3606;
  assign N8143 = N3602 & N3607;
  assign N3603 = ~pe_o_4__6_;
  assign N3604 = ~pe_o_4__4_;
  assign N3605 = ~pe_o_4__2_;
  assign N3606 = ~pe_o_4__0_;
  assign N3607 = ~pe_o_4__1_;
  assign N3608 = N3613 & pe_o_4__5_;
  assign N3609 = N3608 & N3614;
  assign N3610 = N3609 & pe_o_4__3_;
  assign N3611 = N3610 & N3615;
  assign N3612 = N3611 & pe_o_4__0_;
  assign N8145 = N3612 & N3616;
  assign N3613 = ~pe_o_4__6_;
  assign N3614 = ~pe_o_4__4_;
  assign N3615 = ~pe_o_4__2_;
  assign N3616 = ~pe_o_4__1_;
  assign N3617 = N3622 & pe_o_4__5_;
  assign N3618 = N3617 & N3623;
  assign N3619 = N3618 & pe_o_4__3_;
  assign N3620 = N3619 & N3624;
  assign N3621 = N3620 & N3625;
  assign N8147 = N3621 & pe_o_4__1_;
  assign N3622 = ~pe_o_4__6_;
  assign N3623 = ~pe_o_4__4_;
  assign N3624 = ~pe_o_4__2_;
  assign N3625 = ~pe_o_4__0_;
  assign N3626 = N3631 & pe_o_4__5_;
  assign N3627 = N3626 & N3632;
  assign N3628 = N3627 & pe_o_4__3_;
  assign N3629 = N3628 & N3633;
  assign N3630 = N3629 & pe_o_4__0_;
  assign N8149 = N3630 & pe_o_4__1_;
  assign N3631 = ~pe_o_4__6_;
  assign N3632 = ~pe_o_4__4_;
  assign N3633 = ~pe_o_4__2_;
  assign N3634 = N3639 & pe_o_4__5_;
  assign N3635 = N3634 & N3640;
  assign N3636 = N3635 & pe_o_4__3_;
  assign N3637 = N3636 & pe_o_4__2_;
  assign N3638 = N3637 & N3641;
  assign N8151 = N3638 & N3642;
  assign N3639 = ~pe_o_4__6_;
  assign N3640 = ~pe_o_4__4_;
  assign N3641 = ~pe_o_4__0_;
  assign N3642 = ~pe_o_4__1_;
  assign N3643 = N3648 & pe_o_4__5_;
  assign N3644 = N3643 & N3649;
  assign N3645 = N3644 & pe_o_4__3_;
  assign N3646 = N3645 & pe_o_4__2_;
  assign N3647 = N3646 & pe_o_4__0_;
  assign N8153 = N3647 & N3650;
  assign N3648 = ~pe_o_4__6_;
  assign N3649 = ~pe_o_4__4_;
  assign N3650 = ~pe_o_4__1_;
  assign N3651 = N3656 & pe_o_4__5_;
  assign N3652 = N3651 & N3657;
  assign N3653 = N3652 & pe_o_4__3_;
  assign N3654 = N3653 & pe_o_4__2_;
  assign N3655 = N3654 & N3658;
  assign N8155 = N3655 & pe_o_4__1_;
  assign N3656 = ~pe_o_4__6_;
  assign N3657 = ~pe_o_4__4_;
  assign N3658 = ~pe_o_4__0_;
  assign N3659 = N3664 & pe_o_4__5_;
  assign N3660 = N3659 & N3665;
  assign N3661 = N3660 & pe_o_4__3_;
  assign N3662 = N3661 & pe_o_4__2_;
  assign N3663 = N3662 & pe_o_4__0_;
  assign N8157 = N3663 & pe_o_4__1_;
  assign N3664 = ~pe_o_4__6_;
  assign N3665 = ~pe_o_4__4_;
  assign N3666 = N3671 & pe_o_4__5_;
  assign N3667 = N3666 & pe_o_4__4_;
  assign N3668 = N3667 & N3672;
  assign N3669 = N3668 & N3673;
  assign N3670 = N3669 & N3674;
  assign N8159 = N3670 & N3675;
  assign N3671 = ~pe_o_4__6_;
  assign N3672 = ~pe_o_4__3_;
  assign N3673 = ~pe_o_4__2_;
  assign N3674 = ~pe_o_4__0_;
  assign N3675 = ~pe_o_4__1_;
  assign N3676 = N3681 & pe_o_4__5_;
  assign N3677 = N3676 & pe_o_4__4_;
  assign N3678 = N3677 & N3682;
  assign N3679 = N3678 & N3683;
  assign N3680 = N3679 & pe_o_4__0_;
  assign N8161 = N3680 & N3684;
  assign N3681 = ~pe_o_4__6_;
  assign N3682 = ~pe_o_4__3_;
  assign N3683 = ~pe_o_4__2_;
  assign N3684 = ~pe_o_4__1_;
  assign N3685 = N3690 & pe_o_4__5_;
  assign N3686 = N3685 & pe_o_4__4_;
  assign N3687 = N3686 & N3691;
  assign N3688 = N3687 & N3692;
  assign N3689 = N3688 & N3693;
  assign N8163 = N3689 & pe_o_4__1_;
  assign N3690 = ~pe_o_4__6_;
  assign N3691 = ~pe_o_4__3_;
  assign N3692 = ~pe_o_4__2_;
  assign N3693 = ~pe_o_4__0_;
  assign N3694 = N3699 & pe_o_4__5_;
  assign N3695 = N3694 & pe_o_4__4_;
  assign N3696 = N3695 & N3700;
  assign N3697 = N3696 & N3701;
  assign N3698 = N3697 & pe_o_4__0_;
  assign N8165 = N3698 & pe_o_4__1_;
  assign N3699 = ~pe_o_4__6_;
  assign N3700 = ~pe_o_4__3_;
  assign N3701 = ~pe_o_4__2_;
  assign N3702 = N3707 & pe_o_4__5_;
  assign N3703 = N3702 & pe_o_4__4_;
  assign N3704 = N3703 & N3708;
  assign N3705 = N3704 & pe_o_4__2_;
  assign N3706 = N3705 & N3709;
  assign N8167 = N3706 & N3710;
  assign N3707 = ~pe_o_4__6_;
  assign N3708 = ~pe_o_4__3_;
  assign N3709 = ~pe_o_4__0_;
  assign N3710 = ~pe_o_4__1_;
  assign N3711 = N3716 & pe_o_4__5_;
  assign N3712 = N3711 & pe_o_4__4_;
  assign N3713 = N3712 & N3717;
  assign N3714 = N3713 & pe_o_4__2_;
  assign N3715 = N3714 & pe_o_4__0_;
  assign N8169 = N3715 & N3718;
  assign N3716 = ~pe_o_4__6_;
  assign N3717 = ~pe_o_4__3_;
  assign N3718 = ~pe_o_4__1_;
  assign N3719 = N3724 & pe_o_4__5_;
  assign N3720 = N3719 & pe_o_4__4_;
  assign N3721 = N3720 & N3725;
  assign N3722 = N3721 & pe_o_4__2_;
  assign N3723 = N3722 & N3726;
  assign N8171 = N3723 & pe_o_4__1_;
  assign N3724 = ~pe_o_4__6_;
  assign N3725 = ~pe_o_4__3_;
  assign N3726 = ~pe_o_4__0_;
  assign N3727 = N3732 & pe_o_4__5_;
  assign N3728 = N3727 & pe_o_4__4_;
  assign N3729 = N3728 & N3733;
  assign N3730 = N3729 & pe_o_4__2_;
  assign N3731 = N3730 & pe_o_4__0_;
  assign N8173 = N3731 & pe_o_4__1_;
  assign N3732 = ~pe_o_4__6_;
  assign N3733 = ~pe_o_4__3_;
  assign N3734 = N3739 & pe_o_4__5_;
  assign N3735 = N3734 & pe_o_4__4_;
  assign N3736 = N3735 & pe_o_4__3_;
  assign N3737 = N3736 & N3740;
  assign N3738 = N3737 & N3741;
  assign N8175 = N3738 & N3742;
  assign N3739 = ~pe_o_4__6_;
  assign N3740 = ~pe_o_4__2_;
  assign N3741 = ~pe_o_4__0_;
  assign N3742 = ~pe_o_4__1_;
  assign N3743 = N3748 & pe_o_4__5_;
  assign N3744 = N3743 & pe_o_4__4_;
  assign N3745 = N3744 & pe_o_4__3_;
  assign N3746 = N3745 & N3749;
  assign N3747 = N3746 & pe_o_4__0_;
  assign N8177 = N3747 & N3750;
  assign N3748 = ~pe_o_4__6_;
  assign N3749 = ~pe_o_4__2_;
  assign N3750 = ~pe_o_4__1_;
  assign N3751 = N3756 & pe_o_4__5_;
  assign N3752 = N3751 & pe_o_4__4_;
  assign N3753 = N3752 & pe_o_4__3_;
  assign N3754 = N3753 & N3757;
  assign N3755 = N3754 & N3758;
  assign N8179 = N3755 & pe_o_4__1_;
  assign N3756 = ~pe_o_4__6_;
  assign N3757 = ~pe_o_4__2_;
  assign N3758 = ~pe_o_4__0_;
  assign N3759 = N3764 & pe_o_4__5_;
  assign N3760 = N3759 & pe_o_4__4_;
  assign N3761 = N3760 & pe_o_4__3_;
  assign N3762 = N3761 & N3765;
  assign N3763 = N3762 & pe_o_4__0_;
  assign N8181 = N3763 & pe_o_4__1_;
  assign N3764 = ~pe_o_4__6_;
  assign N3765 = ~pe_o_4__2_;
  assign N3766 = N3771 & pe_o_4__5_;
  assign N3767 = N3766 & pe_o_4__4_;
  assign N3768 = N3767 & pe_o_4__3_;
  assign N3769 = N3768 & pe_o_4__2_;
  assign N3770 = N3769 & N3772;
  assign N8183 = N3770 & N3773;
  assign N3771 = ~pe_o_4__6_;
  assign N3772 = ~pe_o_4__0_;
  assign N3773 = ~pe_o_4__1_;
  assign N3774 = N3779 & pe_o_4__5_;
  assign N3775 = N3774 & pe_o_4__4_;
  assign N3776 = N3775 & pe_o_4__3_;
  assign N3777 = N3776 & pe_o_4__2_;
  assign N3778 = N3777 & pe_o_4__0_;
  assign N8185 = N3778 & N3780;
  assign N3779 = ~pe_o_4__6_;
  assign N3780 = ~pe_o_4__1_;
  assign N3781 = N3786 & pe_o_4__5_;
  assign N3782 = N3781 & pe_o_4__4_;
  assign N3783 = N3782 & pe_o_4__3_;
  assign N3784 = N3783 & pe_o_4__2_;
  assign N3785 = N3784 & N3787;
  assign N8187 = N3785 & pe_o_4__1_;
  assign N3786 = ~pe_o_4__6_;
  assign N3787 = ~pe_o_4__0_;
  assign N3788 = pe_o_4__5_ & pe_o_4__4_;
  assign N3789 = N3788 & pe_o_4__3_;
  assign N3790 = N3789 & pe_o_4__2_;
  assign N3791 = N3790 & pe_o_4__0_;
  assign N8189 = N3791 & pe_o_4__1_;
  assign N3792 = pe_o_4__6_ & N3797;
  assign N3793 = N3792 & N3798;
  assign N3794 = N3793 & N3799;
  assign N3795 = N3794 & N3800;
  assign N3796 = N3795 & pe_o_4__0_;
  assign N8066 = N3796 & N3801;
  assign N3797 = ~pe_o_4__5_;
  assign N3798 = ~pe_o_4__4_;
  assign N3799 = ~pe_o_4__3_;
  assign N3800 = ~pe_o_4__2_;
  assign N3801 = ~pe_o_4__1_;
  assign N3802 = pe_o_4__6_ & N3807;
  assign N3803 = N3802 & N3808;
  assign N3804 = N3803 & N3809;
  assign N3805 = N3804 & N3810;
  assign N3806 = N3805 & N3811;
  assign N8068 = N3806 & pe_o_4__1_;
  assign N3807 = ~pe_o_4__5_;
  assign N3808 = ~pe_o_4__4_;
  assign N3809 = ~pe_o_4__3_;
  assign N3810 = ~pe_o_4__2_;
  assign N3811 = ~pe_o_4__0_;
  assign N3812 = pe_o_4__6_ & N3817;
  assign N3813 = N3812 & N3818;
  assign N3814 = N3813 & N3819;
  assign N3815 = N3814 & N3820;
  assign N3816 = N3815 & pe_o_4__0_;
  assign N8070 = N3816 & pe_o_4__1_;
  assign N3817 = ~pe_o_4__5_;
  assign N3818 = ~pe_o_4__4_;
  assign N3819 = ~pe_o_4__3_;
  assign N3820 = ~pe_o_4__2_;
  assign N3821 = pe_o_4__6_ & N3826;
  assign N3822 = N3821 & N3827;
  assign N3823 = N3822 & N3828;
  assign N3824 = N3823 & pe_o_4__2_;
  assign N3825 = N3824 & N3829;
  assign N8072 = N3825 & N3830;
  assign N3826 = ~pe_o_4__5_;
  assign N3827 = ~pe_o_4__4_;
  assign N3828 = ~pe_o_4__3_;
  assign N3829 = ~pe_o_4__0_;
  assign N3830 = ~pe_o_4__1_;
  assign N3831 = pe_o_4__6_ & N3836;
  assign N3832 = N3831 & N3837;
  assign N3833 = N3832 & N3838;
  assign N3834 = N3833 & pe_o_4__2_;
  assign N3835 = N3834 & pe_o_4__0_;
  assign N8074 = N3835 & N3839;
  assign N3836 = ~pe_o_4__5_;
  assign N3837 = ~pe_o_4__4_;
  assign N3838 = ~pe_o_4__3_;
  assign N3839 = ~pe_o_4__1_;
  assign N3840 = pe_o_4__6_ & N3845;
  assign N3841 = N3840 & N3846;
  assign N3842 = N3841 & N3847;
  assign N3843 = N3842 & pe_o_4__2_;
  assign N3844 = N3843 & N3848;
  assign N8076 = N3844 & pe_o_4__1_;
  assign N3845 = ~pe_o_4__5_;
  assign N3846 = ~pe_o_4__4_;
  assign N3847 = ~pe_o_4__3_;
  assign N3848 = ~pe_o_4__0_;
  assign N3849 = pe_o_4__6_ & N3854;
  assign N3850 = N3849 & N3855;
  assign N3851 = N3850 & N3856;
  assign N3852 = N3851 & pe_o_4__2_;
  assign N3853 = N3852 & pe_o_4__0_;
  assign N8078 = N3853 & pe_o_4__1_;
  assign N3854 = ~pe_o_4__5_;
  assign N3855 = ~pe_o_4__4_;
  assign N3856 = ~pe_o_4__3_;
  assign N3857 = pe_o_4__6_ & N3862;
  assign N3858 = N3857 & N3863;
  assign N3859 = N3858 & pe_o_4__3_;
  assign N3860 = N3859 & N3864;
  assign N3861 = N3860 & N3865;
  assign N8080 = N3861 & N3866;
  assign N3862 = ~pe_o_4__5_;
  assign N3863 = ~pe_o_4__4_;
  assign N3864 = ~pe_o_4__2_;
  assign N3865 = ~pe_o_4__0_;
  assign N3866 = ~pe_o_4__1_;
  assign N3867 = pe_o_4__6_ & N3872;
  assign N3868 = N3867 & N3873;
  assign N3869 = N3868 & pe_o_4__3_;
  assign N3870 = N3869 & N3874;
  assign N3871 = N3870 & pe_o_4__0_;
  assign N8082 = N3871 & N3875;
  assign N3872 = ~pe_o_4__5_;
  assign N3873 = ~pe_o_4__4_;
  assign N3874 = ~pe_o_4__2_;
  assign N3875 = ~pe_o_4__1_;
  assign N3876 = pe_o_4__6_ & N3881;
  assign N3877 = N3876 & N3882;
  assign N3878 = N3877 & pe_o_4__3_;
  assign N3879 = N3878 & N3883;
  assign N3880 = N3879 & N3884;
  assign N8084 = N3880 & pe_o_4__1_;
  assign N3881 = ~pe_o_4__5_;
  assign N3882 = ~pe_o_4__4_;
  assign N3883 = ~pe_o_4__2_;
  assign N3884 = ~pe_o_4__0_;
  assign N3885 = pe_o_4__6_ & N3890;
  assign N3886 = N3885 & N3891;
  assign N3887 = N3886 & pe_o_4__3_;
  assign N3888 = N3887 & N3892;
  assign N3889 = N3888 & pe_o_4__0_;
  assign N8086 = N3889 & pe_o_4__1_;
  assign N3890 = ~pe_o_4__5_;
  assign N3891 = ~pe_o_4__4_;
  assign N3892 = ~pe_o_4__2_;
  assign N3893 = pe_o_4__6_ & N3898;
  assign N3894 = N3893 & N3899;
  assign N3895 = N3894 & pe_o_4__3_;
  assign N3896 = N3895 & pe_o_4__2_;
  assign N3897 = N3896 & N3900;
  assign N8088 = N3897 & N3901;
  assign N3898 = ~pe_o_4__5_;
  assign N3899 = ~pe_o_4__4_;
  assign N3900 = ~pe_o_4__0_;
  assign N3901 = ~pe_o_4__1_;
  assign N3902 = pe_o_4__6_ & N3907;
  assign N3903 = N3902 & N3908;
  assign N3904 = N3903 & pe_o_4__3_;
  assign N3905 = N3904 & pe_o_4__2_;
  assign N3906 = N3905 & pe_o_4__0_;
  assign N8090 = N3906 & N3909;
  assign N3907 = ~pe_o_4__5_;
  assign N3908 = ~pe_o_4__4_;
  assign N3909 = ~pe_o_4__1_;
  assign N3910 = pe_o_4__6_ & N3915;
  assign N3911 = N3910 & N3916;
  assign N3912 = N3911 & pe_o_4__3_;
  assign N3913 = N3912 & pe_o_4__2_;
  assign N3914 = N3913 & N3917;
  assign N8092 = N3914 & pe_o_4__1_;
  assign N3915 = ~pe_o_4__5_;
  assign N3916 = ~pe_o_4__4_;
  assign N3917 = ~pe_o_4__0_;
  assign N3918 = pe_o_4__6_ & N3923;
  assign N3919 = N3918 & N3924;
  assign N3920 = N3919 & pe_o_4__3_;
  assign N3921 = N3920 & pe_o_4__2_;
  assign N3922 = N3921 & pe_o_4__0_;
  assign N8094 = N3922 & pe_o_4__1_;
  assign N3923 = ~pe_o_4__5_;
  assign N3924 = ~pe_o_4__4_;
  assign N3925 = pe_o_4__6_ & N3930;
  assign N3926 = N3925 & pe_o_4__4_;
  assign N3927 = N3926 & N3931;
  assign N3928 = N3927 & N3932;
  assign N3929 = N3928 & N3933;
  assign N8096 = N3929 & N3934;
  assign N3930 = ~pe_o_4__5_;
  assign N3931 = ~pe_o_4__3_;
  assign N3932 = ~pe_o_4__2_;
  assign N3933 = ~pe_o_4__0_;
  assign N3934 = ~pe_o_4__1_;
  assign N3935 = pe_o_4__6_ & N3940;
  assign N3936 = N3935 & pe_o_4__4_;
  assign N3937 = N3936 & N3941;
  assign N3938 = N3937 & N3942;
  assign N3939 = N3938 & pe_o_4__0_;
  assign N8098 = N3939 & N3943;
  assign N3940 = ~pe_o_4__5_;
  assign N3941 = ~pe_o_4__3_;
  assign N3942 = ~pe_o_4__2_;
  assign N3943 = ~pe_o_4__1_;
  assign N3944 = pe_o_4__6_ & N3949;
  assign N3945 = N3944 & pe_o_4__4_;
  assign N3946 = N3945 & N3950;
  assign N3947 = N3946 & N3951;
  assign N3948 = N3947 & N3952;
  assign N8100 = N3948 & pe_o_4__1_;
  assign N3949 = ~pe_o_4__5_;
  assign N3950 = ~pe_o_4__3_;
  assign N3951 = ~pe_o_4__2_;
  assign N3952 = ~pe_o_4__0_;
  assign N3953 = pe_o_4__6_ & N3958;
  assign N3954 = N3953 & pe_o_4__4_;
  assign N3955 = N3954 & N3959;
  assign N3956 = N3955 & N3960;
  assign N3957 = N3956 & pe_o_4__0_;
  assign N8102 = N3957 & pe_o_4__1_;
  assign N3958 = ~pe_o_4__5_;
  assign N3959 = ~pe_o_4__3_;
  assign N3960 = ~pe_o_4__2_;
  assign N3961 = pe_o_4__6_ & N3966;
  assign N3962 = N3961 & pe_o_4__4_;
  assign N3963 = N3962 & N3967;
  assign N3964 = N3963 & pe_o_4__2_;
  assign N3965 = N3964 & N3968;
  assign N8104 = N3965 & N3969;
  assign N3966 = ~pe_o_4__5_;
  assign N3967 = ~pe_o_4__3_;
  assign N3968 = ~pe_o_4__0_;
  assign N3969 = ~pe_o_4__1_;
  assign N3970 = pe_o_4__6_ & N3975;
  assign N3971 = N3970 & pe_o_4__4_;
  assign N3972 = N3971 & N3976;
  assign N3973 = N3972 & pe_o_4__2_;
  assign N3974 = N3973 & pe_o_4__0_;
  assign N8106 = N3974 & N3977;
  assign N3975 = ~pe_o_4__5_;
  assign N3976 = ~pe_o_4__3_;
  assign N3977 = ~pe_o_4__1_;
  assign N3978 = pe_o_4__6_ & N3983;
  assign N3979 = N3978 & pe_o_4__4_;
  assign N3980 = N3979 & N3984;
  assign N3981 = N3980 & pe_o_4__2_;
  assign N3982 = N3981 & N3985;
  assign N8108 = N3982 & pe_o_4__1_;
  assign N3983 = ~pe_o_4__5_;
  assign N3984 = ~pe_o_4__3_;
  assign N3985 = ~pe_o_4__0_;
  assign N3986 = pe_o_4__6_ & N3991;
  assign N3987 = N3986 & pe_o_4__4_;
  assign N3988 = N3987 & N3992;
  assign N3989 = N3988 & pe_o_4__2_;
  assign N3990 = N3989 & pe_o_4__0_;
  assign N8110 = N3990 & pe_o_4__1_;
  assign N3991 = ~pe_o_4__5_;
  assign N3992 = ~pe_o_4__3_;
  assign N3993 = pe_o_4__6_ & N3998;
  assign N3994 = N3993 & pe_o_4__4_;
  assign N3995 = N3994 & pe_o_4__3_;
  assign N3996 = N3995 & N3999;
  assign N3997 = N3996 & N4000;
  assign N8112 = N3997 & N4001;
  assign N3998 = ~pe_o_4__5_;
  assign N3999 = ~pe_o_4__2_;
  assign N4000 = ~pe_o_4__0_;
  assign N4001 = ~pe_o_4__1_;
  assign N4002 = pe_o_4__6_ & N4007;
  assign N4003 = N4002 & pe_o_4__4_;
  assign N4004 = N4003 & pe_o_4__3_;
  assign N4005 = N4004 & N4008;
  assign N4006 = N4005 & pe_o_4__0_;
  assign N8114 = N4006 & N4009;
  assign N4007 = ~pe_o_4__5_;
  assign N4008 = ~pe_o_4__2_;
  assign N4009 = ~pe_o_4__1_;
  assign N4010 = pe_o_4__6_ & N4015;
  assign N4011 = N4010 & pe_o_4__4_;
  assign N4012 = N4011 & pe_o_4__3_;
  assign N4013 = N4012 & N4016;
  assign N4014 = N4013 & N4017;
  assign N8116 = N4014 & pe_o_4__1_;
  assign N4015 = ~pe_o_4__5_;
  assign N4016 = ~pe_o_4__2_;
  assign N4017 = ~pe_o_4__0_;
  assign N4018 = pe_o_4__6_ & N4023;
  assign N4019 = N4018 & pe_o_4__4_;
  assign N4020 = N4019 & pe_o_4__3_;
  assign N4021 = N4020 & N4024;
  assign N4022 = N4021 & pe_o_4__0_;
  assign N8118 = N4022 & pe_o_4__1_;
  assign N4023 = ~pe_o_4__5_;
  assign N4024 = ~pe_o_4__2_;
  assign N4025 = pe_o_4__6_ & N4030;
  assign N4026 = N4025 & pe_o_4__4_;
  assign N4027 = N4026 & pe_o_4__3_;
  assign N4028 = N4027 & pe_o_4__2_;
  assign N4029 = N4028 & N4031;
  assign N8120 = N4029 & N4032;
  assign N4030 = ~pe_o_4__5_;
  assign N4031 = ~pe_o_4__0_;
  assign N4032 = ~pe_o_4__1_;
  assign N4033 = pe_o_4__6_ & N4038;
  assign N4034 = N4033 & pe_o_4__4_;
  assign N4035 = N4034 & pe_o_4__3_;
  assign N4036 = N4035 & pe_o_4__2_;
  assign N4037 = N4036 & pe_o_4__0_;
  assign N8122 = N4037 & N4039;
  assign N4038 = ~pe_o_4__5_;
  assign N4039 = ~pe_o_4__1_;
  assign N4040 = pe_o_4__6_ & N4045;
  assign N4041 = N4040 & pe_o_4__4_;
  assign N4042 = N4041 & pe_o_4__3_;
  assign N4043 = N4042 & pe_o_4__2_;
  assign N4044 = N4043 & N4046;
  assign N8124 = N4044 & pe_o_4__1_;
  assign N4045 = ~pe_o_4__5_;
  assign N4046 = ~pe_o_4__0_;
  assign N4047 = pe_o_4__6_ & pe_o_4__4_;
  assign N4048 = N4047 & pe_o_4__3_;
  assign N4049 = N4048 & pe_o_4__2_;
  assign N4050 = N4049 & pe_o_4__0_;
  assign N8126 = N4050 & pe_o_4__1_;
  assign N4051 = pe_o_4__6_ & pe_o_4__5_;
  assign N4052 = N4051 & N4056;
  assign N4053 = N4052 & N4057;
  assign N4054 = N4053 & N4058;
  assign N4055 = N4054 & N4059;
  assign N8128 = N4055 & N4060;
  assign N4056 = ~pe_o_4__4_;
  assign N4057 = ~pe_o_4__3_;
  assign N4058 = ~pe_o_4__2_;
  assign N4059 = ~pe_o_4__0_;
  assign N4060 = ~pe_o_4__1_;
  assign N4061 = pe_o_4__6_ & pe_o_4__5_;
  assign N4062 = N4061 & N4066;
  assign N4063 = N4062 & N4067;
  assign N4064 = N4063 & N4068;
  assign N4065 = N4064 & pe_o_4__0_;
  assign N8130 = N4065 & N4069;
  assign N4066 = ~pe_o_4__4_;
  assign N4067 = ~pe_o_4__3_;
  assign N4068 = ~pe_o_4__2_;
  assign N4069 = ~pe_o_4__1_;
  assign N4070 = pe_o_4__6_ & pe_o_4__5_;
  assign N4071 = N4070 & N4075;
  assign N4072 = N4071 & N4076;
  assign N4073 = N4072 & N4077;
  assign N4074 = N4073 & N4078;
  assign N8132 = N4074 & pe_o_4__1_;
  assign N4075 = ~pe_o_4__4_;
  assign N4076 = ~pe_o_4__3_;
  assign N4077 = ~pe_o_4__2_;
  assign N4078 = ~pe_o_4__0_;
  assign N4079 = pe_o_4__6_ & pe_o_4__5_;
  assign N4080 = N4079 & N4084;
  assign N4081 = N4080 & N4085;
  assign N4082 = N4081 & N4086;
  assign N4083 = N4082 & pe_o_4__0_;
  assign N8134 = N4083 & pe_o_4__1_;
  assign N4084 = ~pe_o_4__4_;
  assign N4085 = ~pe_o_4__3_;
  assign N4086 = ~pe_o_4__2_;
  assign N4087 = pe_o_4__6_ & pe_o_4__5_;
  assign N4088 = N4087 & N4092;
  assign N4089 = N4088 & N4093;
  assign N4090 = N4089 & pe_o_4__2_;
  assign N4091 = N4090 & N4094;
  assign N8136 = N4091 & N4095;
  assign N4092 = ~pe_o_4__4_;
  assign N4093 = ~pe_o_4__3_;
  assign N4094 = ~pe_o_4__0_;
  assign N4095 = ~pe_o_4__1_;
  assign N4096 = pe_o_4__6_ & pe_o_4__5_;
  assign N4097 = N4096 & N4101;
  assign N4098 = N4097 & N4102;
  assign N4099 = N4098 & pe_o_4__2_;
  assign N4100 = N4099 & pe_o_4__0_;
  assign N8138 = N4100 & N4103;
  assign N4101 = ~pe_o_4__4_;
  assign N4102 = ~pe_o_4__3_;
  assign N4103 = ~pe_o_4__1_;
  assign N4104 = pe_o_4__6_ & pe_o_4__5_;
  assign N4105 = N4104 & N4109;
  assign N4106 = N4105 & N4110;
  assign N4107 = N4106 & pe_o_4__2_;
  assign N4108 = N4107 & N4111;
  assign N8140 = N4108 & pe_o_4__1_;
  assign N4109 = ~pe_o_4__4_;
  assign N4110 = ~pe_o_4__3_;
  assign N4111 = ~pe_o_4__0_;
  assign N4112 = pe_o_4__6_ & pe_o_4__5_;
  assign N4113 = N4112 & N4117;
  assign N4114 = N4113 & N4118;
  assign N4115 = N4114 & pe_o_4__2_;
  assign N4116 = N4115 & pe_o_4__0_;
  assign N8142 = N4116 & pe_o_4__1_;
  assign N4117 = ~pe_o_4__4_;
  assign N4118 = ~pe_o_4__3_;
  assign N4119 = pe_o_4__6_ & pe_o_4__5_;
  assign N4120 = N4119 & N4124;
  assign N4121 = N4120 & pe_o_4__3_;
  assign N4122 = N4121 & N4125;
  assign N4123 = N4122 & N4126;
  assign N8144 = N4123 & N4127;
  assign N4124 = ~pe_o_4__4_;
  assign N4125 = ~pe_o_4__2_;
  assign N4126 = ~pe_o_4__0_;
  assign N4127 = ~pe_o_4__1_;
  assign N4128 = pe_o_4__6_ & pe_o_4__5_;
  assign N4129 = N4128 & N4133;
  assign N4130 = N4129 & pe_o_4__3_;
  assign N4131 = N4130 & N4134;
  assign N4132 = N4131 & pe_o_4__0_;
  assign N8146 = N4132 & N4135;
  assign N4133 = ~pe_o_4__4_;
  assign N4134 = ~pe_o_4__2_;
  assign N4135 = ~pe_o_4__1_;
  assign N4136 = pe_o_4__6_ & pe_o_4__5_;
  assign N4137 = N4136 & N4141;
  assign N4138 = N4137 & pe_o_4__3_;
  assign N4139 = N4138 & N4142;
  assign N4140 = N4139 & N4143;
  assign N8148 = N4140 & pe_o_4__1_;
  assign N4141 = ~pe_o_4__4_;
  assign N4142 = ~pe_o_4__2_;
  assign N4143 = ~pe_o_4__0_;
  assign N4144 = pe_o_4__6_ & pe_o_4__5_;
  assign N4145 = N4144 & N4149;
  assign N4146 = N4145 & pe_o_4__3_;
  assign N4147 = N4146 & N4150;
  assign N4148 = N4147 & pe_o_4__0_;
  assign N8150 = N4148 & pe_o_4__1_;
  assign N4149 = ~pe_o_4__4_;
  assign N4150 = ~pe_o_4__2_;
  assign N4151 = pe_o_4__6_ & pe_o_4__5_;
  assign N4152 = N4151 & N4156;
  assign N4153 = N4152 & pe_o_4__3_;
  assign N4154 = N4153 & pe_o_4__2_;
  assign N4155 = N4154 & N4157;
  assign N8152 = N4155 & N4158;
  assign N4156 = ~pe_o_4__4_;
  assign N4157 = ~pe_o_4__0_;
  assign N4158 = ~pe_o_4__1_;
  assign N4159 = pe_o_4__6_ & pe_o_4__5_;
  assign N4160 = N4159 & N4164;
  assign N4161 = N4160 & pe_o_4__3_;
  assign N4162 = N4161 & pe_o_4__2_;
  assign N4163 = N4162 & pe_o_4__0_;
  assign N8154 = N4163 & N4165;
  assign N4164 = ~pe_o_4__4_;
  assign N4165 = ~pe_o_4__1_;
  assign N4166 = pe_o_4__6_ & pe_o_4__5_;
  assign N4167 = N4166 & N4171;
  assign N4168 = N4167 & pe_o_4__3_;
  assign N4169 = N4168 & pe_o_4__2_;
  assign N4170 = N4169 & N4172;
  assign N8156 = N4170 & pe_o_4__1_;
  assign N4171 = ~pe_o_4__4_;
  assign N4172 = ~pe_o_4__0_;
  assign N4173 = pe_o_4__6_ & pe_o_4__5_;
  assign N4174 = N4173 & pe_o_4__3_;
  assign N4175 = N4174 & pe_o_4__2_;
  assign N4176 = N4175 & pe_o_4__0_;
  assign N8158 = N4176 & pe_o_4__1_;
  assign N4177 = pe_o_4__6_ & pe_o_4__5_;
  assign N4178 = N4177 & pe_o_4__4_;
  assign N4179 = N4178 & N4182;
  assign N4180 = N4179 & N4183;
  assign N4181 = N4180 & N4184;
  assign N8160 = N4181 & N4185;
  assign N4182 = ~pe_o_4__3_;
  assign N4183 = ~pe_o_4__2_;
  assign N4184 = ~pe_o_4__0_;
  assign N4185 = ~pe_o_4__1_;
  assign N4186 = pe_o_4__6_ & pe_o_4__5_;
  assign N4187 = N4186 & pe_o_4__4_;
  assign N4188 = N4187 & N4191;
  assign N4189 = N4188 & N4192;
  assign N4190 = N4189 & pe_o_4__0_;
  assign N8162 = N4190 & N4193;
  assign N4191 = ~pe_o_4__3_;
  assign N4192 = ~pe_o_4__2_;
  assign N4193 = ~pe_o_4__1_;
  assign N4194 = pe_o_4__6_ & pe_o_4__5_;
  assign N4195 = N4194 & pe_o_4__4_;
  assign N4196 = N4195 & N4199;
  assign N4197 = N4196 & N4200;
  assign N4198 = N4197 & N4201;
  assign N8164 = N4198 & pe_o_4__1_;
  assign N4199 = ~pe_o_4__3_;
  assign N4200 = ~pe_o_4__2_;
  assign N4201 = ~pe_o_4__0_;
  assign N4202 = pe_o_4__6_ & pe_o_4__5_;
  assign N4203 = N4202 & pe_o_4__4_;
  assign N4204 = N4203 & N4207;
  assign N4205 = N4204 & N4208;
  assign N4206 = N4205 & pe_o_4__0_;
  assign N8166 = N4206 & pe_o_4__1_;
  assign N4207 = ~pe_o_4__3_;
  assign N4208 = ~pe_o_4__2_;
  assign N4209 = pe_o_4__6_ & pe_o_4__5_;
  assign N4210 = N4209 & pe_o_4__4_;
  assign N4211 = N4210 & N4214;
  assign N4212 = N4211 & pe_o_4__2_;
  assign N4213 = N4212 & N4215;
  assign N8168 = N4213 & N4216;
  assign N4214 = ~pe_o_4__3_;
  assign N4215 = ~pe_o_4__0_;
  assign N4216 = ~pe_o_4__1_;
  assign N4217 = pe_o_4__6_ & pe_o_4__5_;
  assign N4218 = N4217 & pe_o_4__4_;
  assign N4219 = N4218 & N4222;
  assign N4220 = N4219 & pe_o_4__2_;
  assign N4221 = N4220 & pe_o_4__0_;
  assign N8170 = N4221 & N4223;
  assign N4222 = ~pe_o_4__3_;
  assign N4223 = ~pe_o_4__1_;
  assign N4224 = pe_o_4__6_ & pe_o_4__5_;
  assign N4225 = N4224 & pe_o_4__4_;
  assign N4226 = N4225 & N4229;
  assign N4227 = N4226 & pe_o_4__2_;
  assign N4228 = N4227 & N4230;
  assign N8172 = N4228 & pe_o_4__1_;
  assign N4229 = ~pe_o_4__3_;
  assign N4230 = ~pe_o_4__0_;
  assign N4231 = pe_o_4__6_ & pe_o_4__5_;
  assign N4232 = N4231 & pe_o_4__4_;
  assign N4233 = N4232 & pe_o_4__2_;
  assign N4234 = N4233 & pe_o_4__0_;
  assign N8174 = N4234 & pe_o_4__1_;
  assign N4235 = pe_o_4__6_ & pe_o_4__5_;
  assign N4236 = N4235 & pe_o_4__4_;
  assign N4237 = N4236 & pe_o_4__3_;
  assign N4238 = N4237 & N4240;
  assign N4239 = N4238 & N4241;
  assign N8176 = N4239 & N4242;
  assign N4240 = ~pe_o_4__2_;
  assign N4241 = ~pe_o_4__0_;
  assign N4242 = ~pe_o_4__1_;
  assign N4243 = pe_o_4__6_ & pe_o_4__5_;
  assign N4244 = N4243 & pe_o_4__4_;
  assign N4245 = N4244 & pe_o_4__3_;
  assign N4246 = N4245 & N4248;
  assign N4247 = N4246 & pe_o_4__0_;
  assign N8178 = N4247 & N4249;
  assign N4248 = ~pe_o_4__2_;
  assign N4249 = ~pe_o_4__1_;
  assign N4250 = pe_o_4__6_ & pe_o_4__5_;
  assign N4251 = N4250 & pe_o_4__4_;
  assign N4252 = N4251 & pe_o_4__3_;
  assign N4253 = N4252 & N4255;
  assign N4254 = N4253 & N4256;
  assign N8180 = N4254 & pe_o_4__1_;
  assign N4255 = ~pe_o_4__2_;
  assign N4256 = ~pe_o_4__0_;
  assign N4257 = pe_o_4__6_ & pe_o_4__5_;
  assign N4258 = N4257 & pe_o_4__4_;
  assign N4259 = N4258 & pe_o_4__3_;
  assign N4260 = N4259 & pe_o_4__0_;
  assign N8182 = N4260 & pe_o_4__1_;
  assign N4261 = pe_o_4__6_ & pe_o_4__5_;
  assign N4262 = N4261 & pe_o_4__4_;
  assign N4263 = N4262 & pe_o_4__3_;
  assign N4264 = N4263 & pe_o_4__2_;
  assign N4265 = N4264 & N4266;
  assign N8184 = N4265 & N4267;
  assign N4266 = ~pe_o_4__0_;
  assign N4267 = ~pe_o_4__1_;
  assign N4268 = pe_o_4__6_ & pe_o_4__5_;
  assign N4269 = N4268 & pe_o_4__4_;
  assign N4270 = N4269 & pe_o_4__3_;
  assign N4271 = N4270 & pe_o_4__2_;
  assign N8186 = N4271 & pe_o_4__0_;
  assign N4272 = pe_o_4__6_ & pe_o_4__5_;
  assign N4273 = N4272 & pe_o_4__4_;
  assign N4274 = N4273 & pe_o_4__3_;
  assign N4275 = N4274 & pe_o_4__2_;
  assign N8188 = N4275 & pe_o_4__1_;
  assign N4276 = N4281 & N4282;
  assign N4277 = N4276 & N4283;
  assign N4278 = N4277 & N4284;
  assign N4279 = N4278 & N4285;
  assign N4280 = N4279 & N4286;
  assign N8317 = N4280 & N4287;
  assign N4281 = ~pe_o_5__6_;
  assign N4282 = ~pe_o_5__5_;
  assign N4283 = ~pe_o_5__4_;
  assign N4284 = ~pe_o_5__3_;
  assign N4285 = ~pe_o_5__2_;
  assign N4286 = ~pe_o_5__0_;
  assign N4287 = ~pe_o_5__1_;
  assign N4288 = pe_o_5__6_ & N4293;
  assign N4289 = N4288 & N4294;
  assign N4290 = N4289 & N4295;
  assign N4291 = N4290 & N4296;
  assign N4292 = N4291 & N4297;
  assign N8318 = N4292 & N4298;
  assign N4293 = ~pe_o_5__5_;
  assign N4294 = ~pe_o_5__4_;
  assign N4295 = ~pe_o_5__3_;
  assign N4296 = ~pe_o_5__2_;
  assign N4297 = ~pe_o_5__0_;
  assign N4298 = ~pe_o_5__1_;
  assign N4299 = N4304 & N4305;
  assign N4300 = N4299 & N4306;
  assign N4301 = N4300 & N4307;
  assign N4302 = N4301 & N4308;
  assign N4303 = N4302 & pe_o_5__0_;
  assign N8319 = N4303 & N4309;
  assign N4304 = ~pe_o_5__6_;
  assign N4305 = ~pe_o_5__5_;
  assign N4306 = ~pe_o_5__4_;
  assign N4307 = ~pe_o_5__3_;
  assign N4308 = ~pe_o_5__2_;
  assign N4309 = ~pe_o_5__1_;
  assign N4310 = N4315 & N4316;
  assign N4311 = N4310 & N4317;
  assign N4312 = N4311 & N4318;
  assign N4313 = N4312 & N4319;
  assign N4314 = N4313 & N4320;
  assign N8321 = N4314 & pe_o_5__1_;
  assign N4315 = ~pe_o_5__6_;
  assign N4316 = ~pe_o_5__5_;
  assign N4317 = ~pe_o_5__4_;
  assign N4318 = ~pe_o_5__3_;
  assign N4319 = ~pe_o_5__2_;
  assign N4320 = ~pe_o_5__0_;
  assign N4321 = N4326 & N4327;
  assign N4322 = N4321 & N4328;
  assign N4323 = N4322 & N4329;
  assign N4324 = N4323 & N4330;
  assign N4325 = N4324 & pe_o_5__0_;
  assign N8323 = N4325 & pe_o_5__1_;
  assign N4326 = ~pe_o_5__6_;
  assign N4327 = ~pe_o_5__5_;
  assign N4328 = ~pe_o_5__4_;
  assign N4329 = ~pe_o_5__3_;
  assign N4330 = ~pe_o_5__2_;
  assign N4331 = N4336 & N4337;
  assign N4332 = N4331 & N4338;
  assign N4333 = N4332 & N4339;
  assign N4334 = N4333 & pe_o_5__2_;
  assign N4335 = N4334 & N4340;
  assign N8325 = N4335 & N4341;
  assign N4336 = ~pe_o_5__6_;
  assign N4337 = ~pe_o_5__5_;
  assign N4338 = ~pe_o_5__4_;
  assign N4339 = ~pe_o_5__3_;
  assign N4340 = ~pe_o_5__0_;
  assign N4341 = ~pe_o_5__1_;
  assign N4342 = N4347 & N4348;
  assign N4343 = N4342 & N4349;
  assign N4344 = N4343 & N4350;
  assign N4345 = N4344 & pe_o_5__2_;
  assign N4346 = N4345 & pe_o_5__0_;
  assign N8327 = N4346 & N4351;
  assign N4347 = ~pe_o_5__6_;
  assign N4348 = ~pe_o_5__5_;
  assign N4349 = ~pe_o_5__4_;
  assign N4350 = ~pe_o_5__3_;
  assign N4351 = ~pe_o_5__1_;
  assign N4352 = N4357 & N4358;
  assign N4353 = N4352 & N4359;
  assign N4354 = N4353 & N4360;
  assign N4355 = N4354 & pe_o_5__2_;
  assign N4356 = N4355 & N4361;
  assign N8329 = N4356 & pe_o_5__1_;
  assign N4357 = ~pe_o_5__6_;
  assign N4358 = ~pe_o_5__5_;
  assign N4359 = ~pe_o_5__4_;
  assign N4360 = ~pe_o_5__3_;
  assign N4361 = ~pe_o_5__0_;
  assign N4362 = N4367 & N4368;
  assign N4363 = N4362 & N4369;
  assign N4364 = N4363 & N4370;
  assign N4365 = N4364 & pe_o_5__2_;
  assign N4366 = N4365 & pe_o_5__0_;
  assign N8331 = N4366 & pe_o_5__1_;
  assign N4367 = ~pe_o_5__6_;
  assign N4368 = ~pe_o_5__5_;
  assign N4369 = ~pe_o_5__4_;
  assign N4370 = ~pe_o_5__3_;
  assign N4371 = N4376 & N4377;
  assign N4372 = N4371 & N4378;
  assign N4373 = N4372 & pe_o_5__3_;
  assign N4374 = N4373 & N4379;
  assign N4375 = N4374 & N4380;
  assign N8333 = N4375 & N4381;
  assign N4376 = ~pe_o_5__6_;
  assign N4377 = ~pe_o_5__5_;
  assign N4378 = ~pe_o_5__4_;
  assign N4379 = ~pe_o_5__2_;
  assign N4380 = ~pe_o_5__0_;
  assign N4381 = ~pe_o_5__1_;
  assign N4382 = N4387 & N4388;
  assign N4383 = N4382 & N4389;
  assign N4384 = N4383 & pe_o_5__3_;
  assign N4385 = N4384 & N4390;
  assign N4386 = N4385 & pe_o_5__0_;
  assign N8335 = N4386 & N4391;
  assign N4387 = ~pe_o_5__6_;
  assign N4388 = ~pe_o_5__5_;
  assign N4389 = ~pe_o_5__4_;
  assign N4390 = ~pe_o_5__2_;
  assign N4391 = ~pe_o_5__1_;
  assign N4392 = N4397 & N4398;
  assign N4393 = N4392 & N4399;
  assign N4394 = N4393 & pe_o_5__3_;
  assign N4395 = N4394 & N4400;
  assign N4396 = N4395 & N4401;
  assign N8337 = N4396 & pe_o_5__1_;
  assign N4397 = ~pe_o_5__6_;
  assign N4398 = ~pe_o_5__5_;
  assign N4399 = ~pe_o_5__4_;
  assign N4400 = ~pe_o_5__2_;
  assign N4401 = ~pe_o_5__0_;
  assign N4402 = N4407 & N4408;
  assign N4403 = N4402 & N4409;
  assign N4404 = N4403 & pe_o_5__3_;
  assign N4405 = N4404 & N4410;
  assign N4406 = N4405 & pe_o_5__0_;
  assign N8339 = N4406 & pe_o_5__1_;
  assign N4407 = ~pe_o_5__6_;
  assign N4408 = ~pe_o_5__5_;
  assign N4409 = ~pe_o_5__4_;
  assign N4410 = ~pe_o_5__2_;
  assign N4411 = N4416 & N4417;
  assign N4412 = N4411 & N4418;
  assign N4413 = N4412 & pe_o_5__3_;
  assign N4414 = N4413 & pe_o_5__2_;
  assign N4415 = N4414 & N4419;
  assign N8341 = N4415 & N4420;
  assign N4416 = ~pe_o_5__6_;
  assign N4417 = ~pe_o_5__5_;
  assign N4418 = ~pe_o_5__4_;
  assign N4419 = ~pe_o_5__0_;
  assign N4420 = ~pe_o_5__1_;
  assign N4421 = N4426 & N4427;
  assign N4422 = N4421 & N4428;
  assign N4423 = N4422 & pe_o_5__3_;
  assign N4424 = N4423 & pe_o_5__2_;
  assign N4425 = N4424 & pe_o_5__0_;
  assign N8343 = N4425 & N4429;
  assign N4426 = ~pe_o_5__6_;
  assign N4427 = ~pe_o_5__5_;
  assign N4428 = ~pe_o_5__4_;
  assign N4429 = ~pe_o_5__1_;
  assign N4430 = N4435 & N4436;
  assign N4431 = N4430 & N4437;
  assign N4432 = N4431 & pe_o_5__3_;
  assign N4433 = N4432 & pe_o_5__2_;
  assign N4434 = N4433 & N4438;
  assign N8345 = N4434 & pe_o_5__1_;
  assign N4435 = ~pe_o_5__6_;
  assign N4436 = ~pe_o_5__5_;
  assign N4437 = ~pe_o_5__4_;
  assign N4438 = ~pe_o_5__0_;
  assign N4439 = N4444 & N4445;
  assign N4440 = N4439 & N4446;
  assign N4441 = N4440 & pe_o_5__3_;
  assign N4442 = N4441 & pe_o_5__2_;
  assign N4443 = N4442 & pe_o_5__0_;
  assign N8347 = N4443 & pe_o_5__1_;
  assign N4444 = ~pe_o_5__6_;
  assign N4445 = ~pe_o_5__5_;
  assign N4446 = ~pe_o_5__4_;
  assign N4447 = N4452 & N4453;
  assign N4448 = N4447 & pe_o_5__4_;
  assign N4449 = N4448 & N4454;
  assign N4450 = N4449 & N4455;
  assign N4451 = N4450 & N4456;
  assign N8349 = N4451 & N4457;
  assign N4452 = ~pe_o_5__6_;
  assign N4453 = ~pe_o_5__5_;
  assign N4454 = ~pe_o_5__3_;
  assign N4455 = ~pe_o_5__2_;
  assign N4456 = ~pe_o_5__0_;
  assign N4457 = ~pe_o_5__1_;
  assign N4458 = N4463 & N4464;
  assign N4459 = N4458 & pe_o_5__4_;
  assign N4460 = N4459 & N4465;
  assign N4461 = N4460 & N4466;
  assign N4462 = N4461 & pe_o_5__0_;
  assign N8351 = N4462 & N4467;
  assign N4463 = ~pe_o_5__6_;
  assign N4464 = ~pe_o_5__5_;
  assign N4465 = ~pe_o_5__3_;
  assign N4466 = ~pe_o_5__2_;
  assign N4467 = ~pe_o_5__1_;
  assign N4468 = N4473 & N4474;
  assign N4469 = N4468 & pe_o_5__4_;
  assign N4470 = N4469 & N4475;
  assign N4471 = N4470 & N4476;
  assign N4472 = N4471 & N4477;
  assign N8353 = N4472 & pe_o_5__1_;
  assign N4473 = ~pe_o_5__6_;
  assign N4474 = ~pe_o_5__5_;
  assign N4475 = ~pe_o_5__3_;
  assign N4476 = ~pe_o_5__2_;
  assign N4477 = ~pe_o_5__0_;
  assign N4478 = N4483 & N4484;
  assign N4479 = N4478 & pe_o_5__4_;
  assign N4480 = N4479 & N4485;
  assign N4481 = N4480 & N4486;
  assign N4482 = N4481 & pe_o_5__0_;
  assign N8355 = N4482 & pe_o_5__1_;
  assign N4483 = ~pe_o_5__6_;
  assign N4484 = ~pe_o_5__5_;
  assign N4485 = ~pe_o_5__3_;
  assign N4486 = ~pe_o_5__2_;
  assign N4487 = N4492 & N4493;
  assign N4488 = N4487 & pe_o_5__4_;
  assign N4489 = N4488 & N4494;
  assign N4490 = N4489 & pe_o_5__2_;
  assign N4491 = N4490 & N4495;
  assign N8357 = N4491 & N4496;
  assign N4492 = ~pe_o_5__6_;
  assign N4493 = ~pe_o_5__5_;
  assign N4494 = ~pe_o_5__3_;
  assign N4495 = ~pe_o_5__0_;
  assign N4496 = ~pe_o_5__1_;
  assign N4497 = N4502 & N4503;
  assign N4498 = N4497 & pe_o_5__4_;
  assign N4499 = N4498 & N4504;
  assign N4500 = N4499 & pe_o_5__2_;
  assign N4501 = N4500 & pe_o_5__0_;
  assign N8359 = N4501 & N4505;
  assign N4502 = ~pe_o_5__6_;
  assign N4503 = ~pe_o_5__5_;
  assign N4504 = ~pe_o_5__3_;
  assign N4505 = ~pe_o_5__1_;
  assign N4506 = N4511 & N4512;
  assign N4507 = N4506 & pe_o_5__4_;
  assign N4508 = N4507 & N4513;
  assign N4509 = N4508 & pe_o_5__2_;
  assign N4510 = N4509 & N4514;
  assign N8361 = N4510 & pe_o_5__1_;
  assign N4511 = ~pe_o_5__6_;
  assign N4512 = ~pe_o_5__5_;
  assign N4513 = ~pe_o_5__3_;
  assign N4514 = ~pe_o_5__0_;
  assign N4515 = N4520 & N4521;
  assign N4516 = N4515 & pe_o_5__4_;
  assign N4517 = N4516 & N4522;
  assign N4518 = N4517 & pe_o_5__2_;
  assign N4519 = N4518 & pe_o_5__0_;
  assign N8363 = N4519 & pe_o_5__1_;
  assign N4520 = ~pe_o_5__6_;
  assign N4521 = ~pe_o_5__5_;
  assign N4522 = ~pe_o_5__3_;
  assign N4523 = N4528 & N4529;
  assign N4524 = N4523 & pe_o_5__4_;
  assign N4525 = N4524 & pe_o_5__3_;
  assign N4526 = N4525 & N4530;
  assign N4527 = N4526 & N4531;
  assign N8365 = N4527 & N4532;
  assign N4528 = ~pe_o_5__6_;
  assign N4529 = ~pe_o_5__5_;
  assign N4530 = ~pe_o_5__2_;
  assign N4531 = ~pe_o_5__0_;
  assign N4532 = ~pe_o_5__1_;
  assign N4533 = N4538 & N4539;
  assign N4534 = N4533 & pe_o_5__4_;
  assign N4535 = N4534 & pe_o_5__3_;
  assign N4536 = N4535 & N4540;
  assign N4537 = N4536 & pe_o_5__0_;
  assign N8367 = N4537 & N4541;
  assign N4538 = ~pe_o_5__6_;
  assign N4539 = ~pe_o_5__5_;
  assign N4540 = ~pe_o_5__2_;
  assign N4541 = ~pe_o_5__1_;
  assign N4542 = N4547 & N4548;
  assign N4543 = N4542 & pe_o_5__4_;
  assign N4544 = N4543 & pe_o_5__3_;
  assign N4545 = N4544 & N4549;
  assign N4546 = N4545 & N4550;
  assign N8369 = N4546 & pe_o_5__1_;
  assign N4547 = ~pe_o_5__6_;
  assign N4548 = ~pe_o_5__5_;
  assign N4549 = ~pe_o_5__2_;
  assign N4550 = ~pe_o_5__0_;
  assign N4551 = N4556 & N4557;
  assign N4552 = N4551 & pe_o_5__4_;
  assign N4553 = N4552 & pe_o_5__3_;
  assign N4554 = N4553 & N4558;
  assign N4555 = N4554 & pe_o_5__0_;
  assign N8371 = N4555 & pe_o_5__1_;
  assign N4556 = ~pe_o_5__6_;
  assign N4557 = ~pe_o_5__5_;
  assign N4558 = ~pe_o_5__2_;
  assign N4559 = N4564 & N4565;
  assign N4560 = N4559 & pe_o_5__4_;
  assign N4561 = N4560 & pe_o_5__3_;
  assign N4562 = N4561 & pe_o_5__2_;
  assign N4563 = N4562 & N4566;
  assign N8373 = N4563 & N4567;
  assign N4564 = ~pe_o_5__6_;
  assign N4565 = ~pe_o_5__5_;
  assign N4566 = ~pe_o_5__0_;
  assign N4567 = ~pe_o_5__1_;
  assign N4568 = N4573 & N4574;
  assign N4569 = N4568 & pe_o_5__4_;
  assign N4570 = N4569 & pe_o_5__3_;
  assign N4571 = N4570 & pe_o_5__2_;
  assign N4572 = N4571 & pe_o_5__0_;
  assign N8375 = N4572 & N4575;
  assign N4573 = ~pe_o_5__6_;
  assign N4574 = ~pe_o_5__5_;
  assign N4575 = ~pe_o_5__1_;
  assign N4576 = N4581 & N4582;
  assign N4577 = N4576 & pe_o_5__4_;
  assign N4578 = N4577 & pe_o_5__3_;
  assign N4579 = N4578 & pe_o_5__2_;
  assign N4580 = N4579 & N4583;
  assign N8377 = N4580 & pe_o_5__1_;
  assign N4581 = ~pe_o_5__6_;
  assign N4582 = ~pe_o_5__5_;
  assign N4583 = ~pe_o_5__0_;
  assign N4584 = N4589 & N4590;
  assign N4585 = N4584 & pe_o_5__4_;
  assign N4586 = N4585 & pe_o_5__3_;
  assign N4587 = N4586 & pe_o_5__2_;
  assign N4588 = N4587 & pe_o_5__0_;
  assign N8379 = N4588 & pe_o_5__1_;
  assign N4589 = ~pe_o_5__6_;
  assign N4590 = ~pe_o_5__5_;
  assign N4591 = N4596 & pe_o_5__5_;
  assign N4592 = N4591 & N4597;
  assign N4593 = N4592 & N4598;
  assign N4594 = N4593 & N4599;
  assign N4595 = N4594 & N4600;
  assign N8381 = N4595 & N4601;
  assign N4596 = ~pe_o_5__6_;
  assign N4597 = ~pe_o_5__4_;
  assign N4598 = ~pe_o_5__3_;
  assign N4599 = ~pe_o_5__2_;
  assign N4600 = ~pe_o_5__0_;
  assign N4601 = ~pe_o_5__1_;
  assign N4602 = N4607 & pe_o_5__5_;
  assign N4603 = N4602 & N4608;
  assign N4604 = N4603 & N4609;
  assign N4605 = N4604 & N4610;
  assign N4606 = N4605 & pe_o_5__0_;
  assign N8383 = N4606 & N4611;
  assign N4607 = ~pe_o_5__6_;
  assign N4608 = ~pe_o_5__4_;
  assign N4609 = ~pe_o_5__3_;
  assign N4610 = ~pe_o_5__2_;
  assign N4611 = ~pe_o_5__1_;
  assign N4612 = N4617 & pe_o_5__5_;
  assign N4613 = N4612 & N4618;
  assign N4614 = N4613 & N4619;
  assign N4615 = N4614 & N4620;
  assign N4616 = N4615 & N4621;
  assign N8385 = N4616 & pe_o_5__1_;
  assign N4617 = ~pe_o_5__6_;
  assign N4618 = ~pe_o_5__4_;
  assign N4619 = ~pe_o_5__3_;
  assign N4620 = ~pe_o_5__2_;
  assign N4621 = ~pe_o_5__0_;
  assign N4622 = N4627 & pe_o_5__5_;
  assign N4623 = N4622 & N4628;
  assign N4624 = N4623 & N4629;
  assign N4625 = N4624 & N4630;
  assign N4626 = N4625 & pe_o_5__0_;
  assign N8387 = N4626 & pe_o_5__1_;
  assign N4627 = ~pe_o_5__6_;
  assign N4628 = ~pe_o_5__4_;
  assign N4629 = ~pe_o_5__3_;
  assign N4630 = ~pe_o_5__2_;
  assign N4631 = N4636 & pe_o_5__5_;
  assign N4632 = N4631 & N4637;
  assign N4633 = N4632 & N4638;
  assign N4634 = N4633 & pe_o_5__2_;
  assign N4635 = N4634 & N4639;
  assign N8389 = N4635 & N4640;
  assign N4636 = ~pe_o_5__6_;
  assign N4637 = ~pe_o_5__4_;
  assign N4638 = ~pe_o_5__3_;
  assign N4639 = ~pe_o_5__0_;
  assign N4640 = ~pe_o_5__1_;
  assign N4641 = N4646 & pe_o_5__5_;
  assign N4642 = N4641 & N4647;
  assign N4643 = N4642 & N4648;
  assign N4644 = N4643 & pe_o_5__2_;
  assign N4645 = N4644 & pe_o_5__0_;
  assign N8391 = N4645 & N4649;
  assign N4646 = ~pe_o_5__6_;
  assign N4647 = ~pe_o_5__4_;
  assign N4648 = ~pe_o_5__3_;
  assign N4649 = ~pe_o_5__1_;
  assign N4650 = N4655 & pe_o_5__5_;
  assign N4651 = N4650 & N4656;
  assign N4652 = N4651 & N4657;
  assign N4653 = N4652 & pe_o_5__2_;
  assign N4654 = N4653 & N4658;
  assign N8393 = N4654 & pe_o_5__1_;
  assign N4655 = ~pe_o_5__6_;
  assign N4656 = ~pe_o_5__4_;
  assign N4657 = ~pe_o_5__3_;
  assign N4658 = ~pe_o_5__0_;
  assign N4659 = N4664 & pe_o_5__5_;
  assign N4660 = N4659 & N4665;
  assign N4661 = N4660 & N4666;
  assign N4662 = N4661 & pe_o_5__2_;
  assign N4663 = N4662 & pe_o_5__0_;
  assign N8395 = N4663 & pe_o_5__1_;
  assign N4664 = ~pe_o_5__6_;
  assign N4665 = ~pe_o_5__4_;
  assign N4666 = ~pe_o_5__3_;
  assign N4667 = N4672 & pe_o_5__5_;
  assign N4668 = N4667 & N4673;
  assign N4669 = N4668 & pe_o_5__3_;
  assign N4670 = N4669 & N4674;
  assign N4671 = N4670 & N4675;
  assign N8397 = N4671 & N4676;
  assign N4672 = ~pe_o_5__6_;
  assign N4673 = ~pe_o_5__4_;
  assign N4674 = ~pe_o_5__2_;
  assign N4675 = ~pe_o_5__0_;
  assign N4676 = ~pe_o_5__1_;
  assign N4677 = N4682 & pe_o_5__5_;
  assign N4678 = N4677 & N4683;
  assign N4679 = N4678 & pe_o_5__3_;
  assign N4680 = N4679 & N4684;
  assign N4681 = N4680 & pe_o_5__0_;
  assign N8399 = N4681 & N4685;
  assign N4682 = ~pe_o_5__6_;
  assign N4683 = ~pe_o_5__4_;
  assign N4684 = ~pe_o_5__2_;
  assign N4685 = ~pe_o_5__1_;
  assign N4686 = N4691 & pe_o_5__5_;
  assign N4687 = N4686 & N4692;
  assign N4688 = N4687 & pe_o_5__3_;
  assign N4689 = N4688 & N4693;
  assign N4690 = N4689 & N4694;
  assign N8401 = N4690 & pe_o_5__1_;
  assign N4691 = ~pe_o_5__6_;
  assign N4692 = ~pe_o_5__4_;
  assign N4693 = ~pe_o_5__2_;
  assign N4694 = ~pe_o_5__0_;
  assign N4695 = N4700 & pe_o_5__5_;
  assign N4696 = N4695 & N4701;
  assign N4697 = N4696 & pe_o_5__3_;
  assign N4698 = N4697 & N4702;
  assign N4699 = N4698 & pe_o_5__0_;
  assign N8403 = N4699 & pe_o_5__1_;
  assign N4700 = ~pe_o_5__6_;
  assign N4701 = ~pe_o_5__4_;
  assign N4702 = ~pe_o_5__2_;
  assign N4703 = N4708 & pe_o_5__5_;
  assign N4704 = N4703 & N4709;
  assign N4705 = N4704 & pe_o_5__3_;
  assign N4706 = N4705 & pe_o_5__2_;
  assign N4707 = N4706 & N4710;
  assign N8405 = N4707 & N4711;
  assign N4708 = ~pe_o_5__6_;
  assign N4709 = ~pe_o_5__4_;
  assign N4710 = ~pe_o_5__0_;
  assign N4711 = ~pe_o_5__1_;
  assign N4712 = N4717 & pe_o_5__5_;
  assign N4713 = N4712 & N4718;
  assign N4714 = N4713 & pe_o_5__3_;
  assign N4715 = N4714 & pe_o_5__2_;
  assign N4716 = N4715 & pe_o_5__0_;
  assign N8407 = N4716 & N4719;
  assign N4717 = ~pe_o_5__6_;
  assign N4718 = ~pe_o_5__4_;
  assign N4719 = ~pe_o_5__1_;
  assign N4720 = N4725 & pe_o_5__5_;
  assign N4721 = N4720 & N4726;
  assign N4722 = N4721 & pe_o_5__3_;
  assign N4723 = N4722 & pe_o_5__2_;
  assign N4724 = N4723 & N4727;
  assign N8409 = N4724 & pe_o_5__1_;
  assign N4725 = ~pe_o_5__6_;
  assign N4726 = ~pe_o_5__4_;
  assign N4727 = ~pe_o_5__0_;
  assign N4728 = N4733 & pe_o_5__5_;
  assign N4729 = N4728 & N4734;
  assign N4730 = N4729 & pe_o_5__3_;
  assign N4731 = N4730 & pe_o_5__2_;
  assign N4732 = N4731 & pe_o_5__0_;
  assign N8411 = N4732 & pe_o_5__1_;
  assign N4733 = ~pe_o_5__6_;
  assign N4734 = ~pe_o_5__4_;
  assign N4735 = N4740 & pe_o_5__5_;
  assign N4736 = N4735 & pe_o_5__4_;
  assign N4737 = N4736 & N4741;
  assign N4738 = N4737 & N4742;
  assign N4739 = N4738 & N4743;
  assign N8413 = N4739 & N4744;
  assign N4740 = ~pe_o_5__6_;
  assign N4741 = ~pe_o_5__3_;
  assign N4742 = ~pe_o_5__2_;
  assign N4743 = ~pe_o_5__0_;
  assign N4744 = ~pe_o_5__1_;
  assign N4745 = N4750 & pe_o_5__5_;
  assign N4746 = N4745 & pe_o_5__4_;
  assign N4747 = N4746 & N4751;
  assign N4748 = N4747 & N4752;
  assign N4749 = N4748 & pe_o_5__0_;
  assign N8415 = N4749 & N4753;
  assign N4750 = ~pe_o_5__6_;
  assign N4751 = ~pe_o_5__3_;
  assign N4752 = ~pe_o_5__2_;
  assign N4753 = ~pe_o_5__1_;
  assign N4754 = N4759 & pe_o_5__5_;
  assign N4755 = N4754 & pe_o_5__4_;
  assign N4756 = N4755 & N4760;
  assign N4757 = N4756 & N4761;
  assign N4758 = N4757 & N4762;
  assign N8417 = N4758 & pe_o_5__1_;
  assign N4759 = ~pe_o_5__6_;
  assign N4760 = ~pe_o_5__3_;
  assign N4761 = ~pe_o_5__2_;
  assign N4762 = ~pe_o_5__0_;
  assign N4763 = N4768 & pe_o_5__5_;
  assign N4764 = N4763 & pe_o_5__4_;
  assign N4765 = N4764 & N4769;
  assign N4766 = N4765 & N4770;
  assign N4767 = N4766 & pe_o_5__0_;
  assign N8419 = N4767 & pe_o_5__1_;
  assign N4768 = ~pe_o_5__6_;
  assign N4769 = ~pe_o_5__3_;
  assign N4770 = ~pe_o_5__2_;
  assign N4771 = N4776 & pe_o_5__5_;
  assign N4772 = N4771 & pe_o_5__4_;
  assign N4773 = N4772 & N4777;
  assign N4774 = N4773 & pe_o_5__2_;
  assign N4775 = N4774 & N4778;
  assign N8421 = N4775 & N4779;
  assign N4776 = ~pe_o_5__6_;
  assign N4777 = ~pe_o_5__3_;
  assign N4778 = ~pe_o_5__0_;
  assign N4779 = ~pe_o_5__1_;
  assign N4780 = N4785 & pe_o_5__5_;
  assign N4781 = N4780 & pe_o_5__4_;
  assign N4782 = N4781 & N4786;
  assign N4783 = N4782 & pe_o_5__2_;
  assign N4784 = N4783 & pe_o_5__0_;
  assign N8423 = N4784 & N4787;
  assign N4785 = ~pe_o_5__6_;
  assign N4786 = ~pe_o_5__3_;
  assign N4787 = ~pe_o_5__1_;
  assign N4788 = N4793 & pe_o_5__5_;
  assign N4789 = N4788 & pe_o_5__4_;
  assign N4790 = N4789 & N4794;
  assign N4791 = N4790 & pe_o_5__2_;
  assign N4792 = N4791 & N4795;
  assign N8425 = N4792 & pe_o_5__1_;
  assign N4793 = ~pe_o_5__6_;
  assign N4794 = ~pe_o_5__3_;
  assign N4795 = ~pe_o_5__0_;
  assign N4796 = N4801 & pe_o_5__5_;
  assign N4797 = N4796 & pe_o_5__4_;
  assign N4798 = N4797 & N4802;
  assign N4799 = N4798 & pe_o_5__2_;
  assign N4800 = N4799 & pe_o_5__0_;
  assign N8427 = N4800 & pe_o_5__1_;
  assign N4801 = ~pe_o_5__6_;
  assign N4802 = ~pe_o_5__3_;
  assign N4803 = N4808 & pe_o_5__5_;
  assign N4804 = N4803 & pe_o_5__4_;
  assign N4805 = N4804 & pe_o_5__3_;
  assign N4806 = N4805 & N4809;
  assign N4807 = N4806 & N4810;
  assign N8429 = N4807 & N4811;
  assign N4808 = ~pe_o_5__6_;
  assign N4809 = ~pe_o_5__2_;
  assign N4810 = ~pe_o_5__0_;
  assign N4811 = ~pe_o_5__1_;
  assign N4812 = N4817 & pe_o_5__5_;
  assign N4813 = N4812 & pe_o_5__4_;
  assign N4814 = N4813 & pe_o_5__3_;
  assign N4815 = N4814 & N4818;
  assign N4816 = N4815 & pe_o_5__0_;
  assign N8431 = N4816 & N4819;
  assign N4817 = ~pe_o_5__6_;
  assign N4818 = ~pe_o_5__2_;
  assign N4819 = ~pe_o_5__1_;
  assign N4820 = N4825 & pe_o_5__5_;
  assign N4821 = N4820 & pe_o_5__4_;
  assign N4822 = N4821 & pe_o_5__3_;
  assign N4823 = N4822 & N4826;
  assign N4824 = N4823 & N4827;
  assign N8433 = N4824 & pe_o_5__1_;
  assign N4825 = ~pe_o_5__6_;
  assign N4826 = ~pe_o_5__2_;
  assign N4827 = ~pe_o_5__0_;
  assign N4828 = N4833 & pe_o_5__5_;
  assign N4829 = N4828 & pe_o_5__4_;
  assign N4830 = N4829 & pe_o_5__3_;
  assign N4831 = N4830 & N4834;
  assign N4832 = N4831 & pe_o_5__0_;
  assign N8435 = N4832 & pe_o_5__1_;
  assign N4833 = ~pe_o_5__6_;
  assign N4834 = ~pe_o_5__2_;
  assign N4835 = N4840 & pe_o_5__5_;
  assign N4836 = N4835 & pe_o_5__4_;
  assign N4837 = N4836 & pe_o_5__3_;
  assign N4838 = N4837 & pe_o_5__2_;
  assign N4839 = N4838 & N4841;
  assign N8437 = N4839 & N4842;
  assign N4840 = ~pe_o_5__6_;
  assign N4841 = ~pe_o_5__0_;
  assign N4842 = ~pe_o_5__1_;
  assign N4843 = N4848 & pe_o_5__5_;
  assign N4844 = N4843 & pe_o_5__4_;
  assign N4845 = N4844 & pe_o_5__3_;
  assign N4846 = N4845 & pe_o_5__2_;
  assign N4847 = N4846 & pe_o_5__0_;
  assign N8439 = N4847 & N4849;
  assign N4848 = ~pe_o_5__6_;
  assign N4849 = ~pe_o_5__1_;
  assign N4850 = N4855 & pe_o_5__5_;
  assign N4851 = N4850 & pe_o_5__4_;
  assign N4852 = N4851 & pe_o_5__3_;
  assign N4853 = N4852 & pe_o_5__2_;
  assign N4854 = N4853 & N4856;
  assign N8441 = N4854 & pe_o_5__1_;
  assign N4855 = ~pe_o_5__6_;
  assign N4856 = ~pe_o_5__0_;
  assign N4857 = pe_o_5__5_ & pe_o_5__4_;
  assign N4858 = N4857 & pe_o_5__3_;
  assign N4859 = N4858 & pe_o_5__2_;
  assign N4860 = N4859 & pe_o_5__0_;
  assign N8443 = N4860 & pe_o_5__1_;
  assign N4861 = pe_o_5__6_ & N4866;
  assign N4862 = N4861 & N4867;
  assign N4863 = N4862 & N4868;
  assign N4864 = N4863 & N4869;
  assign N4865 = N4864 & pe_o_5__0_;
  assign N8320 = N4865 & N4870;
  assign N4866 = ~pe_o_5__5_;
  assign N4867 = ~pe_o_5__4_;
  assign N4868 = ~pe_o_5__3_;
  assign N4869 = ~pe_o_5__2_;
  assign N4870 = ~pe_o_5__1_;
  assign N4871 = pe_o_5__6_ & N4876;
  assign N4872 = N4871 & N4877;
  assign N4873 = N4872 & N4878;
  assign N4874 = N4873 & N4879;
  assign N4875 = N4874 & N4880;
  assign N8322 = N4875 & pe_o_5__1_;
  assign N4876 = ~pe_o_5__5_;
  assign N4877 = ~pe_o_5__4_;
  assign N4878 = ~pe_o_5__3_;
  assign N4879 = ~pe_o_5__2_;
  assign N4880 = ~pe_o_5__0_;
  assign N4881 = pe_o_5__6_ & N4886;
  assign N4882 = N4881 & N4887;
  assign N4883 = N4882 & N4888;
  assign N4884 = N4883 & N4889;
  assign N4885 = N4884 & pe_o_5__0_;
  assign N8324 = N4885 & pe_o_5__1_;
  assign N4886 = ~pe_o_5__5_;
  assign N4887 = ~pe_o_5__4_;
  assign N4888 = ~pe_o_5__3_;
  assign N4889 = ~pe_o_5__2_;
  assign N4890 = pe_o_5__6_ & N4895;
  assign N4891 = N4890 & N4896;
  assign N4892 = N4891 & N4897;
  assign N4893 = N4892 & pe_o_5__2_;
  assign N4894 = N4893 & N4898;
  assign N8326 = N4894 & N4899;
  assign N4895 = ~pe_o_5__5_;
  assign N4896 = ~pe_o_5__4_;
  assign N4897 = ~pe_o_5__3_;
  assign N4898 = ~pe_o_5__0_;
  assign N4899 = ~pe_o_5__1_;
  assign N4900 = pe_o_5__6_ & N4905;
  assign N4901 = N4900 & N4906;
  assign N4902 = N4901 & N4907;
  assign N4903 = N4902 & pe_o_5__2_;
  assign N4904 = N4903 & pe_o_5__0_;
  assign N8328 = N4904 & N4908;
  assign N4905 = ~pe_o_5__5_;
  assign N4906 = ~pe_o_5__4_;
  assign N4907 = ~pe_o_5__3_;
  assign N4908 = ~pe_o_5__1_;
  assign N4909 = pe_o_5__6_ & N4914;
  assign N4910 = N4909 & N4915;
  assign N4911 = N4910 & N4916;
  assign N4912 = N4911 & pe_o_5__2_;
  assign N4913 = N4912 & N4917;
  assign N8330 = N4913 & pe_o_5__1_;
  assign N4914 = ~pe_o_5__5_;
  assign N4915 = ~pe_o_5__4_;
  assign N4916 = ~pe_o_5__3_;
  assign N4917 = ~pe_o_5__0_;
  assign N4918 = pe_o_5__6_ & N4923;
  assign N4919 = N4918 & N4924;
  assign N4920 = N4919 & N4925;
  assign N4921 = N4920 & pe_o_5__2_;
  assign N4922 = N4921 & pe_o_5__0_;
  assign N8332 = N4922 & pe_o_5__1_;
  assign N4923 = ~pe_o_5__5_;
  assign N4924 = ~pe_o_5__4_;
  assign N4925 = ~pe_o_5__3_;
  assign N4926 = pe_o_5__6_ & N4931;
  assign N4927 = N4926 & N4932;
  assign N4928 = N4927 & pe_o_5__3_;
  assign N4929 = N4928 & N4933;
  assign N4930 = N4929 & N4934;
  assign N8334 = N4930 & N4935;
  assign N4931 = ~pe_o_5__5_;
  assign N4932 = ~pe_o_5__4_;
  assign N4933 = ~pe_o_5__2_;
  assign N4934 = ~pe_o_5__0_;
  assign N4935 = ~pe_o_5__1_;
  assign N4936 = pe_o_5__6_ & N4941;
  assign N4937 = N4936 & N4942;
  assign N4938 = N4937 & pe_o_5__3_;
  assign N4939 = N4938 & N4943;
  assign N4940 = N4939 & pe_o_5__0_;
  assign N8336 = N4940 & N4944;
  assign N4941 = ~pe_o_5__5_;
  assign N4942 = ~pe_o_5__4_;
  assign N4943 = ~pe_o_5__2_;
  assign N4944 = ~pe_o_5__1_;
  assign N4945 = pe_o_5__6_ & N4950;
  assign N4946 = N4945 & N4951;
  assign N4947 = N4946 & pe_o_5__3_;
  assign N4948 = N4947 & N4952;
  assign N4949 = N4948 & N4953;
  assign N8338 = N4949 & pe_o_5__1_;
  assign N4950 = ~pe_o_5__5_;
  assign N4951 = ~pe_o_5__4_;
  assign N4952 = ~pe_o_5__2_;
  assign N4953 = ~pe_o_5__0_;
  assign N4954 = pe_o_5__6_ & N4959;
  assign N4955 = N4954 & N4960;
  assign N4956 = N4955 & pe_o_5__3_;
  assign N4957 = N4956 & N4961;
  assign N4958 = N4957 & pe_o_5__0_;
  assign N8340 = N4958 & pe_o_5__1_;
  assign N4959 = ~pe_o_5__5_;
  assign N4960 = ~pe_o_5__4_;
  assign N4961 = ~pe_o_5__2_;
  assign N4962 = pe_o_5__6_ & N4967;
  assign N4963 = N4962 & N4968;
  assign N4964 = N4963 & pe_o_5__3_;
  assign N4965 = N4964 & pe_o_5__2_;
  assign N4966 = N4965 & N4969;
  assign N8342 = N4966 & N4970;
  assign N4967 = ~pe_o_5__5_;
  assign N4968 = ~pe_o_5__4_;
  assign N4969 = ~pe_o_5__0_;
  assign N4970 = ~pe_o_5__1_;
  assign N4971 = pe_o_5__6_ & N4976;
  assign N4972 = N4971 & N4977;
  assign N4973 = N4972 & pe_o_5__3_;
  assign N4974 = N4973 & pe_o_5__2_;
  assign N4975 = N4974 & pe_o_5__0_;
  assign N8344 = N4975 & N4978;
  assign N4976 = ~pe_o_5__5_;
  assign N4977 = ~pe_o_5__4_;
  assign N4978 = ~pe_o_5__1_;
  assign N4979 = pe_o_5__6_ & N4984;
  assign N4980 = N4979 & N4985;
  assign N4981 = N4980 & pe_o_5__3_;
  assign N4982 = N4981 & pe_o_5__2_;
  assign N4983 = N4982 & N4986;
  assign N8346 = N4983 & pe_o_5__1_;
  assign N4984 = ~pe_o_5__5_;
  assign N4985 = ~pe_o_5__4_;
  assign N4986 = ~pe_o_5__0_;
  assign N4987 = pe_o_5__6_ & N4992;
  assign N4988 = N4987 & N4993;
  assign N4989 = N4988 & pe_o_5__3_;
  assign N4990 = N4989 & pe_o_5__2_;
  assign N4991 = N4990 & pe_o_5__0_;
  assign N8348 = N4991 & pe_o_5__1_;
  assign N4992 = ~pe_o_5__5_;
  assign N4993 = ~pe_o_5__4_;
  assign N4994 = pe_o_5__6_ & N4999;
  assign N4995 = N4994 & pe_o_5__4_;
  assign N4996 = N4995 & N5000;
  assign N4997 = N4996 & N5001;
  assign N4998 = N4997 & N5002;
  assign N8350 = N4998 & N5003;
  assign N4999 = ~pe_o_5__5_;
  assign N5000 = ~pe_o_5__3_;
  assign N5001 = ~pe_o_5__2_;
  assign N5002 = ~pe_o_5__0_;
  assign N5003 = ~pe_o_5__1_;
  assign N5004 = pe_o_5__6_ & N5009;
  assign N5005 = N5004 & pe_o_5__4_;
  assign N5006 = N5005 & N5010;
  assign N5007 = N5006 & N5011;
  assign N5008 = N5007 & pe_o_5__0_;
  assign N8352 = N5008 & N5012;
  assign N5009 = ~pe_o_5__5_;
  assign N5010 = ~pe_o_5__3_;
  assign N5011 = ~pe_o_5__2_;
  assign N5012 = ~pe_o_5__1_;
  assign N5013 = pe_o_5__6_ & N5018;
  assign N5014 = N5013 & pe_o_5__4_;
  assign N5015 = N5014 & N5019;
  assign N5016 = N5015 & N5020;
  assign N5017 = N5016 & N5021;
  assign N8354 = N5017 & pe_o_5__1_;
  assign N5018 = ~pe_o_5__5_;
  assign N5019 = ~pe_o_5__3_;
  assign N5020 = ~pe_o_5__2_;
  assign N5021 = ~pe_o_5__0_;
  assign N5022 = pe_o_5__6_ & N5027;
  assign N5023 = N5022 & pe_o_5__4_;
  assign N5024 = N5023 & N5028;
  assign N5025 = N5024 & N5029;
  assign N5026 = N5025 & pe_o_5__0_;
  assign N8356 = N5026 & pe_o_5__1_;
  assign N5027 = ~pe_o_5__5_;
  assign N5028 = ~pe_o_5__3_;
  assign N5029 = ~pe_o_5__2_;
  assign N5030 = pe_o_5__6_ & N5035;
  assign N5031 = N5030 & pe_o_5__4_;
  assign N5032 = N5031 & N5036;
  assign N5033 = N5032 & pe_o_5__2_;
  assign N5034 = N5033 & N5037;
  assign N8358 = N5034 & N5038;
  assign N5035 = ~pe_o_5__5_;
  assign N5036 = ~pe_o_5__3_;
  assign N5037 = ~pe_o_5__0_;
  assign N5038 = ~pe_o_5__1_;
  assign N5039 = pe_o_5__6_ & N5044;
  assign N5040 = N5039 & pe_o_5__4_;
  assign N5041 = N5040 & N5045;
  assign N5042 = N5041 & pe_o_5__2_;
  assign N5043 = N5042 & pe_o_5__0_;
  assign N8360 = N5043 & N5046;
  assign N5044 = ~pe_o_5__5_;
  assign N5045 = ~pe_o_5__3_;
  assign N5046 = ~pe_o_5__1_;
  assign N5047 = pe_o_5__6_ & N5052;
  assign N5048 = N5047 & pe_o_5__4_;
  assign N5049 = N5048 & N5053;
  assign N5050 = N5049 & pe_o_5__2_;
  assign N5051 = N5050 & N5054;
  assign N8362 = N5051 & pe_o_5__1_;
  assign N5052 = ~pe_o_5__5_;
  assign N5053 = ~pe_o_5__3_;
  assign N5054 = ~pe_o_5__0_;
  assign N5055 = pe_o_5__6_ & N5060;
  assign N5056 = N5055 & pe_o_5__4_;
  assign N5057 = N5056 & N5061;
  assign N5058 = N5057 & pe_o_5__2_;
  assign N5059 = N5058 & pe_o_5__0_;
  assign N8364 = N5059 & pe_o_5__1_;
  assign N5060 = ~pe_o_5__5_;
  assign N5061 = ~pe_o_5__3_;
  assign N5062 = pe_o_5__6_ & N5067;
  assign N5063 = N5062 & pe_o_5__4_;
  assign N5064 = N5063 & pe_o_5__3_;
  assign N5065 = N5064 & N5068;
  assign N5066 = N5065 & N5069;
  assign N8366 = N5066 & N5070;
  assign N5067 = ~pe_o_5__5_;
  assign N5068 = ~pe_o_5__2_;
  assign N5069 = ~pe_o_5__0_;
  assign N5070 = ~pe_o_5__1_;
  assign N5071 = pe_o_5__6_ & N5076;
  assign N5072 = N5071 & pe_o_5__4_;
  assign N5073 = N5072 & pe_o_5__3_;
  assign N5074 = N5073 & N5077;
  assign N5075 = N5074 & pe_o_5__0_;
  assign N8368 = N5075 & N5078;
  assign N5076 = ~pe_o_5__5_;
  assign N5077 = ~pe_o_5__2_;
  assign N5078 = ~pe_o_5__1_;
  assign N5079 = pe_o_5__6_ & N5084;
  assign N5080 = N5079 & pe_o_5__4_;
  assign N5081 = N5080 & pe_o_5__3_;
  assign N5082 = N5081 & N5085;
  assign N5083 = N5082 & N5086;
  assign N8370 = N5083 & pe_o_5__1_;
  assign N5084 = ~pe_o_5__5_;
  assign N5085 = ~pe_o_5__2_;
  assign N5086 = ~pe_o_5__0_;
  assign N5087 = pe_o_5__6_ & N5092;
  assign N5088 = N5087 & pe_o_5__4_;
  assign N5089 = N5088 & pe_o_5__3_;
  assign N5090 = N5089 & N5093;
  assign N5091 = N5090 & pe_o_5__0_;
  assign N8372 = N5091 & pe_o_5__1_;
  assign N5092 = ~pe_o_5__5_;
  assign N5093 = ~pe_o_5__2_;
  assign N5094 = pe_o_5__6_ & N5099;
  assign N5095 = N5094 & pe_o_5__4_;
  assign N5096 = N5095 & pe_o_5__3_;
  assign N5097 = N5096 & pe_o_5__2_;
  assign N5098 = N5097 & N5100;
  assign N8374 = N5098 & N5101;
  assign N5099 = ~pe_o_5__5_;
  assign N5100 = ~pe_o_5__0_;
  assign N5101 = ~pe_o_5__1_;
  assign N5102 = pe_o_5__6_ & N5107;
  assign N5103 = N5102 & pe_o_5__4_;
  assign N5104 = N5103 & pe_o_5__3_;
  assign N5105 = N5104 & pe_o_5__2_;
  assign N5106 = N5105 & pe_o_5__0_;
  assign N8376 = N5106 & N5108;
  assign N5107 = ~pe_o_5__5_;
  assign N5108 = ~pe_o_5__1_;
  assign N5109 = pe_o_5__6_ & N5114;
  assign N5110 = N5109 & pe_o_5__4_;
  assign N5111 = N5110 & pe_o_5__3_;
  assign N5112 = N5111 & pe_o_5__2_;
  assign N5113 = N5112 & N5115;
  assign N8378 = N5113 & pe_o_5__1_;
  assign N5114 = ~pe_o_5__5_;
  assign N5115 = ~pe_o_5__0_;
  assign N5116 = pe_o_5__6_ & pe_o_5__4_;
  assign N5117 = N5116 & pe_o_5__3_;
  assign N5118 = N5117 & pe_o_5__2_;
  assign N5119 = N5118 & pe_o_5__0_;
  assign N8380 = N5119 & pe_o_5__1_;
  assign N5120 = pe_o_5__6_ & pe_o_5__5_;
  assign N5121 = N5120 & N5125;
  assign N5122 = N5121 & N5126;
  assign N5123 = N5122 & N5127;
  assign N5124 = N5123 & N5128;
  assign N8382 = N5124 & N5129;
  assign N5125 = ~pe_o_5__4_;
  assign N5126 = ~pe_o_5__3_;
  assign N5127 = ~pe_o_5__2_;
  assign N5128 = ~pe_o_5__0_;
  assign N5129 = ~pe_o_5__1_;
  assign N5130 = pe_o_5__6_ & pe_o_5__5_;
  assign N5131 = N5130 & N5135;
  assign N5132 = N5131 & N5136;
  assign N5133 = N5132 & N5137;
  assign N5134 = N5133 & pe_o_5__0_;
  assign N8384 = N5134 & N5138;
  assign N5135 = ~pe_o_5__4_;
  assign N5136 = ~pe_o_5__3_;
  assign N5137 = ~pe_o_5__2_;
  assign N5138 = ~pe_o_5__1_;
  assign N5139 = pe_o_5__6_ & pe_o_5__5_;
  assign N5140 = N5139 & N5144;
  assign N5141 = N5140 & N5145;
  assign N5142 = N5141 & N5146;
  assign N5143 = N5142 & N5147;
  assign N8386 = N5143 & pe_o_5__1_;
  assign N5144 = ~pe_o_5__4_;
  assign N5145 = ~pe_o_5__3_;
  assign N5146 = ~pe_o_5__2_;
  assign N5147 = ~pe_o_5__0_;
  assign N5148 = pe_o_5__6_ & pe_o_5__5_;
  assign N5149 = N5148 & N5153;
  assign N5150 = N5149 & N5154;
  assign N5151 = N5150 & N5155;
  assign N5152 = N5151 & pe_o_5__0_;
  assign N8388 = N5152 & pe_o_5__1_;
  assign N5153 = ~pe_o_5__4_;
  assign N5154 = ~pe_o_5__3_;
  assign N5155 = ~pe_o_5__2_;
  assign N5156 = pe_o_5__6_ & pe_o_5__5_;
  assign N5157 = N5156 & N5161;
  assign N5158 = N5157 & N5162;
  assign N5159 = N5158 & pe_o_5__2_;
  assign N5160 = N5159 & N5163;
  assign N8390 = N5160 & N5164;
  assign N5161 = ~pe_o_5__4_;
  assign N5162 = ~pe_o_5__3_;
  assign N5163 = ~pe_o_5__0_;
  assign N5164 = ~pe_o_5__1_;
  assign N5165 = pe_o_5__6_ & pe_o_5__5_;
  assign N5166 = N5165 & N5170;
  assign N5167 = N5166 & N5171;
  assign N5168 = N5167 & pe_o_5__2_;
  assign N5169 = N5168 & pe_o_5__0_;
  assign N8392 = N5169 & N5172;
  assign N5170 = ~pe_o_5__4_;
  assign N5171 = ~pe_o_5__3_;
  assign N5172 = ~pe_o_5__1_;
  assign N5173 = pe_o_5__6_ & pe_o_5__5_;
  assign N5174 = N5173 & N5178;
  assign N5175 = N5174 & N5179;
  assign N5176 = N5175 & pe_o_5__2_;
  assign N5177 = N5176 & N5180;
  assign N8394 = N5177 & pe_o_5__1_;
  assign N5178 = ~pe_o_5__4_;
  assign N5179 = ~pe_o_5__3_;
  assign N5180 = ~pe_o_5__0_;
  assign N5181 = pe_o_5__6_ & pe_o_5__5_;
  assign N5182 = N5181 & N5186;
  assign N5183 = N5182 & N5187;
  assign N5184 = N5183 & pe_o_5__2_;
  assign N5185 = N5184 & pe_o_5__0_;
  assign N8396 = N5185 & pe_o_5__1_;
  assign N5186 = ~pe_o_5__4_;
  assign N5187 = ~pe_o_5__3_;
  assign N5188 = pe_o_5__6_ & pe_o_5__5_;
  assign N5189 = N5188 & N5193;
  assign N5190 = N5189 & pe_o_5__3_;
  assign N5191 = N5190 & N5194;
  assign N5192 = N5191 & N5195;
  assign N8398 = N5192 & N5196;
  assign N5193 = ~pe_o_5__4_;
  assign N5194 = ~pe_o_5__2_;
  assign N5195 = ~pe_o_5__0_;
  assign N5196 = ~pe_o_5__1_;
  assign N5197 = pe_o_5__6_ & pe_o_5__5_;
  assign N5198 = N5197 & N5202;
  assign N5199 = N5198 & pe_o_5__3_;
  assign N5200 = N5199 & N5203;
  assign N5201 = N5200 & pe_o_5__0_;
  assign N8400 = N5201 & N5204;
  assign N5202 = ~pe_o_5__4_;
  assign N5203 = ~pe_o_5__2_;
  assign N5204 = ~pe_o_5__1_;
  assign N5205 = pe_o_5__6_ & pe_o_5__5_;
  assign N5206 = N5205 & N5210;
  assign N5207 = N5206 & pe_o_5__3_;
  assign N5208 = N5207 & N5211;
  assign N5209 = N5208 & N5212;
  assign N8402 = N5209 & pe_o_5__1_;
  assign N5210 = ~pe_o_5__4_;
  assign N5211 = ~pe_o_5__2_;
  assign N5212 = ~pe_o_5__0_;
  assign N5213 = pe_o_5__6_ & pe_o_5__5_;
  assign N5214 = N5213 & N5218;
  assign N5215 = N5214 & pe_o_5__3_;
  assign N5216 = N5215 & N5219;
  assign N5217 = N5216 & pe_o_5__0_;
  assign N8404 = N5217 & pe_o_5__1_;
  assign N5218 = ~pe_o_5__4_;
  assign N5219 = ~pe_o_5__2_;
  assign N5220 = pe_o_5__6_ & pe_o_5__5_;
  assign N5221 = N5220 & N5225;
  assign N5222 = N5221 & pe_o_5__3_;
  assign N5223 = N5222 & pe_o_5__2_;
  assign N5224 = N5223 & N5226;
  assign N8406 = N5224 & N5227;
  assign N5225 = ~pe_o_5__4_;
  assign N5226 = ~pe_o_5__0_;
  assign N5227 = ~pe_o_5__1_;
  assign N5228 = pe_o_5__6_ & pe_o_5__5_;
  assign N5229 = N5228 & N5233;
  assign N5230 = N5229 & pe_o_5__3_;
  assign N5231 = N5230 & pe_o_5__2_;
  assign N5232 = N5231 & pe_o_5__0_;
  assign N8408 = N5232 & N5234;
  assign N5233 = ~pe_o_5__4_;
  assign N5234 = ~pe_o_5__1_;
  assign N5235 = pe_o_5__6_ & pe_o_5__5_;
  assign N5236 = N5235 & N5240;
  assign N5237 = N5236 & pe_o_5__3_;
  assign N5238 = N5237 & pe_o_5__2_;
  assign N5239 = N5238 & N5241;
  assign N8410 = N5239 & pe_o_5__1_;
  assign N5240 = ~pe_o_5__4_;
  assign N5241 = ~pe_o_5__0_;
  assign N5242 = pe_o_5__6_ & pe_o_5__5_;
  assign N5243 = N5242 & pe_o_5__3_;
  assign N5244 = N5243 & pe_o_5__2_;
  assign N5245 = N5244 & pe_o_5__0_;
  assign N8412 = N5245 & pe_o_5__1_;
  assign N5246 = pe_o_5__6_ & pe_o_5__5_;
  assign N5247 = N5246 & pe_o_5__4_;
  assign N5248 = N5247 & N5251;
  assign N5249 = N5248 & N5252;
  assign N5250 = N5249 & N5253;
  assign N8414 = N5250 & N5254;
  assign N5251 = ~pe_o_5__3_;
  assign N5252 = ~pe_o_5__2_;
  assign N5253 = ~pe_o_5__0_;
  assign N5254 = ~pe_o_5__1_;
  assign N5255 = pe_o_5__6_ & pe_o_5__5_;
  assign N5256 = N5255 & pe_o_5__4_;
  assign N5257 = N5256 & N5260;
  assign N5258 = N5257 & N5261;
  assign N5259 = N5258 & pe_o_5__0_;
  assign N8416 = N5259 & N5262;
  assign N5260 = ~pe_o_5__3_;
  assign N5261 = ~pe_o_5__2_;
  assign N5262 = ~pe_o_5__1_;
  assign N5263 = pe_o_5__6_ & pe_o_5__5_;
  assign N5264 = N5263 & pe_o_5__4_;
  assign N5265 = N5264 & N5268;
  assign N5266 = N5265 & N5269;
  assign N5267 = N5266 & N5270;
  assign N8418 = N5267 & pe_o_5__1_;
  assign N5268 = ~pe_o_5__3_;
  assign N5269 = ~pe_o_5__2_;
  assign N5270 = ~pe_o_5__0_;
  assign N5271 = pe_o_5__6_ & pe_o_5__5_;
  assign N5272 = N5271 & pe_o_5__4_;
  assign N5273 = N5272 & N5276;
  assign N5274 = N5273 & N5277;
  assign N5275 = N5274 & pe_o_5__0_;
  assign N8420 = N5275 & pe_o_5__1_;
  assign N5276 = ~pe_o_5__3_;
  assign N5277 = ~pe_o_5__2_;
  assign N5278 = pe_o_5__6_ & pe_o_5__5_;
  assign N5279 = N5278 & pe_o_5__4_;
  assign N5280 = N5279 & N5283;
  assign N5281 = N5280 & pe_o_5__2_;
  assign N5282 = N5281 & N5284;
  assign N8422 = N5282 & N5285;
  assign N5283 = ~pe_o_5__3_;
  assign N5284 = ~pe_o_5__0_;
  assign N5285 = ~pe_o_5__1_;
  assign N5286 = pe_o_5__6_ & pe_o_5__5_;
  assign N5287 = N5286 & pe_o_5__4_;
  assign N5288 = N5287 & N5291;
  assign N5289 = N5288 & pe_o_5__2_;
  assign N5290 = N5289 & pe_o_5__0_;
  assign N8424 = N5290 & N5292;
  assign N5291 = ~pe_o_5__3_;
  assign N5292 = ~pe_o_5__1_;
  assign N5293 = pe_o_5__6_ & pe_o_5__5_;
  assign N5294 = N5293 & pe_o_5__4_;
  assign N5295 = N5294 & N5298;
  assign N5296 = N5295 & pe_o_5__2_;
  assign N5297 = N5296 & N5299;
  assign N8426 = N5297 & pe_o_5__1_;
  assign N5298 = ~pe_o_5__3_;
  assign N5299 = ~pe_o_5__0_;
  assign N5300 = pe_o_5__6_ & pe_o_5__5_;
  assign N5301 = N5300 & pe_o_5__4_;
  assign N5302 = N5301 & pe_o_5__2_;
  assign N5303 = N5302 & pe_o_5__0_;
  assign N8428 = N5303 & pe_o_5__1_;
  assign N5304 = pe_o_5__6_ & pe_o_5__5_;
  assign N5305 = N5304 & pe_o_5__4_;
  assign N5306 = N5305 & pe_o_5__3_;
  assign N5307 = N5306 & N5309;
  assign N5308 = N5307 & N5310;
  assign N8430 = N5308 & N5311;
  assign N5309 = ~pe_o_5__2_;
  assign N5310 = ~pe_o_5__0_;
  assign N5311 = ~pe_o_5__1_;
  assign N5312 = pe_o_5__6_ & pe_o_5__5_;
  assign N5313 = N5312 & pe_o_5__4_;
  assign N5314 = N5313 & pe_o_5__3_;
  assign N5315 = N5314 & N5317;
  assign N5316 = N5315 & pe_o_5__0_;
  assign N8432 = N5316 & N5318;
  assign N5317 = ~pe_o_5__2_;
  assign N5318 = ~pe_o_5__1_;
  assign N5319 = pe_o_5__6_ & pe_o_5__5_;
  assign N5320 = N5319 & pe_o_5__4_;
  assign N5321 = N5320 & pe_o_5__3_;
  assign N5322 = N5321 & N5324;
  assign N5323 = N5322 & N5325;
  assign N8434 = N5323 & pe_o_5__1_;
  assign N5324 = ~pe_o_5__2_;
  assign N5325 = ~pe_o_5__0_;
  assign N5326 = pe_o_5__6_ & pe_o_5__5_;
  assign N5327 = N5326 & pe_o_5__4_;
  assign N5328 = N5327 & pe_o_5__3_;
  assign N5329 = N5328 & pe_o_5__0_;
  assign N8436 = N5329 & pe_o_5__1_;
  assign N5330 = pe_o_5__6_ & pe_o_5__5_;
  assign N5331 = N5330 & pe_o_5__4_;
  assign N5332 = N5331 & pe_o_5__3_;
  assign N5333 = N5332 & pe_o_5__2_;
  assign N5334 = N5333 & N5335;
  assign N8438 = N5334 & N5336;
  assign N5335 = ~pe_o_5__0_;
  assign N5336 = ~pe_o_5__1_;
  assign N5337 = pe_o_5__6_ & pe_o_5__5_;
  assign N5338 = N5337 & pe_o_5__4_;
  assign N5339 = N5338 & pe_o_5__3_;
  assign N5340 = N5339 & pe_o_5__2_;
  assign N8440 = N5340 & pe_o_5__0_;
  assign N5341 = pe_o_5__6_ & pe_o_5__5_;
  assign N5342 = N5341 & pe_o_5__4_;
  assign N5343 = N5342 & pe_o_5__3_;
  assign N5344 = N5343 & pe_o_5__2_;
  assign N8442 = N5344 & pe_o_5__1_;
  assign N5345 = N5350 & N5351;
  assign N5346 = N5345 & N5352;
  assign N5347 = N5346 & N5353;
  assign N5348 = N5347 & N5354;
  assign N5349 = N5348 & N5355;
  assign N8571 = N5349 & N5356;
  assign N5350 = ~pe_o_6__6_;
  assign N5351 = ~pe_o_6__5_;
  assign N5352 = ~pe_o_6__4_;
  assign N5353 = ~pe_o_6__3_;
  assign N5354 = ~pe_o_6__2_;
  assign N5355 = ~pe_o_6__0_;
  assign N5356 = ~pe_o_6__1_;
  assign N5357 = pe_o_6__6_ & N5362;
  assign N5358 = N5357 & N5363;
  assign N5359 = N5358 & N5364;
  assign N5360 = N5359 & N5365;
  assign N5361 = N5360 & N5366;
  assign N8572 = N5361 & N5367;
  assign N5362 = ~pe_o_6__5_;
  assign N5363 = ~pe_o_6__4_;
  assign N5364 = ~pe_o_6__3_;
  assign N5365 = ~pe_o_6__2_;
  assign N5366 = ~pe_o_6__0_;
  assign N5367 = ~pe_o_6__1_;
  assign N5368 = N5373 & N5374;
  assign N5369 = N5368 & N5375;
  assign N5370 = N5369 & N5376;
  assign N5371 = N5370 & N5377;
  assign N5372 = N5371 & pe_o_6__0_;
  assign N8573 = N5372 & N5378;
  assign N5373 = ~pe_o_6__6_;
  assign N5374 = ~pe_o_6__5_;
  assign N5375 = ~pe_o_6__4_;
  assign N5376 = ~pe_o_6__3_;
  assign N5377 = ~pe_o_6__2_;
  assign N5378 = ~pe_o_6__1_;
  assign N5379 = N5384 & N5385;
  assign N5380 = N5379 & N5386;
  assign N5381 = N5380 & N5387;
  assign N5382 = N5381 & N5388;
  assign N5383 = N5382 & N5389;
  assign N8575 = N5383 & pe_o_6__1_;
  assign N5384 = ~pe_o_6__6_;
  assign N5385 = ~pe_o_6__5_;
  assign N5386 = ~pe_o_6__4_;
  assign N5387 = ~pe_o_6__3_;
  assign N5388 = ~pe_o_6__2_;
  assign N5389 = ~pe_o_6__0_;
  assign N5390 = N5395 & N5396;
  assign N5391 = N5390 & N5397;
  assign N5392 = N5391 & N5398;
  assign N5393 = N5392 & N5399;
  assign N5394 = N5393 & pe_o_6__0_;
  assign N8577 = N5394 & pe_o_6__1_;
  assign N5395 = ~pe_o_6__6_;
  assign N5396 = ~pe_o_6__5_;
  assign N5397 = ~pe_o_6__4_;
  assign N5398 = ~pe_o_6__3_;
  assign N5399 = ~pe_o_6__2_;
  assign N5400 = N5405 & N5406;
  assign N5401 = N5400 & N5407;
  assign N5402 = N5401 & N5408;
  assign N5403 = N5402 & pe_o_6__2_;
  assign N5404 = N5403 & N5409;
  assign N8579 = N5404 & N5410;
  assign N5405 = ~pe_o_6__6_;
  assign N5406 = ~pe_o_6__5_;
  assign N5407 = ~pe_o_6__4_;
  assign N5408 = ~pe_o_6__3_;
  assign N5409 = ~pe_o_6__0_;
  assign N5410 = ~pe_o_6__1_;
  assign N5411 = N5416 & N5417;
  assign N5412 = N5411 & N5418;
  assign N5413 = N5412 & N5419;
  assign N5414 = N5413 & pe_o_6__2_;
  assign N5415 = N5414 & pe_o_6__0_;
  assign N8581 = N5415 & N5420;
  assign N5416 = ~pe_o_6__6_;
  assign N5417 = ~pe_o_6__5_;
  assign N5418 = ~pe_o_6__4_;
  assign N5419 = ~pe_o_6__3_;
  assign N5420 = ~pe_o_6__1_;
  assign N5421 = N5426 & N5427;
  assign N5422 = N5421 & N5428;
  assign N5423 = N5422 & N5429;
  assign N5424 = N5423 & pe_o_6__2_;
  assign N5425 = N5424 & N5430;
  assign N8583 = N5425 & pe_o_6__1_;
  assign N5426 = ~pe_o_6__6_;
  assign N5427 = ~pe_o_6__5_;
  assign N5428 = ~pe_o_6__4_;
  assign N5429 = ~pe_o_6__3_;
  assign N5430 = ~pe_o_6__0_;
  assign N5431 = N5436 & N5437;
  assign N5432 = N5431 & N5438;
  assign N5433 = N5432 & N5439;
  assign N5434 = N5433 & pe_o_6__2_;
  assign N5435 = N5434 & pe_o_6__0_;
  assign N8585 = N5435 & pe_o_6__1_;
  assign N5436 = ~pe_o_6__6_;
  assign N5437 = ~pe_o_6__5_;
  assign N5438 = ~pe_o_6__4_;
  assign N5439 = ~pe_o_6__3_;
  assign N5440 = N5445 & N5446;
  assign N5441 = N5440 & N5447;
  assign N5442 = N5441 & pe_o_6__3_;
  assign N5443 = N5442 & N5448;
  assign N5444 = N5443 & N5449;
  assign N8587 = N5444 & N5450;
  assign N5445 = ~pe_o_6__6_;
  assign N5446 = ~pe_o_6__5_;
  assign N5447 = ~pe_o_6__4_;
  assign N5448 = ~pe_o_6__2_;
  assign N5449 = ~pe_o_6__0_;
  assign N5450 = ~pe_o_6__1_;
  assign N5451 = N5456 & N5457;
  assign N5452 = N5451 & N5458;
  assign N5453 = N5452 & pe_o_6__3_;
  assign N5454 = N5453 & N5459;
  assign N5455 = N5454 & pe_o_6__0_;
  assign N8589 = N5455 & N5460;
  assign N5456 = ~pe_o_6__6_;
  assign N5457 = ~pe_o_6__5_;
  assign N5458 = ~pe_o_6__4_;
  assign N5459 = ~pe_o_6__2_;
  assign N5460 = ~pe_o_6__1_;
  assign N5461 = N5466 & N5467;
  assign N5462 = N5461 & N5468;
  assign N5463 = N5462 & pe_o_6__3_;
  assign N5464 = N5463 & N5469;
  assign N5465 = N5464 & N5470;
  assign N8591 = N5465 & pe_o_6__1_;
  assign N5466 = ~pe_o_6__6_;
  assign N5467 = ~pe_o_6__5_;
  assign N5468 = ~pe_o_6__4_;
  assign N5469 = ~pe_o_6__2_;
  assign N5470 = ~pe_o_6__0_;
  assign N5471 = N5476 & N5477;
  assign N5472 = N5471 & N5478;
  assign N5473 = N5472 & pe_o_6__3_;
  assign N5474 = N5473 & N5479;
  assign N5475 = N5474 & pe_o_6__0_;
  assign N8593 = N5475 & pe_o_6__1_;
  assign N5476 = ~pe_o_6__6_;
  assign N5477 = ~pe_o_6__5_;
  assign N5478 = ~pe_o_6__4_;
  assign N5479 = ~pe_o_6__2_;
  assign N5480 = N5485 & N5486;
  assign N5481 = N5480 & N5487;
  assign N5482 = N5481 & pe_o_6__3_;
  assign N5483 = N5482 & pe_o_6__2_;
  assign N5484 = N5483 & N5488;
  assign N8595 = N5484 & N5489;
  assign N5485 = ~pe_o_6__6_;
  assign N5486 = ~pe_o_6__5_;
  assign N5487 = ~pe_o_6__4_;
  assign N5488 = ~pe_o_6__0_;
  assign N5489 = ~pe_o_6__1_;
  assign N5490 = N5495 & N5496;
  assign N5491 = N5490 & N5497;
  assign N5492 = N5491 & pe_o_6__3_;
  assign N5493 = N5492 & pe_o_6__2_;
  assign N5494 = N5493 & pe_o_6__0_;
  assign N8597 = N5494 & N5498;
  assign N5495 = ~pe_o_6__6_;
  assign N5496 = ~pe_o_6__5_;
  assign N5497 = ~pe_o_6__4_;
  assign N5498 = ~pe_o_6__1_;
  assign N5499 = N5504 & N5505;
  assign N5500 = N5499 & N5506;
  assign N5501 = N5500 & pe_o_6__3_;
  assign N5502 = N5501 & pe_o_6__2_;
  assign N5503 = N5502 & N5507;
  assign N8599 = N5503 & pe_o_6__1_;
  assign N5504 = ~pe_o_6__6_;
  assign N5505 = ~pe_o_6__5_;
  assign N5506 = ~pe_o_6__4_;
  assign N5507 = ~pe_o_6__0_;
  assign N5508 = N5513 & N5514;
  assign N5509 = N5508 & N5515;
  assign N5510 = N5509 & pe_o_6__3_;
  assign N5511 = N5510 & pe_o_6__2_;
  assign N5512 = N5511 & pe_o_6__0_;
  assign N8601 = N5512 & pe_o_6__1_;
  assign N5513 = ~pe_o_6__6_;
  assign N5514 = ~pe_o_6__5_;
  assign N5515 = ~pe_o_6__4_;
  assign N5516 = N5521 & N5522;
  assign N5517 = N5516 & pe_o_6__4_;
  assign N5518 = N5517 & N5523;
  assign N5519 = N5518 & N5524;
  assign N5520 = N5519 & N5525;
  assign N8603 = N5520 & N5526;
  assign N5521 = ~pe_o_6__6_;
  assign N5522 = ~pe_o_6__5_;
  assign N5523 = ~pe_o_6__3_;
  assign N5524 = ~pe_o_6__2_;
  assign N5525 = ~pe_o_6__0_;
  assign N5526 = ~pe_o_6__1_;
  assign N5527 = N5532 & N5533;
  assign N5528 = N5527 & pe_o_6__4_;
  assign N5529 = N5528 & N5534;
  assign N5530 = N5529 & N5535;
  assign N5531 = N5530 & pe_o_6__0_;
  assign N8605 = N5531 & N5536;
  assign N5532 = ~pe_o_6__6_;
  assign N5533 = ~pe_o_6__5_;
  assign N5534 = ~pe_o_6__3_;
  assign N5535 = ~pe_o_6__2_;
  assign N5536 = ~pe_o_6__1_;
  assign N5537 = N5542 & N5543;
  assign N5538 = N5537 & pe_o_6__4_;
  assign N5539 = N5538 & N5544;
  assign N5540 = N5539 & N5545;
  assign N5541 = N5540 & N5546;
  assign N8607 = N5541 & pe_o_6__1_;
  assign N5542 = ~pe_o_6__6_;
  assign N5543 = ~pe_o_6__5_;
  assign N5544 = ~pe_o_6__3_;
  assign N5545 = ~pe_o_6__2_;
  assign N5546 = ~pe_o_6__0_;
  assign N5547 = N5552 & N5553;
  assign N5548 = N5547 & pe_o_6__4_;
  assign N5549 = N5548 & N5554;
  assign N5550 = N5549 & N5555;
  assign N5551 = N5550 & pe_o_6__0_;
  assign N8609 = N5551 & pe_o_6__1_;
  assign N5552 = ~pe_o_6__6_;
  assign N5553 = ~pe_o_6__5_;
  assign N5554 = ~pe_o_6__3_;
  assign N5555 = ~pe_o_6__2_;
  assign N5556 = N5561 & N5562;
  assign N5557 = N5556 & pe_o_6__4_;
  assign N5558 = N5557 & N5563;
  assign N5559 = N5558 & pe_o_6__2_;
  assign N5560 = N5559 & N5564;
  assign N8611 = N5560 & N5565;
  assign N5561 = ~pe_o_6__6_;
  assign N5562 = ~pe_o_6__5_;
  assign N5563 = ~pe_o_6__3_;
  assign N5564 = ~pe_o_6__0_;
  assign N5565 = ~pe_o_6__1_;
  assign N5566 = N5571 & N5572;
  assign N5567 = N5566 & pe_o_6__4_;
  assign N5568 = N5567 & N5573;
  assign N5569 = N5568 & pe_o_6__2_;
  assign N5570 = N5569 & pe_o_6__0_;
  assign N8613 = N5570 & N5574;
  assign N5571 = ~pe_o_6__6_;
  assign N5572 = ~pe_o_6__5_;
  assign N5573 = ~pe_o_6__3_;
  assign N5574 = ~pe_o_6__1_;
  assign N5575 = N5580 & N5581;
  assign N5576 = N5575 & pe_o_6__4_;
  assign N5577 = N5576 & N5582;
  assign N5578 = N5577 & pe_o_6__2_;
  assign N5579 = N5578 & N5583;
  assign N8615 = N5579 & pe_o_6__1_;
  assign N5580 = ~pe_o_6__6_;
  assign N5581 = ~pe_o_6__5_;
  assign N5582 = ~pe_o_6__3_;
  assign N5583 = ~pe_o_6__0_;
  assign N5584 = N5589 & N5590;
  assign N5585 = N5584 & pe_o_6__4_;
  assign N5586 = N5585 & N5591;
  assign N5587 = N5586 & pe_o_6__2_;
  assign N5588 = N5587 & pe_o_6__0_;
  assign N8617 = N5588 & pe_o_6__1_;
  assign N5589 = ~pe_o_6__6_;
  assign N5590 = ~pe_o_6__5_;
  assign N5591 = ~pe_o_6__3_;
  assign N5592 = N5597 & N5598;
  assign N5593 = N5592 & pe_o_6__4_;
  assign N5594 = N5593 & pe_o_6__3_;
  assign N5595 = N5594 & N5599;
  assign N5596 = N5595 & N5600;
  assign N8619 = N5596 & N5601;
  assign N5597 = ~pe_o_6__6_;
  assign N5598 = ~pe_o_6__5_;
  assign N5599 = ~pe_o_6__2_;
  assign N5600 = ~pe_o_6__0_;
  assign N5601 = ~pe_o_6__1_;
  assign N5602 = N5607 & N5608;
  assign N5603 = N5602 & pe_o_6__4_;
  assign N5604 = N5603 & pe_o_6__3_;
  assign N5605 = N5604 & N5609;
  assign N5606 = N5605 & pe_o_6__0_;
  assign N8621 = N5606 & N5610;
  assign N5607 = ~pe_o_6__6_;
  assign N5608 = ~pe_o_6__5_;
  assign N5609 = ~pe_o_6__2_;
  assign N5610 = ~pe_o_6__1_;
  assign N5611 = N5616 & N5617;
  assign N5612 = N5611 & pe_o_6__4_;
  assign N5613 = N5612 & pe_o_6__3_;
  assign N5614 = N5613 & N5618;
  assign N5615 = N5614 & N5619;
  assign N8623 = N5615 & pe_o_6__1_;
  assign N5616 = ~pe_o_6__6_;
  assign N5617 = ~pe_o_6__5_;
  assign N5618 = ~pe_o_6__2_;
  assign N5619 = ~pe_o_6__0_;
  assign N5620 = N5625 & N5626;
  assign N5621 = N5620 & pe_o_6__4_;
  assign N5622 = N5621 & pe_o_6__3_;
  assign N5623 = N5622 & N5627;
  assign N5624 = N5623 & pe_o_6__0_;
  assign N8625 = N5624 & pe_o_6__1_;
  assign N5625 = ~pe_o_6__6_;
  assign N5626 = ~pe_o_6__5_;
  assign N5627 = ~pe_o_6__2_;
  assign N5628 = N5633 & N5634;
  assign N5629 = N5628 & pe_o_6__4_;
  assign N5630 = N5629 & pe_o_6__3_;
  assign N5631 = N5630 & pe_o_6__2_;
  assign N5632 = N5631 & N5635;
  assign N8627 = N5632 & N5636;
  assign N5633 = ~pe_o_6__6_;
  assign N5634 = ~pe_o_6__5_;
  assign N5635 = ~pe_o_6__0_;
  assign N5636 = ~pe_o_6__1_;
  assign N5637 = N5642 & N5643;
  assign N5638 = N5637 & pe_o_6__4_;
  assign N5639 = N5638 & pe_o_6__3_;
  assign N5640 = N5639 & pe_o_6__2_;
  assign N5641 = N5640 & pe_o_6__0_;
  assign N8629 = N5641 & N5644;
  assign N5642 = ~pe_o_6__6_;
  assign N5643 = ~pe_o_6__5_;
  assign N5644 = ~pe_o_6__1_;
  assign N5645 = N5650 & N5651;
  assign N5646 = N5645 & pe_o_6__4_;
  assign N5647 = N5646 & pe_o_6__3_;
  assign N5648 = N5647 & pe_o_6__2_;
  assign N5649 = N5648 & N5652;
  assign N8631 = N5649 & pe_o_6__1_;
  assign N5650 = ~pe_o_6__6_;
  assign N5651 = ~pe_o_6__5_;
  assign N5652 = ~pe_o_6__0_;
  assign N5653 = N5658 & N5659;
  assign N5654 = N5653 & pe_o_6__4_;
  assign N5655 = N5654 & pe_o_6__3_;
  assign N5656 = N5655 & pe_o_6__2_;
  assign N5657 = N5656 & pe_o_6__0_;
  assign N8633 = N5657 & pe_o_6__1_;
  assign N5658 = ~pe_o_6__6_;
  assign N5659 = ~pe_o_6__5_;
  assign N5660 = N5665 & pe_o_6__5_;
  assign N5661 = N5660 & N5666;
  assign N5662 = N5661 & N5667;
  assign N5663 = N5662 & N5668;
  assign N5664 = N5663 & N5669;
  assign N8635 = N5664 & N5670;
  assign N5665 = ~pe_o_6__6_;
  assign N5666 = ~pe_o_6__4_;
  assign N5667 = ~pe_o_6__3_;
  assign N5668 = ~pe_o_6__2_;
  assign N5669 = ~pe_o_6__0_;
  assign N5670 = ~pe_o_6__1_;
  assign N5671 = N5676 & pe_o_6__5_;
  assign N5672 = N5671 & N5677;
  assign N5673 = N5672 & N5678;
  assign N5674 = N5673 & N5679;
  assign N5675 = N5674 & pe_o_6__0_;
  assign N8637 = N5675 & N5680;
  assign N5676 = ~pe_o_6__6_;
  assign N5677 = ~pe_o_6__4_;
  assign N5678 = ~pe_o_6__3_;
  assign N5679 = ~pe_o_6__2_;
  assign N5680 = ~pe_o_6__1_;
  assign N5681 = N5686 & pe_o_6__5_;
  assign N5682 = N5681 & N5687;
  assign N5683 = N5682 & N5688;
  assign N5684 = N5683 & N5689;
  assign N5685 = N5684 & N5690;
  assign N8639 = N5685 & pe_o_6__1_;
  assign N5686 = ~pe_o_6__6_;
  assign N5687 = ~pe_o_6__4_;
  assign N5688 = ~pe_o_6__3_;
  assign N5689 = ~pe_o_6__2_;
  assign N5690 = ~pe_o_6__0_;
  assign N5691 = N5696 & pe_o_6__5_;
  assign N5692 = N5691 & N5697;
  assign N5693 = N5692 & N5698;
  assign N5694 = N5693 & N5699;
  assign N5695 = N5694 & pe_o_6__0_;
  assign N8641 = N5695 & pe_o_6__1_;
  assign N5696 = ~pe_o_6__6_;
  assign N5697 = ~pe_o_6__4_;
  assign N5698 = ~pe_o_6__3_;
  assign N5699 = ~pe_o_6__2_;
  assign N5700 = N5705 & pe_o_6__5_;
  assign N5701 = N5700 & N5706;
  assign N5702 = N5701 & N5707;
  assign N5703 = N5702 & pe_o_6__2_;
  assign N5704 = N5703 & N5708;
  assign N8643 = N5704 & N5709;
  assign N5705 = ~pe_o_6__6_;
  assign N5706 = ~pe_o_6__4_;
  assign N5707 = ~pe_o_6__3_;
  assign N5708 = ~pe_o_6__0_;
  assign N5709 = ~pe_o_6__1_;
  assign N5710 = N5715 & pe_o_6__5_;
  assign N5711 = N5710 & N5716;
  assign N5712 = N5711 & N5717;
  assign N5713 = N5712 & pe_o_6__2_;
  assign N5714 = N5713 & pe_o_6__0_;
  assign N8645 = N5714 & N5718;
  assign N5715 = ~pe_o_6__6_;
  assign N5716 = ~pe_o_6__4_;
  assign N5717 = ~pe_o_6__3_;
  assign N5718 = ~pe_o_6__1_;
  assign N5719 = N5724 & pe_o_6__5_;
  assign N5720 = N5719 & N5725;
  assign N5721 = N5720 & N5726;
  assign N5722 = N5721 & pe_o_6__2_;
  assign N5723 = N5722 & N5727;
  assign N8647 = N5723 & pe_o_6__1_;
  assign N5724 = ~pe_o_6__6_;
  assign N5725 = ~pe_o_6__4_;
  assign N5726 = ~pe_o_6__3_;
  assign N5727 = ~pe_o_6__0_;
  assign N5728 = N5733 & pe_o_6__5_;
  assign N5729 = N5728 & N5734;
  assign N5730 = N5729 & N5735;
  assign N5731 = N5730 & pe_o_6__2_;
  assign N5732 = N5731 & pe_o_6__0_;
  assign N8649 = N5732 & pe_o_6__1_;
  assign N5733 = ~pe_o_6__6_;
  assign N5734 = ~pe_o_6__4_;
  assign N5735 = ~pe_o_6__3_;
  assign N5736 = N5741 & pe_o_6__5_;
  assign N5737 = N5736 & N5742;
  assign N5738 = N5737 & pe_o_6__3_;
  assign N5739 = N5738 & N5743;
  assign N5740 = N5739 & N5744;
  assign N8651 = N5740 & N5745;
  assign N5741 = ~pe_o_6__6_;
  assign N5742 = ~pe_o_6__4_;
  assign N5743 = ~pe_o_6__2_;
  assign N5744 = ~pe_o_6__0_;
  assign N5745 = ~pe_o_6__1_;
  assign N5746 = N5751 & pe_o_6__5_;
  assign N5747 = N5746 & N5752;
  assign N5748 = N5747 & pe_o_6__3_;
  assign N5749 = N5748 & N5753;
  assign N5750 = N5749 & pe_o_6__0_;
  assign N8653 = N5750 & N5754;
  assign N5751 = ~pe_o_6__6_;
  assign N5752 = ~pe_o_6__4_;
  assign N5753 = ~pe_o_6__2_;
  assign N5754 = ~pe_o_6__1_;
  assign N5755 = N5760 & pe_o_6__5_;
  assign N5756 = N5755 & N5761;
  assign N5757 = N5756 & pe_o_6__3_;
  assign N5758 = N5757 & N5762;
  assign N5759 = N5758 & N5763;
  assign N8655 = N5759 & pe_o_6__1_;
  assign N5760 = ~pe_o_6__6_;
  assign N5761 = ~pe_o_6__4_;
  assign N5762 = ~pe_o_6__2_;
  assign N5763 = ~pe_o_6__0_;
  assign N5764 = N5769 & pe_o_6__5_;
  assign N5765 = N5764 & N5770;
  assign N5766 = N5765 & pe_o_6__3_;
  assign N5767 = N5766 & N5771;
  assign N5768 = N5767 & pe_o_6__0_;
  assign N8657 = N5768 & pe_o_6__1_;
  assign N5769 = ~pe_o_6__6_;
  assign N5770 = ~pe_o_6__4_;
  assign N5771 = ~pe_o_6__2_;
  assign N5772 = N5777 & pe_o_6__5_;
  assign N5773 = N5772 & N5778;
  assign N5774 = N5773 & pe_o_6__3_;
  assign N5775 = N5774 & pe_o_6__2_;
  assign N5776 = N5775 & N5779;
  assign N8659 = N5776 & N5780;
  assign N5777 = ~pe_o_6__6_;
  assign N5778 = ~pe_o_6__4_;
  assign N5779 = ~pe_o_6__0_;
  assign N5780 = ~pe_o_6__1_;
  assign N5781 = N5786 & pe_o_6__5_;
  assign N5782 = N5781 & N5787;
  assign N5783 = N5782 & pe_o_6__3_;
  assign N5784 = N5783 & pe_o_6__2_;
  assign N5785 = N5784 & pe_o_6__0_;
  assign N8661 = N5785 & N5788;
  assign N5786 = ~pe_o_6__6_;
  assign N5787 = ~pe_o_6__4_;
  assign N5788 = ~pe_o_6__1_;
  assign N5789 = N5794 & pe_o_6__5_;
  assign N5790 = N5789 & N5795;
  assign N5791 = N5790 & pe_o_6__3_;
  assign N5792 = N5791 & pe_o_6__2_;
  assign N5793 = N5792 & N5796;
  assign N8663 = N5793 & pe_o_6__1_;
  assign N5794 = ~pe_o_6__6_;
  assign N5795 = ~pe_o_6__4_;
  assign N5796 = ~pe_o_6__0_;
  assign N5797 = N5802 & pe_o_6__5_;
  assign N5798 = N5797 & N5803;
  assign N5799 = N5798 & pe_o_6__3_;
  assign N5800 = N5799 & pe_o_6__2_;
  assign N5801 = N5800 & pe_o_6__0_;
  assign N8665 = N5801 & pe_o_6__1_;
  assign N5802 = ~pe_o_6__6_;
  assign N5803 = ~pe_o_6__4_;
  assign N5804 = N5809 & pe_o_6__5_;
  assign N5805 = N5804 & pe_o_6__4_;
  assign N5806 = N5805 & N5810;
  assign N5807 = N5806 & N5811;
  assign N5808 = N5807 & N5812;
  assign N8667 = N5808 & N5813;
  assign N5809 = ~pe_o_6__6_;
  assign N5810 = ~pe_o_6__3_;
  assign N5811 = ~pe_o_6__2_;
  assign N5812 = ~pe_o_6__0_;
  assign N5813 = ~pe_o_6__1_;
  assign N5814 = N5819 & pe_o_6__5_;
  assign N5815 = N5814 & pe_o_6__4_;
  assign N5816 = N5815 & N5820;
  assign N5817 = N5816 & N5821;
  assign N5818 = N5817 & pe_o_6__0_;
  assign N8669 = N5818 & N5822;
  assign N5819 = ~pe_o_6__6_;
  assign N5820 = ~pe_o_6__3_;
  assign N5821 = ~pe_o_6__2_;
  assign N5822 = ~pe_o_6__1_;
  assign N5823 = N5828 & pe_o_6__5_;
  assign N5824 = N5823 & pe_o_6__4_;
  assign N5825 = N5824 & N5829;
  assign N5826 = N5825 & N5830;
  assign N5827 = N5826 & N5831;
  assign N8671 = N5827 & pe_o_6__1_;
  assign N5828 = ~pe_o_6__6_;
  assign N5829 = ~pe_o_6__3_;
  assign N5830 = ~pe_o_6__2_;
  assign N5831 = ~pe_o_6__0_;
  assign N5832 = N5837 & pe_o_6__5_;
  assign N5833 = N5832 & pe_o_6__4_;
  assign N5834 = N5833 & N5838;
  assign N5835 = N5834 & N5839;
  assign N5836 = N5835 & pe_o_6__0_;
  assign N8673 = N5836 & pe_o_6__1_;
  assign N5837 = ~pe_o_6__6_;
  assign N5838 = ~pe_o_6__3_;
  assign N5839 = ~pe_o_6__2_;
  assign N5840 = N5845 & pe_o_6__5_;
  assign N5841 = N5840 & pe_o_6__4_;
  assign N5842 = N5841 & N5846;
  assign N5843 = N5842 & pe_o_6__2_;
  assign N5844 = N5843 & N5847;
  assign N8675 = N5844 & N5848;
  assign N5845 = ~pe_o_6__6_;
  assign N5846 = ~pe_o_6__3_;
  assign N5847 = ~pe_o_6__0_;
  assign N5848 = ~pe_o_6__1_;
  assign N5849 = N5854 & pe_o_6__5_;
  assign N5850 = N5849 & pe_o_6__4_;
  assign N5851 = N5850 & N5855;
  assign N5852 = N5851 & pe_o_6__2_;
  assign N5853 = N5852 & pe_o_6__0_;
  assign N8677 = N5853 & N5856;
  assign N5854 = ~pe_o_6__6_;
  assign N5855 = ~pe_o_6__3_;
  assign N5856 = ~pe_o_6__1_;
  assign N5857 = N5862 & pe_o_6__5_;
  assign N5858 = N5857 & pe_o_6__4_;
  assign N5859 = N5858 & N5863;
  assign N5860 = N5859 & pe_o_6__2_;
  assign N5861 = N5860 & N5864;
  assign N8679 = N5861 & pe_o_6__1_;
  assign N5862 = ~pe_o_6__6_;
  assign N5863 = ~pe_o_6__3_;
  assign N5864 = ~pe_o_6__0_;
  assign N5865 = N5870 & pe_o_6__5_;
  assign N5866 = N5865 & pe_o_6__4_;
  assign N5867 = N5866 & N5871;
  assign N5868 = N5867 & pe_o_6__2_;
  assign N5869 = N5868 & pe_o_6__0_;
  assign N8681 = N5869 & pe_o_6__1_;
  assign N5870 = ~pe_o_6__6_;
  assign N5871 = ~pe_o_6__3_;
  assign N5872 = N5877 & pe_o_6__5_;
  assign N5873 = N5872 & pe_o_6__4_;
  assign N5874 = N5873 & pe_o_6__3_;
  assign N5875 = N5874 & N5878;
  assign N5876 = N5875 & N5879;
  assign N8683 = N5876 & N5880;
  assign N5877 = ~pe_o_6__6_;
  assign N5878 = ~pe_o_6__2_;
  assign N5879 = ~pe_o_6__0_;
  assign N5880 = ~pe_o_6__1_;
  assign N5881 = N5886 & pe_o_6__5_;
  assign N5882 = N5881 & pe_o_6__4_;
  assign N5883 = N5882 & pe_o_6__3_;
  assign N5884 = N5883 & N5887;
  assign N5885 = N5884 & pe_o_6__0_;
  assign N8685 = N5885 & N5888;
  assign N5886 = ~pe_o_6__6_;
  assign N5887 = ~pe_o_6__2_;
  assign N5888 = ~pe_o_6__1_;
  assign N5889 = N5894 & pe_o_6__5_;
  assign N5890 = N5889 & pe_o_6__4_;
  assign N5891 = N5890 & pe_o_6__3_;
  assign N5892 = N5891 & N5895;
  assign N5893 = N5892 & N5896;
  assign N8687 = N5893 & pe_o_6__1_;
  assign N5894 = ~pe_o_6__6_;
  assign N5895 = ~pe_o_6__2_;
  assign N5896 = ~pe_o_6__0_;
  assign N5897 = N5902 & pe_o_6__5_;
  assign N5898 = N5897 & pe_o_6__4_;
  assign N5899 = N5898 & pe_o_6__3_;
  assign N5900 = N5899 & N5903;
  assign N5901 = N5900 & pe_o_6__0_;
  assign N8689 = N5901 & pe_o_6__1_;
  assign N5902 = ~pe_o_6__6_;
  assign N5903 = ~pe_o_6__2_;
  assign N5904 = N5909 & pe_o_6__5_;
  assign N5905 = N5904 & pe_o_6__4_;
  assign N5906 = N5905 & pe_o_6__3_;
  assign N5907 = N5906 & pe_o_6__2_;
  assign N5908 = N5907 & N5910;
  assign N8691 = N5908 & N5911;
  assign N5909 = ~pe_o_6__6_;
  assign N5910 = ~pe_o_6__0_;
  assign N5911 = ~pe_o_6__1_;
  assign N5912 = N5917 & pe_o_6__5_;
  assign N5913 = N5912 & pe_o_6__4_;
  assign N5914 = N5913 & pe_o_6__3_;
  assign N5915 = N5914 & pe_o_6__2_;
  assign N5916 = N5915 & pe_o_6__0_;
  assign N8693 = N5916 & N5918;
  assign N5917 = ~pe_o_6__6_;
  assign N5918 = ~pe_o_6__1_;
  assign N5919 = N5924 & pe_o_6__5_;
  assign N5920 = N5919 & pe_o_6__4_;
  assign N5921 = N5920 & pe_o_6__3_;
  assign N5922 = N5921 & pe_o_6__2_;
  assign N5923 = N5922 & N5925;
  assign N8695 = N5923 & pe_o_6__1_;
  assign N5924 = ~pe_o_6__6_;
  assign N5925 = ~pe_o_6__0_;
  assign N5926 = pe_o_6__5_ & pe_o_6__4_;
  assign N5927 = N5926 & pe_o_6__3_;
  assign N5928 = N5927 & pe_o_6__2_;
  assign N5929 = N5928 & pe_o_6__0_;
  assign N8697 = N5929 & pe_o_6__1_;
  assign N5930 = pe_o_6__6_ & N5935;
  assign N5931 = N5930 & N5936;
  assign N5932 = N5931 & N5937;
  assign N5933 = N5932 & N5938;
  assign N5934 = N5933 & pe_o_6__0_;
  assign N8574 = N5934 & N5939;
  assign N5935 = ~pe_o_6__5_;
  assign N5936 = ~pe_o_6__4_;
  assign N5937 = ~pe_o_6__3_;
  assign N5938 = ~pe_o_6__2_;
  assign N5939 = ~pe_o_6__1_;
  assign N5940 = pe_o_6__6_ & N5945;
  assign N5941 = N5940 & N5946;
  assign N5942 = N5941 & N5947;
  assign N5943 = N5942 & N5948;
  assign N5944 = N5943 & N5949;
  assign N8576 = N5944 & pe_o_6__1_;
  assign N5945 = ~pe_o_6__5_;
  assign N5946 = ~pe_o_6__4_;
  assign N5947 = ~pe_o_6__3_;
  assign N5948 = ~pe_o_6__2_;
  assign N5949 = ~pe_o_6__0_;
  assign N5950 = pe_o_6__6_ & N5955;
  assign N5951 = N5950 & N5956;
  assign N5952 = N5951 & N5957;
  assign N5953 = N5952 & N5958;
  assign N5954 = N5953 & pe_o_6__0_;
  assign N8578 = N5954 & pe_o_6__1_;
  assign N5955 = ~pe_o_6__5_;
  assign N5956 = ~pe_o_6__4_;
  assign N5957 = ~pe_o_6__3_;
  assign N5958 = ~pe_o_6__2_;
  assign N5959 = pe_o_6__6_ & N5964;
  assign N5960 = N5959 & N5965;
  assign N5961 = N5960 & N5966;
  assign N5962 = N5961 & pe_o_6__2_;
  assign N5963 = N5962 & N5967;
  assign N8580 = N5963 & N5968;
  assign N5964 = ~pe_o_6__5_;
  assign N5965 = ~pe_o_6__4_;
  assign N5966 = ~pe_o_6__3_;
  assign N5967 = ~pe_o_6__0_;
  assign N5968 = ~pe_o_6__1_;
  assign N5969 = pe_o_6__6_ & N5974;
  assign N5970 = N5969 & N5975;
  assign N5971 = N5970 & N5976;
  assign N5972 = N5971 & pe_o_6__2_;
  assign N5973 = N5972 & pe_o_6__0_;
  assign N8582 = N5973 & N5977;
  assign N5974 = ~pe_o_6__5_;
  assign N5975 = ~pe_o_6__4_;
  assign N5976 = ~pe_o_6__3_;
  assign N5977 = ~pe_o_6__1_;
  assign N5978 = pe_o_6__6_ & N5983;
  assign N5979 = N5978 & N5984;
  assign N5980 = N5979 & N5985;
  assign N5981 = N5980 & pe_o_6__2_;
  assign N5982 = N5981 & N5986;
  assign N8584 = N5982 & pe_o_6__1_;
  assign N5983 = ~pe_o_6__5_;
  assign N5984 = ~pe_o_6__4_;
  assign N5985 = ~pe_o_6__3_;
  assign N5986 = ~pe_o_6__0_;
  assign N5987 = pe_o_6__6_ & N5992;
  assign N5988 = N5987 & N5993;
  assign N5989 = N5988 & N5994;
  assign N5990 = N5989 & pe_o_6__2_;
  assign N5991 = N5990 & pe_o_6__0_;
  assign N8586 = N5991 & pe_o_6__1_;
  assign N5992 = ~pe_o_6__5_;
  assign N5993 = ~pe_o_6__4_;
  assign N5994 = ~pe_o_6__3_;
  assign N5995 = pe_o_6__6_ & N6000;
  assign N5996 = N5995 & N6001;
  assign N5997 = N5996 & pe_o_6__3_;
  assign N5998 = N5997 & N6002;
  assign N5999 = N5998 & N6003;
  assign N8588 = N5999 & N6004;
  assign N6000 = ~pe_o_6__5_;
  assign N6001 = ~pe_o_6__4_;
  assign N6002 = ~pe_o_6__2_;
  assign N6003 = ~pe_o_6__0_;
  assign N6004 = ~pe_o_6__1_;
  assign N6005 = pe_o_6__6_ & N6010;
  assign N6006 = N6005 & N6011;
  assign N6007 = N6006 & pe_o_6__3_;
  assign N6008 = N6007 & N6012;
  assign N6009 = N6008 & pe_o_6__0_;
  assign N8590 = N6009 & N6013;
  assign N6010 = ~pe_o_6__5_;
  assign N6011 = ~pe_o_6__4_;
  assign N6012 = ~pe_o_6__2_;
  assign N6013 = ~pe_o_6__1_;
  assign N6014 = pe_o_6__6_ & N6019;
  assign N6015 = N6014 & N6020;
  assign N6016 = N6015 & pe_o_6__3_;
  assign N6017 = N6016 & N6021;
  assign N6018 = N6017 & N6022;
  assign N8592 = N6018 & pe_o_6__1_;
  assign N6019 = ~pe_o_6__5_;
  assign N6020 = ~pe_o_6__4_;
  assign N6021 = ~pe_o_6__2_;
  assign N6022 = ~pe_o_6__0_;
  assign N6023 = pe_o_6__6_ & N6028;
  assign N6024 = N6023 & N6029;
  assign N6025 = N6024 & pe_o_6__3_;
  assign N6026 = N6025 & N6030;
  assign N6027 = N6026 & pe_o_6__0_;
  assign N8594 = N6027 & pe_o_6__1_;
  assign N6028 = ~pe_o_6__5_;
  assign N6029 = ~pe_o_6__4_;
  assign N6030 = ~pe_o_6__2_;
  assign N6031 = pe_o_6__6_ & N6036;
  assign N6032 = N6031 & N6037;
  assign N6033 = N6032 & pe_o_6__3_;
  assign N6034 = N6033 & pe_o_6__2_;
  assign N6035 = N6034 & N6038;
  assign N8596 = N6035 & N6039;
  assign N6036 = ~pe_o_6__5_;
  assign N6037 = ~pe_o_6__4_;
  assign N6038 = ~pe_o_6__0_;
  assign N6039 = ~pe_o_6__1_;
  assign N6040 = pe_o_6__6_ & N6045;
  assign N6041 = N6040 & N6046;
  assign N6042 = N6041 & pe_o_6__3_;
  assign N6043 = N6042 & pe_o_6__2_;
  assign N6044 = N6043 & pe_o_6__0_;
  assign N8598 = N6044 & N6047;
  assign N6045 = ~pe_o_6__5_;
  assign N6046 = ~pe_o_6__4_;
  assign N6047 = ~pe_o_6__1_;
  assign N6048 = pe_o_6__6_ & N6053;
  assign N6049 = N6048 & N6054;
  assign N6050 = N6049 & pe_o_6__3_;
  assign N6051 = N6050 & pe_o_6__2_;
  assign N6052 = N6051 & N6055;
  assign N8600 = N6052 & pe_o_6__1_;
  assign N6053 = ~pe_o_6__5_;
  assign N6054 = ~pe_o_6__4_;
  assign N6055 = ~pe_o_6__0_;
  assign N6056 = pe_o_6__6_ & N6061;
  assign N6057 = N6056 & N6062;
  assign N6058 = N6057 & pe_o_6__3_;
  assign N6059 = N6058 & pe_o_6__2_;
  assign N6060 = N6059 & pe_o_6__0_;
  assign N8602 = N6060 & pe_o_6__1_;
  assign N6061 = ~pe_o_6__5_;
  assign N6062 = ~pe_o_6__4_;
  assign N6063 = pe_o_6__6_ & N6068;
  assign N6064 = N6063 & pe_o_6__4_;
  assign N6065 = N6064 & N6069;
  assign N6066 = N6065 & N6070;
  assign N6067 = N6066 & N6071;
  assign N8604 = N6067 & N6072;
  assign N6068 = ~pe_o_6__5_;
  assign N6069 = ~pe_o_6__3_;
  assign N6070 = ~pe_o_6__2_;
  assign N6071 = ~pe_o_6__0_;
  assign N6072 = ~pe_o_6__1_;
  assign N6073 = pe_o_6__6_ & N6078;
  assign N6074 = N6073 & pe_o_6__4_;
  assign N6075 = N6074 & N6079;
  assign N6076 = N6075 & N6080;
  assign N6077 = N6076 & pe_o_6__0_;
  assign N8606 = N6077 & N6081;
  assign N6078 = ~pe_o_6__5_;
  assign N6079 = ~pe_o_6__3_;
  assign N6080 = ~pe_o_6__2_;
  assign N6081 = ~pe_o_6__1_;
  assign N6082 = pe_o_6__6_ & N6087;
  assign N6083 = N6082 & pe_o_6__4_;
  assign N6084 = N6083 & N6088;
  assign N6085 = N6084 & N6089;
  assign N6086 = N6085 & N6090;
  assign N8608 = N6086 & pe_o_6__1_;
  assign N6087 = ~pe_o_6__5_;
  assign N6088 = ~pe_o_6__3_;
  assign N6089 = ~pe_o_6__2_;
  assign N6090 = ~pe_o_6__0_;
  assign N6091 = pe_o_6__6_ & N6096;
  assign N6092 = N6091 & pe_o_6__4_;
  assign N6093 = N6092 & N6097;
  assign N6094 = N6093 & N6098;
  assign N6095 = N6094 & pe_o_6__0_;
  assign N8610 = N6095 & pe_o_6__1_;
  assign N6096 = ~pe_o_6__5_;
  assign N6097 = ~pe_o_6__3_;
  assign N6098 = ~pe_o_6__2_;
  assign N6099 = pe_o_6__6_ & N6104;
  assign N6100 = N6099 & pe_o_6__4_;
  assign N6101 = N6100 & N6105;
  assign N6102 = N6101 & pe_o_6__2_;
  assign N6103 = N6102 & N6106;
  assign N8612 = N6103 & N6107;
  assign N6104 = ~pe_o_6__5_;
  assign N6105 = ~pe_o_6__3_;
  assign N6106 = ~pe_o_6__0_;
  assign N6107 = ~pe_o_6__1_;
  assign N6108 = pe_o_6__6_ & N6113;
  assign N6109 = N6108 & pe_o_6__4_;
  assign N6110 = N6109 & N6114;
  assign N6111 = N6110 & pe_o_6__2_;
  assign N6112 = N6111 & pe_o_6__0_;
  assign N8614 = N6112 & N6115;
  assign N6113 = ~pe_o_6__5_;
  assign N6114 = ~pe_o_6__3_;
  assign N6115 = ~pe_o_6__1_;
  assign N6116 = pe_o_6__6_ & N6121;
  assign N6117 = N6116 & pe_o_6__4_;
  assign N6118 = N6117 & N6122;
  assign N6119 = N6118 & pe_o_6__2_;
  assign N6120 = N6119 & N6123;
  assign N8616 = N6120 & pe_o_6__1_;
  assign N6121 = ~pe_o_6__5_;
  assign N6122 = ~pe_o_6__3_;
  assign N6123 = ~pe_o_6__0_;
  assign N6124 = pe_o_6__6_ & N6129;
  assign N6125 = N6124 & pe_o_6__4_;
  assign N6126 = N6125 & N6130;
  assign N6127 = N6126 & pe_o_6__2_;
  assign N6128 = N6127 & pe_o_6__0_;
  assign N8618 = N6128 & pe_o_6__1_;
  assign N6129 = ~pe_o_6__5_;
  assign N6130 = ~pe_o_6__3_;
  assign N6131 = pe_o_6__6_ & N6136;
  assign N6132 = N6131 & pe_o_6__4_;
  assign N6133 = N6132 & pe_o_6__3_;
  assign N6134 = N6133 & N6137;
  assign N6135 = N6134 & N6138;
  assign N8620 = N6135 & N6139;
  assign N6136 = ~pe_o_6__5_;
  assign N6137 = ~pe_o_6__2_;
  assign N6138 = ~pe_o_6__0_;
  assign N6139 = ~pe_o_6__1_;
  assign N6140 = pe_o_6__6_ & N6145;
  assign N6141 = N6140 & pe_o_6__4_;
  assign N6142 = N6141 & pe_o_6__3_;
  assign N6143 = N6142 & N6146;
  assign N6144 = N6143 & pe_o_6__0_;
  assign N8622 = N6144 & N6147;
  assign N6145 = ~pe_o_6__5_;
  assign N6146 = ~pe_o_6__2_;
  assign N6147 = ~pe_o_6__1_;
  assign N6148 = pe_o_6__6_ & N6153;
  assign N6149 = N6148 & pe_o_6__4_;
  assign N6150 = N6149 & pe_o_6__3_;
  assign N6151 = N6150 & N6154;
  assign N6152 = N6151 & N6155;
  assign N8624 = N6152 & pe_o_6__1_;
  assign N6153 = ~pe_o_6__5_;
  assign N6154 = ~pe_o_6__2_;
  assign N6155 = ~pe_o_6__0_;
  assign N6156 = pe_o_6__6_ & N6161;
  assign N6157 = N6156 & pe_o_6__4_;
  assign N6158 = N6157 & pe_o_6__3_;
  assign N6159 = N6158 & N6162;
  assign N6160 = N6159 & pe_o_6__0_;
  assign N8626 = N6160 & pe_o_6__1_;
  assign N6161 = ~pe_o_6__5_;
  assign N6162 = ~pe_o_6__2_;
  assign N6163 = pe_o_6__6_ & N6168;
  assign N6164 = N6163 & pe_o_6__4_;
  assign N6165 = N6164 & pe_o_6__3_;
  assign N6166 = N6165 & pe_o_6__2_;
  assign N6167 = N6166 & N6169;
  assign N8628 = N6167 & N6170;
  assign N6168 = ~pe_o_6__5_;
  assign N6169 = ~pe_o_6__0_;
  assign N6170 = ~pe_o_6__1_;
  assign N6171 = pe_o_6__6_ & N6176;
  assign N6172 = N6171 & pe_o_6__4_;
  assign N6173 = N6172 & pe_o_6__3_;
  assign N6174 = N6173 & pe_o_6__2_;
  assign N6175 = N6174 & pe_o_6__0_;
  assign N8630 = N6175 & N6177;
  assign N6176 = ~pe_o_6__5_;
  assign N6177 = ~pe_o_6__1_;
  assign N6178 = pe_o_6__6_ & N6183;
  assign N6179 = N6178 & pe_o_6__4_;
  assign N6180 = N6179 & pe_o_6__3_;
  assign N6181 = N6180 & pe_o_6__2_;
  assign N6182 = N6181 & N6184;
  assign N8632 = N6182 & pe_o_6__1_;
  assign N6183 = ~pe_o_6__5_;
  assign N6184 = ~pe_o_6__0_;
  assign N6185 = pe_o_6__6_ & pe_o_6__4_;
  assign N6186 = N6185 & pe_o_6__3_;
  assign N6187 = N6186 & pe_o_6__2_;
  assign N6188 = N6187 & pe_o_6__0_;
  assign N8634 = N6188 & pe_o_6__1_;
  assign N6189 = pe_o_6__6_ & pe_o_6__5_;
  assign N6190 = N6189 & N6194;
  assign N6191 = N6190 & N6195;
  assign N6192 = N6191 & N6196;
  assign N6193 = N6192 & N6197;
  assign N8636 = N6193 & N6198;
  assign N6194 = ~pe_o_6__4_;
  assign N6195 = ~pe_o_6__3_;
  assign N6196 = ~pe_o_6__2_;
  assign N6197 = ~pe_o_6__0_;
  assign N6198 = ~pe_o_6__1_;
  assign N6199 = pe_o_6__6_ & pe_o_6__5_;
  assign N6200 = N6199 & N6204;
  assign N6201 = N6200 & N6205;
  assign N6202 = N6201 & N6206;
  assign N6203 = N6202 & pe_o_6__0_;
  assign N8638 = N6203 & N6207;
  assign N6204 = ~pe_o_6__4_;
  assign N6205 = ~pe_o_6__3_;
  assign N6206 = ~pe_o_6__2_;
  assign N6207 = ~pe_o_6__1_;
  assign N6208 = pe_o_6__6_ & pe_o_6__5_;
  assign N6209 = N6208 & N6213;
  assign N6210 = N6209 & N6214;
  assign N6211 = N6210 & N6215;
  assign N6212 = N6211 & N6216;
  assign N8640 = N6212 & pe_o_6__1_;
  assign N6213 = ~pe_o_6__4_;
  assign N6214 = ~pe_o_6__3_;
  assign N6215 = ~pe_o_6__2_;
  assign N6216 = ~pe_o_6__0_;
  assign N6217 = pe_o_6__6_ & pe_o_6__5_;
  assign N6218 = N6217 & N6222;
  assign N6219 = N6218 & N6223;
  assign N6220 = N6219 & N6224;
  assign N6221 = N6220 & pe_o_6__0_;
  assign N8642 = N6221 & pe_o_6__1_;
  assign N6222 = ~pe_o_6__4_;
  assign N6223 = ~pe_o_6__3_;
  assign N6224 = ~pe_o_6__2_;
  assign N6225 = pe_o_6__6_ & pe_o_6__5_;
  assign N6226 = N6225 & N6230;
  assign N6227 = N6226 & N6231;
  assign N6228 = N6227 & pe_o_6__2_;
  assign N6229 = N6228 & N6232;
  assign N8644 = N6229 & N6233;
  assign N6230 = ~pe_o_6__4_;
  assign N6231 = ~pe_o_6__3_;
  assign N6232 = ~pe_o_6__0_;
  assign N6233 = ~pe_o_6__1_;
  assign N6234 = pe_o_6__6_ & pe_o_6__5_;
  assign N6235 = N6234 & N6239;
  assign N6236 = N6235 & N6240;
  assign N6237 = N6236 & pe_o_6__2_;
  assign N6238 = N6237 & pe_o_6__0_;
  assign N8646 = N6238 & N6241;
  assign N6239 = ~pe_o_6__4_;
  assign N6240 = ~pe_o_6__3_;
  assign N6241 = ~pe_o_6__1_;
  assign N6242 = pe_o_6__6_ & pe_o_6__5_;
  assign N6243 = N6242 & N6247;
  assign N6244 = N6243 & N6248;
  assign N6245 = N6244 & pe_o_6__2_;
  assign N6246 = N6245 & N6249;
  assign N8648 = N6246 & pe_o_6__1_;
  assign N6247 = ~pe_o_6__4_;
  assign N6248 = ~pe_o_6__3_;
  assign N6249 = ~pe_o_6__0_;
  assign N6250 = pe_o_6__6_ & pe_o_6__5_;
  assign N6251 = N6250 & N6255;
  assign N6252 = N6251 & N6256;
  assign N6253 = N6252 & pe_o_6__2_;
  assign N6254 = N6253 & pe_o_6__0_;
  assign N8650 = N6254 & pe_o_6__1_;
  assign N6255 = ~pe_o_6__4_;
  assign N6256 = ~pe_o_6__3_;
  assign N6257 = pe_o_6__6_ & pe_o_6__5_;
  assign N6258 = N6257 & N6262;
  assign N6259 = N6258 & pe_o_6__3_;
  assign N6260 = N6259 & N6263;
  assign N6261 = N6260 & N6264;
  assign N8652 = N6261 & N6265;
  assign N6262 = ~pe_o_6__4_;
  assign N6263 = ~pe_o_6__2_;
  assign N6264 = ~pe_o_6__0_;
  assign N6265 = ~pe_o_6__1_;
  assign N6266 = pe_o_6__6_ & pe_o_6__5_;
  assign N6267 = N6266 & N6271;
  assign N6268 = N6267 & pe_o_6__3_;
  assign N6269 = N6268 & N6272;
  assign N6270 = N6269 & pe_o_6__0_;
  assign N8654 = N6270 & N6273;
  assign N6271 = ~pe_o_6__4_;
  assign N6272 = ~pe_o_6__2_;
  assign N6273 = ~pe_o_6__1_;
  assign N6274 = pe_o_6__6_ & pe_o_6__5_;
  assign N6275 = N6274 & N6279;
  assign N6276 = N6275 & pe_o_6__3_;
  assign N6277 = N6276 & N6280;
  assign N6278 = N6277 & N6281;
  assign N8656 = N6278 & pe_o_6__1_;
  assign N6279 = ~pe_o_6__4_;
  assign N6280 = ~pe_o_6__2_;
  assign N6281 = ~pe_o_6__0_;
  assign N6282 = pe_o_6__6_ & pe_o_6__5_;
  assign N6283 = N6282 & N6287;
  assign N6284 = N6283 & pe_o_6__3_;
  assign N6285 = N6284 & N6288;
  assign N6286 = N6285 & pe_o_6__0_;
  assign N8658 = N6286 & pe_o_6__1_;
  assign N6287 = ~pe_o_6__4_;
  assign N6288 = ~pe_o_6__2_;
  assign N6289 = pe_o_6__6_ & pe_o_6__5_;
  assign N6290 = N6289 & N6294;
  assign N6291 = N6290 & pe_o_6__3_;
  assign N6292 = N6291 & pe_o_6__2_;
  assign N6293 = N6292 & N6295;
  assign N8660 = N6293 & N6296;
  assign N6294 = ~pe_o_6__4_;
  assign N6295 = ~pe_o_6__0_;
  assign N6296 = ~pe_o_6__1_;
  assign N6297 = pe_o_6__6_ & pe_o_6__5_;
  assign N6298 = N6297 & N6302;
  assign N6299 = N6298 & pe_o_6__3_;
  assign N6300 = N6299 & pe_o_6__2_;
  assign N6301 = N6300 & pe_o_6__0_;
  assign N8662 = N6301 & N6303;
  assign N6302 = ~pe_o_6__4_;
  assign N6303 = ~pe_o_6__1_;
  assign N6304 = pe_o_6__6_ & pe_o_6__5_;
  assign N6305 = N6304 & N6309;
  assign N6306 = N6305 & pe_o_6__3_;
  assign N6307 = N6306 & pe_o_6__2_;
  assign N6308 = N6307 & N6310;
  assign N8664 = N6308 & pe_o_6__1_;
  assign N6309 = ~pe_o_6__4_;
  assign N6310 = ~pe_o_6__0_;
  assign N6311 = pe_o_6__6_ & pe_o_6__5_;
  assign N6312 = N6311 & pe_o_6__3_;
  assign N6313 = N6312 & pe_o_6__2_;
  assign N6314 = N6313 & pe_o_6__0_;
  assign N8666 = N6314 & pe_o_6__1_;
  assign N6315 = pe_o_6__6_ & pe_o_6__5_;
  assign N6316 = N6315 & pe_o_6__4_;
  assign N6317 = N6316 & N6320;
  assign N6318 = N6317 & N6321;
  assign N6319 = N6318 & N6322;
  assign N8668 = N6319 & N6323;
  assign N6320 = ~pe_o_6__3_;
  assign N6321 = ~pe_o_6__2_;
  assign N6322 = ~pe_o_6__0_;
  assign N6323 = ~pe_o_6__1_;
  assign N6324 = pe_o_6__6_ & pe_o_6__5_;
  assign N6325 = N6324 & pe_o_6__4_;
  assign N6326 = N6325 & N6329;
  assign N6327 = N6326 & N6330;
  assign N6328 = N6327 & pe_o_6__0_;
  assign N8670 = N6328 & N6331;
  assign N6329 = ~pe_o_6__3_;
  assign N6330 = ~pe_o_6__2_;
  assign N6331 = ~pe_o_6__1_;
  assign N6332 = pe_o_6__6_ & pe_o_6__5_;
  assign N6333 = N6332 & pe_o_6__4_;
  assign N6334 = N6333 & N6337;
  assign N6335 = N6334 & N6338;
  assign N6336 = N6335 & N6339;
  assign N8672 = N6336 & pe_o_6__1_;
  assign N6337 = ~pe_o_6__3_;
  assign N6338 = ~pe_o_6__2_;
  assign N6339 = ~pe_o_6__0_;
  assign N6340 = pe_o_6__6_ & pe_o_6__5_;
  assign N6341 = N6340 & pe_o_6__4_;
  assign N6342 = N6341 & N6345;
  assign N6343 = N6342 & N6346;
  assign N6344 = N6343 & pe_o_6__0_;
  assign N8674 = N6344 & pe_o_6__1_;
  assign N6345 = ~pe_o_6__3_;
  assign N6346 = ~pe_o_6__2_;
  assign N6347 = pe_o_6__6_ & pe_o_6__5_;
  assign N6348 = N6347 & pe_o_6__4_;
  assign N6349 = N6348 & N6352;
  assign N6350 = N6349 & pe_o_6__2_;
  assign N6351 = N6350 & N6353;
  assign N8676 = N6351 & N6354;
  assign N6352 = ~pe_o_6__3_;
  assign N6353 = ~pe_o_6__0_;
  assign N6354 = ~pe_o_6__1_;
  assign N6355 = pe_o_6__6_ & pe_o_6__5_;
  assign N6356 = N6355 & pe_o_6__4_;
  assign N6357 = N6356 & N6360;
  assign N6358 = N6357 & pe_o_6__2_;
  assign N6359 = N6358 & pe_o_6__0_;
  assign N8678 = N6359 & N6361;
  assign N6360 = ~pe_o_6__3_;
  assign N6361 = ~pe_o_6__1_;
  assign N6362 = pe_o_6__6_ & pe_o_6__5_;
  assign N6363 = N6362 & pe_o_6__4_;
  assign N6364 = N6363 & N6367;
  assign N6365 = N6364 & pe_o_6__2_;
  assign N6366 = N6365 & N6368;
  assign N8680 = N6366 & pe_o_6__1_;
  assign N6367 = ~pe_o_6__3_;
  assign N6368 = ~pe_o_6__0_;
  assign N6369 = pe_o_6__6_ & pe_o_6__5_;
  assign N6370 = N6369 & pe_o_6__4_;
  assign N6371 = N6370 & pe_o_6__2_;
  assign N6372 = N6371 & pe_o_6__0_;
  assign N8682 = N6372 & pe_o_6__1_;
  assign N6373 = pe_o_6__6_ & pe_o_6__5_;
  assign N6374 = N6373 & pe_o_6__4_;
  assign N6375 = N6374 & pe_o_6__3_;
  assign N6376 = N6375 & N6378;
  assign N6377 = N6376 & N6379;
  assign N8684 = N6377 & N6380;
  assign N6378 = ~pe_o_6__2_;
  assign N6379 = ~pe_o_6__0_;
  assign N6380 = ~pe_o_6__1_;
  assign N6381 = pe_o_6__6_ & pe_o_6__5_;
  assign N6382 = N6381 & pe_o_6__4_;
  assign N6383 = N6382 & pe_o_6__3_;
  assign N6384 = N6383 & N6386;
  assign N6385 = N6384 & pe_o_6__0_;
  assign N8686 = N6385 & N6387;
  assign N6386 = ~pe_o_6__2_;
  assign N6387 = ~pe_o_6__1_;
  assign N6388 = pe_o_6__6_ & pe_o_6__5_;
  assign N6389 = N6388 & pe_o_6__4_;
  assign N6390 = N6389 & pe_o_6__3_;
  assign N6391 = N6390 & N6393;
  assign N6392 = N6391 & N6394;
  assign N8688 = N6392 & pe_o_6__1_;
  assign N6393 = ~pe_o_6__2_;
  assign N6394 = ~pe_o_6__0_;
  assign N6395 = pe_o_6__6_ & pe_o_6__5_;
  assign N6396 = N6395 & pe_o_6__4_;
  assign N6397 = N6396 & pe_o_6__3_;
  assign N6398 = N6397 & pe_o_6__0_;
  assign N8690 = N6398 & pe_o_6__1_;
  assign N6399 = pe_o_6__6_ & pe_o_6__5_;
  assign N6400 = N6399 & pe_o_6__4_;
  assign N6401 = N6400 & pe_o_6__3_;
  assign N6402 = N6401 & pe_o_6__2_;
  assign N6403 = N6402 & N6404;
  assign N8692 = N6403 & N6405;
  assign N6404 = ~pe_o_6__0_;
  assign N6405 = ~pe_o_6__1_;
  assign N6406 = pe_o_6__6_ & pe_o_6__5_;
  assign N6407 = N6406 & pe_o_6__4_;
  assign N6408 = N6407 & pe_o_6__3_;
  assign N6409 = N6408 & pe_o_6__2_;
  assign N8694 = N6409 & pe_o_6__0_;
  assign N6410 = pe_o_6__6_ & pe_o_6__5_;
  assign N6411 = N6410 & pe_o_6__4_;
  assign N6412 = N6411 & pe_o_6__3_;
  assign N6413 = N6412 & pe_o_6__2_;
  assign N8696 = N6413 & pe_o_6__1_;
  assign way_id_o[5] = (N6414)? lru_i[0] : 
                       (N6415)? lru_i[1] : 
                       (N6416)? lru_i[2] : 
                       (N6417)? lru_i[3] : 
                       (N6418)? lru_i[4] : 
                       (N6419)? lru_i[5] : 
                       (N6420)? lru_i[6] : 
                       (N6421)? lru_i[7] : 
                       (N6422)? lru_i[8] : 
                       (N6423)? lru_i[9] : 
                       (N6424)? lru_i[10] : 
                       (N6425)? lru_i[11] : 
                       (N6426)? lru_i[12] : 
                       (N6427)? lru_i[13] : 
                       (N6428)? lru_i[14] : 
                       (N6429)? lru_i[15] : 
                       (N6430)? lru_i[16] : 
                       (N6431)? lru_i[17] : 
                       (N6432)? lru_i[18] : 
                       (N6433)? lru_i[19] : 
                       (N6434)? lru_i[20] : 
                       (N6435)? lru_i[21] : 
                       (N6436)? lru_i[22] : 
                       (N6437)? lru_i[23] : 
                       (N6438)? lru_i[24] : 
                       (N6439)? lru_i[25] : 
                       (N6440)? lru_i[26] : 
                       (N6441)? lru_i[27] : 
                       (N6442)? lru_i[28] : 
                       (N6443)? lru_i[29] : 
                       (N6444)? lru_i[30] : 
                       (N6445)? lru_i[31] : 
                       (N6446)? lru_i[32] : 
                       (N6447)? lru_i[33] : 
                       (N6448)? lru_i[34] : 
                       (N6449)? lru_i[35] : 
                       (N6450)? lru_i[36] : 
                       (N6451)? lru_i[37] : 
                       (N6452)? lru_i[38] : 
                       (N6453)? lru_i[39] : 
                       (N6454)? lru_i[40] : 
                       (N6455)? lru_i[41] : 
                       (N6456)? lru_i[42] : 
                       (N6457)? lru_i[43] : 
                       (N6458)? lru_i[44] : 
                       (N6459)? lru_i[45] : 
                       (N6460)? lru_i[46] : 
                       (N6461)? lru_i[47] : 
                       (N6462)? lru_i[48] : 
                       (N6463)? lru_i[49] : 
                       (N6464)? lru_i[50] : 
                       (N6465)? lru_i[51] : 
                       (N6466)? lru_i[52] : 
                       (N6467)? lru_i[53] : 
                       (N6468)? lru_i[54] : 
                       (N6469)? lru_i[55] : 
                       (N6470)? lru_i[56] : 
                       (N6471)? lru_i[57] : 
                       (N6472)? lru_i[58] : 
                       (N6473)? lru_i[59] : 
                       (N6474)? lru_i[60] : 
                       (N6475)? lru_i[61] : 
                       (N6476)? lru_i[62] : 
                       (N6477)? lru_i[63] : 
                       (N6478)? lru_i[64] : 
                       (N6479)? lru_i[65] : 
                       (N6480)? lru_i[66] : 
                       (N6481)? lru_i[67] : 
                       (N6482)? lru_i[68] : 
                       (N6483)? lru_i[69] : 
                       (N6484)? lru_i[70] : 
                       (N6485)? lru_i[71] : 
                       (N6486)? lru_i[72] : 
                       (N6487)? lru_i[73] : 
                       (N6488)? lru_i[74] : 
                       (N6489)? lru_i[75] : 
                       (N6490)? lru_i[76] : 
                       (N6491)? lru_i[77] : 
                       (N6492)? lru_i[78] : 
                       (N6493)? lru_i[79] : 
                       (N6494)? lru_i[80] : 
                       (N6495)? lru_i[81] : 
                       (N6496)? lru_i[82] : 
                       (N6497)? lru_i[83] : 
                       (N6498)? lru_i[84] : 
                       (N6499)? lru_i[85] : 
                       (N6500)? lru_i[86] : 
                       (N6501)? lru_i[87] : 
                       (N6502)? lru_i[88] : 
                       (N6503)? lru_i[89] : 
                       (N6504)? lru_i[90] : 
                       (N6505)? lru_i[91] : 
                       (N6506)? lru_i[92] : 
                       (N6507)? lru_i[93] : 
                       (N6508)? lru_i[94] : 
                       (N6509)? lru_i[95] : 
                       (N6510)? lru_i[96] : 
                       (N6511)? lru_i[97] : 
                       (N6512)? lru_i[98] : 
                       (N6513)? lru_i[99] : 
                       (N6514)? lru_i[100] : 
                       (N6515)? lru_i[101] : 
                       (N6516)? lru_i[102] : 
                       (N6517)? lru_i[103] : 
                       (N6518)? lru_i[104] : 
                       (N6519)? lru_i[105] : 
                       (N6520)? lru_i[106] : 
                       (N6521)? lru_i[107] : 
                       (N6522)? lru_i[108] : 
                       (N6523)? lru_i[109] : 
                       (N6524)? lru_i[110] : 
                       (N6525)? lru_i[111] : 
                       (N6526)? lru_i[112] : 
                       (N6527)? lru_i[113] : 
                       (N6528)? lru_i[114] : 
                       (N6529)? lru_i[115] : 
                       (N6530)? lru_i[116] : 
                       (N6531)? lru_i[117] : 
                       (N6532)? lru_i[118] : 
                       (N6533)? lru_i[119] : 
                       (N6534)? lru_i[120] : 
                       (N6535)? lru_i[121] : 
                       (N6536)? lru_i[122] : 
                       (N6537)? lru_i[123] : 
                       (N6538)? lru_i[124] : 
                       (N6539)? lru_i[125] : 
                       (N6540)? lru_i[126] : 1'b0;
  assign N6414 = N7428;
  assign N6415 = N7430;
  assign N6416 = N7432;
  assign N6417 = N7434;
  assign N6418 = N7436;
  assign N6419 = N7438;
  assign N6420 = N7440;
  assign N6421 = N7442;
  assign N6422 = N7444;
  assign N6423 = N7446;
  assign N6424 = N7448;
  assign N6425 = N7450;
  assign N6426 = N7452;
  assign N6427 = N7454;
  assign N6428 = N7456;
  assign N6429 = N7458;
  assign N6430 = N7460;
  assign N6431 = N7462;
  assign N6432 = N7464;
  assign N6433 = N7466;
  assign N6434 = N7468;
  assign N6435 = N7470;
  assign N6436 = N7472;
  assign N6437 = N7474;
  assign N6438 = N7476;
  assign N6439 = N7478;
  assign N6440 = N7480;
  assign N6441 = N7482;
  assign N6442 = N7484;
  assign N6443 = N7486;
  assign N6444 = N7488;
  assign N6445 = N7490;
  assign N6446 = N7492;
  assign N6447 = N7494;
  assign N6448 = N7496;
  assign N6449 = N7498;
  assign N6450 = N7500;
  assign N6451 = N7502;
  assign N6452 = N7504;
  assign N6453 = N7506;
  assign N6454 = N7508;
  assign N6455 = N7510;
  assign N6456 = N7512;
  assign N6457 = N7514;
  assign N6458 = N7516;
  assign N6459 = N7518;
  assign N6460 = N7520;
  assign N6461 = N7522;
  assign N6462 = N7524;
  assign N6463 = N7526;
  assign N6464 = N7528;
  assign N6465 = N7530;
  assign N6466 = N7532;
  assign N6467 = N7534;
  assign N6468 = N7536;
  assign N6469 = N7538;
  assign N6470 = N7540;
  assign N6471 = N7542;
  assign N6472 = N7544;
  assign N6473 = N7546;
  assign N6474 = N7548;
  assign N6475 = N7550;
  assign N6476 = N7552;
  assign N6477 = N7554;
  assign N6478 = N7429;
  assign N6479 = N7431;
  assign N6480 = N7433;
  assign N6481 = N7435;
  assign N6482 = N7437;
  assign N6483 = N7439;
  assign N6484 = N7441;
  assign N6485 = N7443;
  assign N6486 = N7445;
  assign N6487 = N7447;
  assign N6488 = N7449;
  assign N6489 = N7451;
  assign N6490 = N7453;
  assign N6491 = N7455;
  assign N6492 = N7457;
  assign N6493 = N7459;
  assign N6494 = N7461;
  assign N6495 = N7463;
  assign N6496 = N7465;
  assign N6497 = N7467;
  assign N6498 = N7469;
  assign N6499 = N7471;
  assign N6500 = N7473;
  assign N6501 = N7475;
  assign N6502 = N7477;
  assign N6503 = N7479;
  assign N6504 = N7481;
  assign N6505 = N7483;
  assign N6506 = N7485;
  assign N6507 = N7487;
  assign N6508 = N7489;
  assign N6509 = N7491;
  assign N6510 = N7493;
  assign N6511 = N7495;
  assign N6512 = N7497;
  assign N6513 = N7499;
  assign N6514 = N7501;
  assign N6515 = N7503;
  assign N6516 = N7505;
  assign N6517 = N7507;
  assign N6518 = N7509;
  assign N6519 = N7511;
  assign N6520 = N7513;
  assign N6521 = N7515;
  assign N6522 = N7517;
  assign N6523 = N7519;
  assign N6524 = N7521;
  assign N6525 = N7523;
  assign N6526 = N7525;
  assign N6527 = N7527;
  assign N6528 = N7529;
  assign N6529 = N7531;
  assign N6530 = N7533;
  assign N6531 = N7535;
  assign N6532 = N7537;
  assign N6533 = N7539;
  assign N6534 = N7541;
  assign N6535 = N7543;
  assign N6536 = N7545;
  assign N6537 = N7547;
  assign N6538 = N7549;
  assign N6539 = N7551;
  assign N6540 = N7553;
  assign way_id_o[4] = (N6541)? lru_i[0] : 
                       (N6542)? lru_i[1] : 
                       (N6543)? lru_i[2] : 
                       (N6544)? lru_i[3] : 
                       (N6545)? lru_i[4] : 
                       (N6546)? lru_i[5] : 
                       (N6547)? lru_i[6] : 
                       (N6548)? lru_i[7] : 
                       (N6549)? lru_i[8] : 
                       (N6550)? lru_i[9] : 
                       (N6551)? lru_i[10] : 
                       (N6552)? lru_i[11] : 
                       (N6553)? lru_i[12] : 
                       (N6554)? lru_i[13] : 
                       (N6555)? lru_i[14] : 
                       (N6556)? lru_i[15] : 
                       (N6557)? lru_i[16] : 
                       (N6558)? lru_i[17] : 
                       (N6559)? lru_i[18] : 
                       (N6560)? lru_i[19] : 
                       (N6561)? lru_i[20] : 
                       (N6562)? lru_i[21] : 
                       (N6563)? lru_i[22] : 
                       (N6564)? lru_i[23] : 
                       (N6565)? lru_i[24] : 
                       (N6566)? lru_i[25] : 
                       (N6567)? lru_i[26] : 
                       (N6568)? lru_i[27] : 
                       (N6569)? lru_i[28] : 
                       (N6570)? lru_i[29] : 
                       (N6571)? lru_i[30] : 
                       (N6572)? lru_i[31] : 
                       (N6573)? lru_i[32] : 
                       (N6574)? lru_i[33] : 
                       (N6575)? lru_i[34] : 
                       (N6576)? lru_i[35] : 
                       (N6577)? lru_i[36] : 
                       (N6578)? lru_i[37] : 
                       (N6579)? lru_i[38] : 
                       (N6580)? lru_i[39] : 
                       (N6581)? lru_i[40] : 
                       (N6582)? lru_i[41] : 
                       (N6583)? lru_i[42] : 
                       (N6584)? lru_i[43] : 
                       (N6585)? lru_i[44] : 
                       (N6586)? lru_i[45] : 
                       (N6587)? lru_i[46] : 
                       (N6588)? lru_i[47] : 
                       (N6589)? lru_i[48] : 
                       (N6590)? lru_i[49] : 
                       (N6591)? lru_i[50] : 
                       (N6592)? lru_i[51] : 
                       (N6593)? lru_i[52] : 
                       (N6594)? lru_i[53] : 
                       (N6595)? lru_i[54] : 
                       (N6596)? lru_i[55] : 
                       (N6597)? lru_i[56] : 
                       (N6598)? lru_i[57] : 
                       (N6599)? lru_i[58] : 
                       (N6600)? lru_i[59] : 
                       (N6601)? lru_i[60] : 
                       (N6602)? lru_i[61] : 
                       (N6603)? lru_i[62] : 
                       (N6604)? lru_i[63] : 
                       (N6605)? lru_i[64] : 
                       (N6606)? lru_i[65] : 
                       (N6607)? lru_i[66] : 
                       (N6608)? lru_i[67] : 
                       (N6609)? lru_i[68] : 
                       (N6610)? lru_i[69] : 
                       (N6611)? lru_i[70] : 
                       (N6612)? lru_i[71] : 
                       (N6613)? lru_i[72] : 
                       (N6614)? lru_i[73] : 
                       (N6615)? lru_i[74] : 
                       (N6616)? lru_i[75] : 
                       (N6617)? lru_i[76] : 
                       (N6618)? lru_i[77] : 
                       (N6619)? lru_i[78] : 
                       (N6620)? lru_i[79] : 
                       (N6621)? lru_i[80] : 
                       (N6622)? lru_i[81] : 
                       (N6623)? lru_i[82] : 
                       (N6624)? lru_i[83] : 
                       (N6625)? lru_i[84] : 
                       (N6626)? lru_i[85] : 
                       (N6627)? lru_i[86] : 
                       (N6628)? lru_i[87] : 
                       (N6629)? lru_i[88] : 
                       (N6630)? lru_i[89] : 
                       (N6631)? lru_i[90] : 
                       (N6632)? lru_i[91] : 
                       (N6633)? lru_i[92] : 
                       (N6634)? lru_i[93] : 
                       (N6635)? lru_i[94] : 
                       (N6636)? lru_i[95] : 
                       (N6637)? lru_i[96] : 
                       (N6638)? lru_i[97] : 
                       (N6639)? lru_i[98] : 
                       (N6640)? lru_i[99] : 
                       (N6641)? lru_i[100] : 
                       (N6642)? lru_i[101] : 
                       (N6643)? lru_i[102] : 
                       (N6644)? lru_i[103] : 
                       (N6645)? lru_i[104] : 
                       (N6646)? lru_i[105] : 
                       (N6647)? lru_i[106] : 
                       (N6648)? lru_i[107] : 
                       (N6649)? lru_i[108] : 
                       (N6650)? lru_i[109] : 
                       (N6651)? lru_i[110] : 
                       (N6652)? lru_i[111] : 
                       (N6653)? lru_i[112] : 
                       (N6654)? lru_i[113] : 
                       (N6655)? lru_i[114] : 
                       (N6656)? lru_i[115] : 
                       (N6657)? lru_i[116] : 
                       (N6658)? lru_i[117] : 
                       (N6659)? lru_i[118] : 
                       (N6660)? lru_i[119] : 
                       (N6661)? lru_i[120] : 
                       (N6662)? lru_i[121] : 
                       (N6663)? lru_i[122] : 
                       (N6664)? lru_i[123] : 
                       (N6665)? lru_i[124] : 
                       (N6666)? lru_i[125] : 
                       (N6667)? lru_i[126] : 1'b0;
  assign N6541 = N7555;
  assign N6542 = N7557;
  assign N6543 = N7559;
  assign N6544 = N7561;
  assign N6545 = N7563;
  assign N6546 = N7565;
  assign N6547 = N7567;
  assign N6548 = N7569;
  assign N6549 = N7571;
  assign N6550 = N7573;
  assign N6551 = N7575;
  assign N6552 = N7577;
  assign N6553 = N7579;
  assign N6554 = N7581;
  assign N6555 = N7583;
  assign N6556 = N7585;
  assign N6557 = N7587;
  assign N6558 = N7589;
  assign N6559 = N7591;
  assign N6560 = N7593;
  assign N6561 = N7595;
  assign N6562 = N7597;
  assign N6563 = N7599;
  assign N6564 = N7601;
  assign N6565 = N7603;
  assign N6566 = N7605;
  assign N6567 = N7607;
  assign N6568 = N7609;
  assign N6569 = N7611;
  assign N6570 = N7613;
  assign N6571 = N7615;
  assign N6572 = N7617;
  assign N6573 = N7619;
  assign N6574 = N7621;
  assign N6575 = N7623;
  assign N6576 = N7625;
  assign N6577 = N7627;
  assign N6578 = N7629;
  assign N6579 = N7631;
  assign N6580 = N7633;
  assign N6581 = N7635;
  assign N6582 = N7637;
  assign N6583 = N7639;
  assign N6584 = N7641;
  assign N6585 = N7643;
  assign N6586 = N7645;
  assign N6587 = N7647;
  assign N6588 = N7649;
  assign N6589 = N7651;
  assign N6590 = N7653;
  assign N6591 = N7655;
  assign N6592 = N7657;
  assign N6593 = N7659;
  assign N6594 = N7661;
  assign N6595 = N7663;
  assign N6596 = N7665;
  assign N6597 = N7667;
  assign N6598 = N7669;
  assign N6599 = N7671;
  assign N6600 = N7673;
  assign N6601 = N7675;
  assign N6602 = N7677;
  assign N6603 = N7679;
  assign N6604 = N7681;
  assign N6605 = N7556;
  assign N6606 = N7558;
  assign N6607 = N7560;
  assign N6608 = N7562;
  assign N6609 = N7564;
  assign N6610 = N7566;
  assign N6611 = N7568;
  assign N6612 = N7570;
  assign N6613 = N7572;
  assign N6614 = N7574;
  assign N6615 = N7576;
  assign N6616 = N7578;
  assign N6617 = N7580;
  assign N6618 = N7582;
  assign N6619 = N7584;
  assign N6620 = N7586;
  assign N6621 = N7588;
  assign N6622 = N7590;
  assign N6623 = N7592;
  assign N6624 = N7594;
  assign N6625 = N7596;
  assign N6626 = N7598;
  assign N6627 = N7600;
  assign N6628 = N7602;
  assign N6629 = N7604;
  assign N6630 = N7606;
  assign N6631 = N7608;
  assign N6632 = N7610;
  assign N6633 = N7612;
  assign N6634 = N7614;
  assign N6635 = N7616;
  assign N6636 = N7618;
  assign N6637 = N7620;
  assign N6638 = N7622;
  assign N6639 = N7624;
  assign N6640 = N7626;
  assign N6641 = N7628;
  assign N6642 = N7630;
  assign N6643 = N7632;
  assign N6644 = N7634;
  assign N6645 = N7636;
  assign N6646 = N7638;
  assign N6647 = N7640;
  assign N6648 = N7642;
  assign N6649 = N7644;
  assign N6650 = N7646;
  assign N6651 = N7648;
  assign N6652 = N7650;
  assign N6653 = N7652;
  assign N6654 = N7654;
  assign N6655 = N7656;
  assign N6656 = N7658;
  assign N6657 = N7660;
  assign N6658 = N7662;
  assign N6659 = N7664;
  assign N6660 = N7666;
  assign N6661 = N7668;
  assign N6662 = N7670;
  assign N6663 = N7672;
  assign N6664 = N7674;
  assign N6665 = N7676;
  assign N6666 = N7678;
  assign N6667 = N7680;
  assign way_id_o[3] = (N6668)? lru_i[0] : 
                       (N6669)? lru_i[1] : 
                       (N6670)? lru_i[2] : 
                       (N6671)? lru_i[3] : 
                       (N6672)? lru_i[4] : 
                       (N6673)? lru_i[5] : 
                       (N6674)? lru_i[6] : 
                       (N6675)? lru_i[7] : 
                       (N6676)? lru_i[8] : 
                       (N6677)? lru_i[9] : 
                       (N6678)? lru_i[10] : 
                       (N6679)? lru_i[11] : 
                       (N6680)? lru_i[12] : 
                       (N6681)? lru_i[13] : 
                       (N6682)? lru_i[14] : 
                       (N6683)? lru_i[15] : 
                       (N6684)? lru_i[16] : 
                       (N6685)? lru_i[17] : 
                       (N6686)? lru_i[18] : 
                       (N6687)? lru_i[19] : 
                       (N6688)? lru_i[20] : 
                       (N6689)? lru_i[21] : 
                       (N6690)? lru_i[22] : 
                       (N6691)? lru_i[23] : 
                       (N6692)? lru_i[24] : 
                       (N6693)? lru_i[25] : 
                       (N6694)? lru_i[26] : 
                       (N6695)? lru_i[27] : 
                       (N6696)? lru_i[28] : 
                       (N6697)? lru_i[29] : 
                       (N6698)? lru_i[30] : 
                       (N6699)? lru_i[31] : 
                       (N6700)? lru_i[32] : 
                       (N6701)? lru_i[33] : 
                       (N6702)? lru_i[34] : 
                       (N6703)? lru_i[35] : 
                       (N6704)? lru_i[36] : 
                       (N6705)? lru_i[37] : 
                       (N6706)? lru_i[38] : 
                       (N6707)? lru_i[39] : 
                       (N6708)? lru_i[40] : 
                       (N6709)? lru_i[41] : 
                       (N6710)? lru_i[42] : 
                       (N6711)? lru_i[43] : 
                       (N6712)? lru_i[44] : 
                       (N6713)? lru_i[45] : 
                       (N6714)? lru_i[46] : 
                       (N6715)? lru_i[47] : 
                       (N6716)? lru_i[48] : 
                       (N6717)? lru_i[49] : 
                       (N6718)? lru_i[50] : 
                       (N6719)? lru_i[51] : 
                       (N6720)? lru_i[52] : 
                       (N6721)? lru_i[53] : 
                       (N6722)? lru_i[54] : 
                       (N6723)? lru_i[55] : 
                       (N6724)? lru_i[56] : 
                       (N6725)? lru_i[57] : 
                       (N6726)? lru_i[58] : 
                       (N6727)? lru_i[59] : 
                       (N6728)? lru_i[60] : 
                       (N6729)? lru_i[61] : 
                       (N6730)? lru_i[62] : 
                       (N6731)? lru_i[63] : 
                       (N6732)? lru_i[64] : 
                       (N6733)? lru_i[65] : 
                       (N6734)? lru_i[66] : 
                       (N6735)? lru_i[67] : 
                       (N6736)? lru_i[68] : 
                       (N6737)? lru_i[69] : 
                       (N6738)? lru_i[70] : 
                       (N6739)? lru_i[71] : 
                       (N6740)? lru_i[72] : 
                       (N6741)? lru_i[73] : 
                       (N6742)? lru_i[74] : 
                       (N6743)? lru_i[75] : 
                       (N6744)? lru_i[76] : 
                       (N6745)? lru_i[77] : 
                       (N6746)? lru_i[78] : 
                       (N6747)? lru_i[79] : 
                       (N6748)? lru_i[80] : 
                       (N6749)? lru_i[81] : 
                       (N6750)? lru_i[82] : 
                       (N6751)? lru_i[83] : 
                       (N6752)? lru_i[84] : 
                       (N6753)? lru_i[85] : 
                       (N6754)? lru_i[86] : 
                       (N6755)? lru_i[87] : 
                       (N6756)? lru_i[88] : 
                       (N6757)? lru_i[89] : 
                       (N6758)? lru_i[90] : 
                       (N6759)? lru_i[91] : 
                       (N6760)? lru_i[92] : 
                       (N6761)? lru_i[93] : 
                       (N6762)? lru_i[94] : 
                       (N6763)? lru_i[95] : 
                       (N6764)? lru_i[96] : 
                       (N6765)? lru_i[97] : 
                       (N6766)? lru_i[98] : 
                       (N6767)? lru_i[99] : 
                       (N6768)? lru_i[100] : 
                       (N6769)? lru_i[101] : 
                       (N6770)? lru_i[102] : 
                       (N6771)? lru_i[103] : 
                       (N6772)? lru_i[104] : 
                       (N6773)? lru_i[105] : 
                       (N6774)? lru_i[106] : 
                       (N6775)? lru_i[107] : 
                       (N6776)? lru_i[108] : 
                       (N6777)? lru_i[109] : 
                       (N6778)? lru_i[110] : 
                       (N6779)? lru_i[111] : 
                       (N6780)? lru_i[112] : 
                       (N6781)? lru_i[113] : 
                       (N6782)? lru_i[114] : 
                       (N6783)? lru_i[115] : 
                       (N6784)? lru_i[116] : 
                       (N6785)? lru_i[117] : 
                       (N6786)? lru_i[118] : 
                       (N6787)? lru_i[119] : 
                       (N6788)? lru_i[120] : 
                       (N6789)? lru_i[121] : 
                       (N6790)? lru_i[122] : 
                       (N6791)? lru_i[123] : 
                       (N6792)? lru_i[124] : 
                       (N6793)? lru_i[125] : 
                       (N6794)? lru_i[126] : 1'b0;
  assign N6668 = N7809;
  assign N6669 = N7811;
  assign N6670 = N7813;
  assign N6671 = N7815;
  assign N6672 = N7817;
  assign N6673 = N7819;
  assign N6674 = N7821;
  assign N6675 = N7823;
  assign N6676 = N7825;
  assign N6677 = N7827;
  assign N6678 = N7829;
  assign N6679 = N7831;
  assign N6680 = N7833;
  assign N6681 = N7835;
  assign N6682 = N7837;
  assign N6683 = N7839;
  assign N6684 = N7841;
  assign N6685 = N7843;
  assign N6686 = N7845;
  assign N6687 = N7847;
  assign N6688 = N7849;
  assign N6689 = N7851;
  assign N6690 = N7853;
  assign N6691 = N7855;
  assign N6692 = N7857;
  assign N6693 = N7859;
  assign N6694 = N7861;
  assign N6695 = N7863;
  assign N6696 = N7865;
  assign N6697 = N7867;
  assign N6698 = N7869;
  assign N6699 = N7871;
  assign N6700 = N7873;
  assign N6701 = N7875;
  assign N6702 = N7877;
  assign N6703 = N7879;
  assign N6704 = N7881;
  assign N6705 = N7883;
  assign N6706 = N7885;
  assign N6707 = N7887;
  assign N6708 = N7889;
  assign N6709 = N7891;
  assign N6710 = N7893;
  assign N6711 = N7895;
  assign N6712 = N7897;
  assign N6713 = N7899;
  assign N6714 = N7901;
  assign N6715 = N7903;
  assign N6716 = N7905;
  assign N6717 = N7907;
  assign N6718 = N7909;
  assign N6719 = N7911;
  assign N6720 = N7913;
  assign N6721 = N7915;
  assign N6722 = N7917;
  assign N6723 = N7919;
  assign N6724 = N7921;
  assign N6725 = N7923;
  assign N6726 = N7925;
  assign N6727 = N7927;
  assign N6728 = N7929;
  assign N6729 = N7931;
  assign N6730 = N7933;
  assign N6731 = N7935;
  assign N6732 = N7810;
  assign N6733 = N7812;
  assign N6734 = N7814;
  assign N6735 = N7816;
  assign N6736 = N7818;
  assign N6737 = N7820;
  assign N6738 = N7822;
  assign N6739 = N7824;
  assign N6740 = N7826;
  assign N6741 = N7828;
  assign N6742 = N7830;
  assign N6743 = N7832;
  assign N6744 = N7834;
  assign N6745 = N7836;
  assign N6746 = N7838;
  assign N6747 = N7840;
  assign N6748 = N7842;
  assign N6749 = N7844;
  assign N6750 = N7846;
  assign N6751 = N7848;
  assign N6752 = N7850;
  assign N6753 = N7852;
  assign N6754 = N7854;
  assign N6755 = N7856;
  assign N6756 = N7858;
  assign N6757 = N7860;
  assign N6758 = N7862;
  assign N6759 = N7864;
  assign N6760 = N7866;
  assign N6761 = N7868;
  assign N6762 = N7870;
  assign N6763 = N7872;
  assign N6764 = N7874;
  assign N6765 = N7876;
  assign N6766 = N7878;
  assign N6767 = N7880;
  assign N6768 = N7882;
  assign N6769 = N7884;
  assign N6770 = N7886;
  assign N6771 = N7888;
  assign N6772 = N7890;
  assign N6773 = N7892;
  assign N6774 = N7894;
  assign N6775 = N7896;
  assign N6776 = N7898;
  assign N6777 = N7900;
  assign N6778 = N7902;
  assign N6779 = N7904;
  assign N6780 = N7906;
  assign N6781 = N7908;
  assign N6782 = N7910;
  assign N6783 = N7912;
  assign N6784 = N7914;
  assign N6785 = N7916;
  assign N6786 = N7918;
  assign N6787 = N7920;
  assign N6788 = N7922;
  assign N6789 = N7924;
  assign N6790 = N7926;
  assign N6791 = N7928;
  assign N6792 = N7930;
  assign N6793 = N7932;
  assign N6794 = N7934;
  assign way_id_o[2] = (N6795)? lru_i[0] : 
                       (N6796)? lru_i[1] : 
                       (N6797)? lru_i[2] : 
                       (N6798)? lru_i[3] : 
                       (N6799)? lru_i[4] : 
                       (N6800)? lru_i[5] : 
                       (N6801)? lru_i[6] : 
                       (N6802)? lru_i[7] : 
                       (N6803)? lru_i[8] : 
                       (N6804)? lru_i[9] : 
                       (N6805)? lru_i[10] : 
                       (N6806)? lru_i[11] : 
                       (N6807)? lru_i[12] : 
                       (N6808)? lru_i[13] : 
                       (N6809)? lru_i[14] : 
                       (N6810)? lru_i[15] : 
                       (N6811)? lru_i[16] : 
                       (N6812)? lru_i[17] : 
                       (N6813)? lru_i[18] : 
                       (N6814)? lru_i[19] : 
                       (N6815)? lru_i[20] : 
                       (N6816)? lru_i[21] : 
                       (N6817)? lru_i[22] : 
                       (N6818)? lru_i[23] : 
                       (N6819)? lru_i[24] : 
                       (N6820)? lru_i[25] : 
                       (N6821)? lru_i[26] : 
                       (N6822)? lru_i[27] : 
                       (N6823)? lru_i[28] : 
                       (N6824)? lru_i[29] : 
                       (N6825)? lru_i[30] : 
                       (N6826)? lru_i[31] : 
                       (N6827)? lru_i[32] : 
                       (N6828)? lru_i[33] : 
                       (N6829)? lru_i[34] : 
                       (N6830)? lru_i[35] : 
                       (N6831)? lru_i[36] : 
                       (N6832)? lru_i[37] : 
                       (N6833)? lru_i[38] : 
                       (N6834)? lru_i[39] : 
                       (N6835)? lru_i[40] : 
                       (N6836)? lru_i[41] : 
                       (N6837)? lru_i[42] : 
                       (N6838)? lru_i[43] : 
                       (N6839)? lru_i[44] : 
                       (N6840)? lru_i[45] : 
                       (N6841)? lru_i[46] : 
                       (N6842)? lru_i[47] : 
                       (N6843)? lru_i[48] : 
                       (N6844)? lru_i[49] : 
                       (N6845)? lru_i[50] : 
                       (N6846)? lru_i[51] : 
                       (N6847)? lru_i[52] : 
                       (N6848)? lru_i[53] : 
                       (N6849)? lru_i[54] : 
                       (N6850)? lru_i[55] : 
                       (N6851)? lru_i[56] : 
                       (N6852)? lru_i[57] : 
                       (N6853)? lru_i[58] : 
                       (N6854)? lru_i[59] : 
                       (N6855)? lru_i[60] : 
                       (N6856)? lru_i[61] : 
                       (N6857)? lru_i[62] : 
                       (N6858)? lru_i[63] : 
                       (N6859)? lru_i[64] : 
                       (N6860)? lru_i[65] : 
                       (N6861)? lru_i[66] : 
                       (N6862)? lru_i[67] : 
                       (N6863)? lru_i[68] : 
                       (N6864)? lru_i[69] : 
                       (N6865)? lru_i[70] : 
                       (N6866)? lru_i[71] : 
                       (N6867)? lru_i[72] : 
                       (N6868)? lru_i[73] : 
                       (N6869)? lru_i[74] : 
                       (N6870)? lru_i[75] : 
                       (N6871)? lru_i[76] : 
                       (N6872)? lru_i[77] : 
                       (N6873)? lru_i[78] : 
                       (N6874)? lru_i[79] : 
                       (N6875)? lru_i[80] : 
                       (N6876)? lru_i[81] : 
                       (N6877)? lru_i[82] : 
                       (N6878)? lru_i[83] : 
                       (N6879)? lru_i[84] : 
                       (N6880)? lru_i[85] : 
                       (N6881)? lru_i[86] : 
                       (N6882)? lru_i[87] : 
                       (N6883)? lru_i[88] : 
                       (N6884)? lru_i[89] : 
                       (N6885)? lru_i[90] : 
                       (N6886)? lru_i[91] : 
                       (N6887)? lru_i[92] : 
                       (N6888)? lru_i[93] : 
                       (N6889)? lru_i[94] : 
                       (N6890)? lru_i[95] : 
                       (N6891)? lru_i[96] : 
                       (N6892)? lru_i[97] : 
                       (N6893)? lru_i[98] : 
                       (N6894)? lru_i[99] : 
                       (N6895)? lru_i[100] : 
                       (N6896)? lru_i[101] : 
                       (N6897)? lru_i[102] : 
                       (N6898)? lru_i[103] : 
                       (N6899)? lru_i[104] : 
                       (N6900)? lru_i[105] : 
                       (N6901)? lru_i[106] : 
                       (N6902)? lru_i[107] : 
                       (N6903)? lru_i[108] : 
                       (N6904)? lru_i[109] : 
                       (N6905)? lru_i[110] : 
                       (N6906)? lru_i[111] : 
                       (N6907)? lru_i[112] : 
                       (N6908)? lru_i[113] : 
                       (N6909)? lru_i[114] : 
                       (N6910)? lru_i[115] : 
                       (N6911)? lru_i[116] : 
                       (N6912)? lru_i[117] : 
                       (N6913)? lru_i[118] : 
                       (N6914)? lru_i[119] : 
                       (N6915)? lru_i[120] : 
                       (N6916)? lru_i[121] : 
                       (N6917)? lru_i[122] : 
                       (N6918)? lru_i[123] : 
                       (N6919)? lru_i[124] : 
                       (N6920)? lru_i[125] : 
                       (N6921)? lru_i[126] : 1'b0;
  assign N6795 = N8063;
  assign N6796 = N8065;
  assign N6797 = N8067;
  assign N6798 = N8069;
  assign N6799 = N8071;
  assign N6800 = N8073;
  assign N6801 = N8075;
  assign N6802 = N8077;
  assign N6803 = N8079;
  assign N6804 = N8081;
  assign N6805 = N8083;
  assign N6806 = N8085;
  assign N6807 = N8087;
  assign N6808 = N8089;
  assign N6809 = N8091;
  assign N6810 = N8093;
  assign N6811 = N8095;
  assign N6812 = N8097;
  assign N6813 = N8099;
  assign N6814 = N8101;
  assign N6815 = N8103;
  assign N6816 = N8105;
  assign N6817 = N8107;
  assign N6818 = N8109;
  assign N6819 = N8111;
  assign N6820 = N8113;
  assign N6821 = N8115;
  assign N6822 = N8117;
  assign N6823 = N8119;
  assign N6824 = N8121;
  assign N6825 = N8123;
  assign N6826 = N8125;
  assign N6827 = N8127;
  assign N6828 = N8129;
  assign N6829 = N8131;
  assign N6830 = N8133;
  assign N6831 = N8135;
  assign N6832 = N8137;
  assign N6833 = N8139;
  assign N6834 = N8141;
  assign N6835 = N8143;
  assign N6836 = N8145;
  assign N6837 = N8147;
  assign N6838 = N8149;
  assign N6839 = N8151;
  assign N6840 = N8153;
  assign N6841 = N8155;
  assign N6842 = N8157;
  assign N6843 = N8159;
  assign N6844 = N8161;
  assign N6845 = N8163;
  assign N6846 = N8165;
  assign N6847 = N8167;
  assign N6848 = N8169;
  assign N6849 = N8171;
  assign N6850 = N8173;
  assign N6851 = N8175;
  assign N6852 = N8177;
  assign N6853 = N8179;
  assign N6854 = N8181;
  assign N6855 = N8183;
  assign N6856 = N8185;
  assign N6857 = N8187;
  assign N6858 = N8189;
  assign N6859 = N8064;
  assign N6860 = N8066;
  assign N6861 = N8068;
  assign N6862 = N8070;
  assign N6863 = N8072;
  assign N6864 = N8074;
  assign N6865 = N8076;
  assign N6866 = N8078;
  assign N6867 = N8080;
  assign N6868 = N8082;
  assign N6869 = N8084;
  assign N6870 = N8086;
  assign N6871 = N8088;
  assign N6872 = N8090;
  assign N6873 = N8092;
  assign N6874 = N8094;
  assign N6875 = N8096;
  assign N6876 = N8098;
  assign N6877 = N8100;
  assign N6878 = N8102;
  assign N6879 = N8104;
  assign N6880 = N8106;
  assign N6881 = N8108;
  assign N6882 = N8110;
  assign N6883 = N8112;
  assign N6884 = N8114;
  assign N6885 = N8116;
  assign N6886 = N8118;
  assign N6887 = N8120;
  assign N6888 = N8122;
  assign N6889 = N8124;
  assign N6890 = N8126;
  assign N6891 = N8128;
  assign N6892 = N8130;
  assign N6893 = N8132;
  assign N6894 = N8134;
  assign N6895 = N8136;
  assign N6896 = N8138;
  assign N6897 = N8140;
  assign N6898 = N8142;
  assign N6899 = N8144;
  assign N6900 = N8146;
  assign N6901 = N8148;
  assign N6902 = N8150;
  assign N6903 = N8152;
  assign N6904 = N8154;
  assign N6905 = N8156;
  assign N6906 = N8158;
  assign N6907 = N8160;
  assign N6908 = N8162;
  assign N6909 = N8164;
  assign N6910 = N8166;
  assign N6911 = N8168;
  assign N6912 = N8170;
  assign N6913 = N8172;
  assign N6914 = N8174;
  assign N6915 = N8176;
  assign N6916 = N8178;
  assign N6917 = N8180;
  assign N6918 = N8182;
  assign N6919 = N8184;
  assign N6920 = N8186;
  assign N6921 = N8188;
  assign way_id_o[1] = (N6922)? lru_i[0] : 
                       (N6923)? lru_i[1] : 
                       (N6924)? lru_i[2] : 
                       (N6925)? lru_i[3] : 
                       (N6926)? lru_i[4] : 
                       (N6927)? lru_i[5] : 
                       (N6928)? lru_i[6] : 
                       (N6929)? lru_i[7] : 
                       (N6930)? lru_i[8] : 
                       (N6931)? lru_i[9] : 
                       (N6932)? lru_i[10] : 
                       (N6933)? lru_i[11] : 
                       (N6934)? lru_i[12] : 
                       (N6935)? lru_i[13] : 
                       (N6936)? lru_i[14] : 
                       (N6937)? lru_i[15] : 
                       (N6938)? lru_i[16] : 
                       (N6939)? lru_i[17] : 
                       (N6940)? lru_i[18] : 
                       (N6941)? lru_i[19] : 
                       (N6942)? lru_i[20] : 
                       (N6943)? lru_i[21] : 
                       (N6944)? lru_i[22] : 
                       (N6945)? lru_i[23] : 
                       (N6946)? lru_i[24] : 
                       (N6947)? lru_i[25] : 
                       (N6948)? lru_i[26] : 
                       (N6949)? lru_i[27] : 
                       (N6950)? lru_i[28] : 
                       (N6951)? lru_i[29] : 
                       (N6952)? lru_i[30] : 
                       (N6953)? lru_i[31] : 
                       (N6954)? lru_i[32] : 
                       (N6955)? lru_i[33] : 
                       (N6956)? lru_i[34] : 
                       (N6957)? lru_i[35] : 
                       (N6958)? lru_i[36] : 
                       (N6959)? lru_i[37] : 
                       (N6960)? lru_i[38] : 
                       (N6961)? lru_i[39] : 
                       (N6962)? lru_i[40] : 
                       (N6963)? lru_i[41] : 
                       (N6964)? lru_i[42] : 
                       (N6965)? lru_i[43] : 
                       (N6966)? lru_i[44] : 
                       (N6967)? lru_i[45] : 
                       (N6968)? lru_i[46] : 
                       (N6969)? lru_i[47] : 
                       (N6970)? lru_i[48] : 
                       (N6971)? lru_i[49] : 
                       (N6972)? lru_i[50] : 
                       (N6973)? lru_i[51] : 
                       (N6974)? lru_i[52] : 
                       (N6975)? lru_i[53] : 
                       (N6976)? lru_i[54] : 
                       (N6977)? lru_i[55] : 
                       (N6978)? lru_i[56] : 
                       (N6979)? lru_i[57] : 
                       (N6980)? lru_i[58] : 
                       (N6981)? lru_i[59] : 
                       (N6982)? lru_i[60] : 
                       (N6983)? lru_i[61] : 
                       (N6984)? lru_i[62] : 
                       (N6985)? lru_i[63] : 
                       (N6986)? lru_i[64] : 
                       (N6987)? lru_i[65] : 
                       (N6988)? lru_i[66] : 
                       (N6989)? lru_i[67] : 
                       (N6990)? lru_i[68] : 
                       (N6991)? lru_i[69] : 
                       (N6992)? lru_i[70] : 
                       (N6993)? lru_i[71] : 
                       (N6994)? lru_i[72] : 
                       (N6995)? lru_i[73] : 
                       (N6996)? lru_i[74] : 
                       (N6997)? lru_i[75] : 
                       (N6998)? lru_i[76] : 
                       (N6999)? lru_i[77] : 
                       (N7000)? lru_i[78] : 
                       (N7001)? lru_i[79] : 
                       (N7002)? lru_i[80] : 
                       (N7003)? lru_i[81] : 
                       (N7004)? lru_i[82] : 
                       (N7005)? lru_i[83] : 
                       (N7006)? lru_i[84] : 
                       (N7007)? lru_i[85] : 
                       (N7008)? lru_i[86] : 
                       (N7009)? lru_i[87] : 
                       (N7010)? lru_i[88] : 
                       (N7011)? lru_i[89] : 
                       (N7012)? lru_i[90] : 
                       (N7013)? lru_i[91] : 
                       (N7014)? lru_i[92] : 
                       (N7015)? lru_i[93] : 
                       (N7016)? lru_i[94] : 
                       (N7017)? lru_i[95] : 
                       (N7018)? lru_i[96] : 
                       (N7019)? lru_i[97] : 
                       (N7020)? lru_i[98] : 
                       (N7021)? lru_i[99] : 
                       (N7022)? lru_i[100] : 
                       (N7023)? lru_i[101] : 
                       (N7024)? lru_i[102] : 
                       (N7025)? lru_i[103] : 
                       (N7026)? lru_i[104] : 
                       (N7027)? lru_i[105] : 
                       (N7028)? lru_i[106] : 
                       (N7029)? lru_i[107] : 
                       (N7030)? lru_i[108] : 
                       (N7031)? lru_i[109] : 
                       (N7032)? lru_i[110] : 
                       (N7033)? lru_i[111] : 
                       (N7034)? lru_i[112] : 
                       (N7035)? lru_i[113] : 
                       (N7036)? lru_i[114] : 
                       (N7037)? lru_i[115] : 
                       (N7038)? lru_i[116] : 
                       (N7039)? lru_i[117] : 
                       (N7040)? lru_i[118] : 
                       (N7041)? lru_i[119] : 
                       (N7042)? lru_i[120] : 
                       (N7043)? lru_i[121] : 
                       (N7044)? lru_i[122] : 
                       (N7045)? lru_i[123] : 
                       (N7046)? lru_i[124] : 
                       (N7047)? lru_i[125] : 
                       (N7048)? lru_i[126] : 1'b0;
  assign N6922 = N8317;
  assign N6923 = N8319;
  assign N6924 = N8321;
  assign N6925 = N8323;
  assign N6926 = N8325;
  assign N6927 = N8327;
  assign N6928 = N8329;
  assign N6929 = N8331;
  assign N6930 = N8333;
  assign N6931 = N8335;
  assign N6932 = N8337;
  assign N6933 = N8339;
  assign N6934 = N8341;
  assign N6935 = N8343;
  assign N6936 = N8345;
  assign N6937 = N8347;
  assign N6938 = N8349;
  assign N6939 = N8351;
  assign N6940 = N8353;
  assign N6941 = N8355;
  assign N6942 = N8357;
  assign N6943 = N8359;
  assign N6944 = N8361;
  assign N6945 = N8363;
  assign N6946 = N8365;
  assign N6947 = N8367;
  assign N6948 = N8369;
  assign N6949 = N8371;
  assign N6950 = N8373;
  assign N6951 = N8375;
  assign N6952 = N8377;
  assign N6953 = N8379;
  assign N6954 = N8381;
  assign N6955 = N8383;
  assign N6956 = N8385;
  assign N6957 = N8387;
  assign N6958 = N8389;
  assign N6959 = N8391;
  assign N6960 = N8393;
  assign N6961 = N8395;
  assign N6962 = N8397;
  assign N6963 = N8399;
  assign N6964 = N8401;
  assign N6965 = N8403;
  assign N6966 = N8405;
  assign N6967 = N8407;
  assign N6968 = N8409;
  assign N6969 = N8411;
  assign N6970 = N8413;
  assign N6971 = N8415;
  assign N6972 = N8417;
  assign N6973 = N8419;
  assign N6974 = N8421;
  assign N6975 = N8423;
  assign N6976 = N8425;
  assign N6977 = N8427;
  assign N6978 = N8429;
  assign N6979 = N8431;
  assign N6980 = N8433;
  assign N6981 = N8435;
  assign N6982 = N8437;
  assign N6983 = N8439;
  assign N6984 = N8441;
  assign N6985 = N8443;
  assign N6986 = N8318;
  assign N6987 = N8320;
  assign N6988 = N8322;
  assign N6989 = N8324;
  assign N6990 = N8326;
  assign N6991 = N8328;
  assign N6992 = N8330;
  assign N6993 = N8332;
  assign N6994 = N8334;
  assign N6995 = N8336;
  assign N6996 = N8338;
  assign N6997 = N8340;
  assign N6998 = N8342;
  assign N6999 = N8344;
  assign N7000 = N8346;
  assign N7001 = N8348;
  assign N7002 = N8350;
  assign N7003 = N8352;
  assign N7004 = N8354;
  assign N7005 = N8356;
  assign N7006 = N8358;
  assign N7007 = N8360;
  assign N7008 = N8362;
  assign N7009 = N8364;
  assign N7010 = N8366;
  assign N7011 = N8368;
  assign N7012 = N8370;
  assign N7013 = N8372;
  assign N7014 = N8374;
  assign N7015 = N8376;
  assign N7016 = N8378;
  assign N7017 = N8380;
  assign N7018 = N8382;
  assign N7019 = N8384;
  assign N7020 = N8386;
  assign N7021 = N8388;
  assign N7022 = N8390;
  assign N7023 = N8392;
  assign N7024 = N8394;
  assign N7025 = N8396;
  assign N7026 = N8398;
  assign N7027 = N8400;
  assign N7028 = N8402;
  assign N7029 = N8404;
  assign N7030 = N8406;
  assign N7031 = N8408;
  assign N7032 = N8410;
  assign N7033 = N8412;
  assign N7034 = N8414;
  assign N7035 = N8416;
  assign N7036 = N8418;
  assign N7037 = N8420;
  assign N7038 = N8422;
  assign N7039 = N8424;
  assign N7040 = N8426;
  assign N7041 = N8428;
  assign N7042 = N8430;
  assign N7043 = N8432;
  assign N7044 = N8434;
  assign N7045 = N8436;
  assign N7046 = N8438;
  assign N7047 = N8440;
  assign N7048 = N8442;
  assign way_id_o[0] = (N7049)? lru_i[0] : 
                       (N7050)? lru_i[1] : 
                       (N7051)? lru_i[2] : 
                       (N7052)? lru_i[3] : 
                       (N7053)? lru_i[4] : 
                       (N7054)? lru_i[5] : 
                       (N7055)? lru_i[6] : 
                       (N7056)? lru_i[7] : 
                       (N7057)? lru_i[8] : 
                       (N7058)? lru_i[9] : 
                       (N7059)? lru_i[10] : 
                       (N7060)? lru_i[11] : 
                       (N7061)? lru_i[12] : 
                       (N7062)? lru_i[13] : 
                       (N7063)? lru_i[14] : 
                       (N7064)? lru_i[15] : 
                       (N7065)? lru_i[16] : 
                       (N7066)? lru_i[17] : 
                       (N7067)? lru_i[18] : 
                       (N7068)? lru_i[19] : 
                       (N7069)? lru_i[20] : 
                       (N7070)? lru_i[21] : 
                       (N7071)? lru_i[22] : 
                       (N7072)? lru_i[23] : 
                       (N7073)? lru_i[24] : 
                       (N7074)? lru_i[25] : 
                       (N7075)? lru_i[26] : 
                       (N7076)? lru_i[27] : 
                       (N7077)? lru_i[28] : 
                       (N7078)? lru_i[29] : 
                       (N7079)? lru_i[30] : 
                       (N7080)? lru_i[31] : 
                       (N7081)? lru_i[32] : 
                       (N7082)? lru_i[33] : 
                       (N7083)? lru_i[34] : 
                       (N7084)? lru_i[35] : 
                       (N7085)? lru_i[36] : 
                       (N7086)? lru_i[37] : 
                       (N7087)? lru_i[38] : 
                       (N7088)? lru_i[39] : 
                       (N7089)? lru_i[40] : 
                       (N7090)? lru_i[41] : 
                       (N7091)? lru_i[42] : 
                       (N7092)? lru_i[43] : 
                       (N7093)? lru_i[44] : 
                       (N7094)? lru_i[45] : 
                       (N7095)? lru_i[46] : 
                       (N7096)? lru_i[47] : 
                       (N7097)? lru_i[48] : 
                       (N7098)? lru_i[49] : 
                       (N7099)? lru_i[50] : 
                       (N7100)? lru_i[51] : 
                       (N7101)? lru_i[52] : 
                       (N7102)? lru_i[53] : 
                       (N7103)? lru_i[54] : 
                       (N7104)? lru_i[55] : 
                       (N7105)? lru_i[56] : 
                       (N7106)? lru_i[57] : 
                       (N7107)? lru_i[58] : 
                       (N7108)? lru_i[59] : 
                       (N7109)? lru_i[60] : 
                       (N7110)? lru_i[61] : 
                       (N7111)? lru_i[62] : 
                       (N7112)? lru_i[63] : 
                       (N7113)? lru_i[64] : 
                       (N7114)? lru_i[65] : 
                       (N7115)? lru_i[66] : 
                       (N7116)? lru_i[67] : 
                       (N7117)? lru_i[68] : 
                       (N7118)? lru_i[69] : 
                       (N7119)? lru_i[70] : 
                       (N7120)? lru_i[71] : 
                       (N7121)? lru_i[72] : 
                       (N7122)? lru_i[73] : 
                       (N7123)? lru_i[74] : 
                       (N7124)? lru_i[75] : 
                       (N7125)? lru_i[76] : 
                       (N7126)? lru_i[77] : 
                       (N7127)? lru_i[78] : 
                       (N7128)? lru_i[79] : 
                       (N7129)? lru_i[80] : 
                       (N7130)? lru_i[81] : 
                       (N7131)? lru_i[82] : 
                       (N7132)? lru_i[83] : 
                       (N7133)? lru_i[84] : 
                       (N7134)? lru_i[85] : 
                       (N7135)? lru_i[86] : 
                       (N7136)? lru_i[87] : 
                       (N7137)? lru_i[88] : 
                       (N7138)? lru_i[89] : 
                       (N7139)? lru_i[90] : 
                       (N7140)? lru_i[91] : 
                       (N7141)? lru_i[92] : 
                       (N7142)? lru_i[93] : 
                       (N7143)? lru_i[94] : 
                       (N7144)? lru_i[95] : 
                       (N7145)? lru_i[96] : 
                       (N7146)? lru_i[97] : 
                       (N7147)? lru_i[98] : 
                       (N7148)? lru_i[99] : 
                       (N7149)? lru_i[100] : 
                       (N7150)? lru_i[101] : 
                       (N7151)? lru_i[102] : 
                       (N7152)? lru_i[103] : 
                       (N7153)? lru_i[104] : 
                       (N7154)? lru_i[105] : 
                       (N7155)? lru_i[106] : 
                       (N7156)? lru_i[107] : 
                       (N7157)? lru_i[108] : 
                       (N7158)? lru_i[109] : 
                       (N7159)? lru_i[110] : 
                       (N7160)? lru_i[111] : 
                       (N7161)? lru_i[112] : 
                       (N7162)? lru_i[113] : 
                       (N7163)? lru_i[114] : 
                       (N7164)? lru_i[115] : 
                       (N7165)? lru_i[116] : 
                       (N7166)? lru_i[117] : 
                       (N7167)? lru_i[118] : 
                       (N7168)? lru_i[119] : 
                       (N7169)? lru_i[120] : 
                       (N7170)? lru_i[121] : 
                       (N7171)? lru_i[122] : 
                       (N7172)? lru_i[123] : 
                       (N7173)? lru_i[124] : 
                       (N7174)? lru_i[125] : 
                       (N7175)? lru_i[126] : 1'b0;
  assign N7049 = N8571;
  assign N7050 = N8573;
  assign N7051 = N8575;
  assign N7052 = N8577;
  assign N7053 = N8579;
  assign N7054 = N8581;
  assign N7055 = N8583;
  assign N7056 = N8585;
  assign N7057 = N8587;
  assign N7058 = N8589;
  assign N7059 = N8591;
  assign N7060 = N8593;
  assign N7061 = N8595;
  assign N7062 = N8597;
  assign N7063 = N8599;
  assign N7064 = N8601;
  assign N7065 = N8603;
  assign N7066 = N8605;
  assign N7067 = N8607;
  assign N7068 = N8609;
  assign N7069 = N8611;
  assign N7070 = N8613;
  assign N7071 = N8615;
  assign N7072 = N8617;
  assign N7073 = N8619;
  assign N7074 = N8621;
  assign N7075 = N8623;
  assign N7076 = N8625;
  assign N7077 = N8627;
  assign N7078 = N8629;
  assign N7079 = N8631;
  assign N7080 = N8633;
  assign N7081 = N8635;
  assign N7082 = N8637;
  assign N7083 = N8639;
  assign N7084 = N8641;
  assign N7085 = N8643;
  assign N7086 = N8645;
  assign N7087 = N8647;
  assign N7088 = N8649;
  assign N7089 = N8651;
  assign N7090 = N8653;
  assign N7091 = N8655;
  assign N7092 = N8657;
  assign N7093 = N8659;
  assign N7094 = N8661;
  assign N7095 = N8663;
  assign N7096 = N8665;
  assign N7097 = N8667;
  assign N7098 = N8669;
  assign N7099 = N8671;
  assign N7100 = N8673;
  assign N7101 = N8675;
  assign N7102 = N8677;
  assign N7103 = N8679;
  assign N7104 = N8681;
  assign N7105 = N8683;
  assign N7106 = N8685;
  assign N7107 = N8687;
  assign N7108 = N8689;
  assign N7109 = N8691;
  assign N7110 = N8693;
  assign N7111 = N8695;
  assign N7112 = N8697;
  assign N7113 = N8572;
  assign N7114 = N8574;
  assign N7115 = N8576;
  assign N7116 = N8578;
  assign N7117 = N8580;
  assign N7118 = N8582;
  assign N7119 = N8584;
  assign N7120 = N8586;
  assign N7121 = N8588;
  assign N7122 = N8590;
  assign N7123 = N8592;
  assign N7124 = N8594;
  assign N7125 = N8596;
  assign N7126 = N8598;
  assign N7127 = N8600;
  assign N7128 = N8602;
  assign N7129 = N8604;
  assign N7130 = N8606;
  assign N7131 = N8608;
  assign N7132 = N8610;
  assign N7133 = N8612;
  assign N7134 = N8614;
  assign N7135 = N8616;
  assign N7136 = N8618;
  assign N7137 = N8620;
  assign N7138 = N8622;
  assign N7139 = N8624;
  assign N7140 = N8626;
  assign N7141 = N8628;
  assign N7142 = N8630;
  assign N7143 = N8632;
  assign N7144 = N8634;
  assign N7145 = N8636;
  assign N7146 = N8638;
  assign N7147 = N8640;
  assign N7148 = N8642;
  assign N7149 = N8644;
  assign N7150 = N8646;
  assign N7151 = N8648;
  assign N7152 = N8650;
  assign N7153 = N8652;
  assign N7154 = N8654;
  assign N7155 = N8656;
  assign N7156 = N8658;
  assign N7157 = N8660;
  assign N7158 = N8662;
  assign N7159 = N8664;
  assign N7160 = N8666;
  assign N7161 = N8668;
  assign N7162 = N8670;
  assign N7163 = N8672;
  assign N7164 = N8674;
  assign N7165 = N8676;
  assign N7166 = N8678;
  assign N7167 = N8680;
  assign N7168 = N8682;
  assign N7169 = N8684;
  assign N7170 = N8686;
  assign N7171 = N8688;
  assign N7172 = N8690;
  assign N7173 = N8692;
  assign N7174 = N8694;
  assign N7175 = N8696;
  assign way_id_o[6] = (N7301)? lru_i[0] : 
                       (N7303)? lru_i[1] : 
                       (N7305)? lru_i[2] : 
                       (N7307)? lru_i[3] : 
                       (N7309)? lru_i[4] : 
                       (N7311)? lru_i[5] : 
                       (N7313)? lru_i[6] : 
                       (N7315)? lru_i[7] : 
                       (N7317)? lru_i[8] : 
                       (N7319)? lru_i[9] : 
                       (N7321)? lru_i[10] : 
                       (N7323)? lru_i[11] : 
                       (N7325)? lru_i[12] : 
                       (N7327)? lru_i[13] : 
                       (N7329)? lru_i[14] : 
                       (N7331)? lru_i[15] : 
                       (N7333)? lru_i[16] : 
                       (N7335)? lru_i[17] : 
                       (N7337)? lru_i[18] : 
                       (N7339)? lru_i[19] : 
                       (N7341)? lru_i[20] : 
                       (N7343)? lru_i[21] : 
                       (N7345)? lru_i[22] : 
                       (N7347)? lru_i[23] : 
                       (N7349)? lru_i[24] : 
                       (N7351)? lru_i[25] : 
                       (N7353)? lru_i[26] : 
                       (N7355)? lru_i[27] : 
                       (N7357)? lru_i[28] : 
                       (N7359)? lru_i[29] : 
                       (N7361)? lru_i[30] : 
                       (N7363)? lru_i[31] : 
                       (N7365)? lru_i[32] : 
                       (N7367)? lru_i[33] : 
                       (N7369)? lru_i[34] : 
                       (N7371)? lru_i[35] : 
                       (N7373)? lru_i[36] : 
                       (N7375)? lru_i[37] : 
                       (N7377)? lru_i[38] : 
                       (N7379)? lru_i[39] : 
                       (N7381)? lru_i[40] : 
                       (N7383)? lru_i[41] : 
                       (N7385)? lru_i[42] : 
                       (N7387)? lru_i[43] : 
                       (N7389)? lru_i[44] : 
                       (N7391)? lru_i[45] : 
                       (N7393)? lru_i[46] : 
                       (N7395)? lru_i[47] : 
                       (N7397)? lru_i[48] : 
                       (N7399)? lru_i[49] : 
                       (N7401)? lru_i[50] : 
                       (N7403)? lru_i[51] : 
                       (N7405)? lru_i[52] : 
                       (N7407)? lru_i[53] : 
                       (N7409)? lru_i[54] : 
                       (N7411)? lru_i[55] : 
                       (N7413)? lru_i[56] : 
                       (N7415)? lru_i[57] : 
                       (N7417)? lru_i[58] : 
                       (N7419)? lru_i[59] : 
                       (N7421)? lru_i[60] : 
                       (N7423)? lru_i[61] : 
                       (N7425)? lru_i[62] : 
                       (N7427)? lru_i[63] : 
                       (N7302)? lru_i[64] : 
                       (N7304)? lru_i[65] : 
                       (N7306)? lru_i[66] : 
                       (N7308)? lru_i[67] : 
                       (N7310)? lru_i[68] : 
                       (N7312)? lru_i[69] : 
                       (N7314)? lru_i[70] : 
                       (N7316)? lru_i[71] : 
                       (N7318)? lru_i[72] : 
                       (N7320)? lru_i[73] : 
                       (N7322)? lru_i[74] : 
                       (N7324)? lru_i[75] : 
                       (N7326)? lru_i[76] : 
                       (N7328)? lru_i[77] : 
                       (N7330)? lru_i[78] : 
                       (N7332)? lru_i[79] : 
                       (N7334)? lru_i[80] : 
                       (N7336)? lru_i[81] : 
                       (N7338)? lru_i[82] : 
                       (N7340)? lru_i[83] : 
                       (N7342)? lru_i[84] : 
                       (N7344)? lru_i[85] : 
                       (N7346)? lru_i[86] : 
                       (N7348)? lru_i[87] : 
                       (N7350)? lru_i[88] : 
                       (N7352)? lru_i[89] : 
                       (N7354)? lru_i[90] : 
                       (N7356)? lru_i[91] : 
                       (N7358)? lru_i[92] : 
                       (N7360)? lru_i[93] : 
                       (N7362)? lru_i[94] : 
                       (N7364)? lru_i[95] : 
                       (N7366)? lru_i[96] : 
                       (N7368)? lru_i[97] : 
                       (N7370)? lru_i[98] : 
                       (N7372)? lru_i[99] : 
                       (N7374)? lru_i[100] : 
                       (N7376)? lru_i[101] : 
                       (N7378)? lru_i[102] : 
                       (N7380)? lru_i[103] : 
                       (N7382)? lru_i[104] : 
                       (N7384)? lru_i[105] : 
                       (N7386)? lru_i[106] : 
                       (N7388)? lru_i[107] : 
                       (N7390)? lru_i[108] : 
                       (N7392)? lru_i[109] : 
                       (N7394)? lru_i[110] : 
                       (N7396)? lru_i[111] : 
                       (N7398)? lru_i[112] : 
                       (N7400)? lru_i[113] : 
                       (N7402)? lru_i[114] : 
                       (N7404)? lru_i[115] : 
                       (N7406)? lru_i[116] : 
                       (N7408)? lru_i[117] : 
                       (N7410)? lru_i[118] : 
                       (N7412)? lru_i[119] : 
                       (N7414)? lru_i[120] : 
                       (N7416)? lru_i[121] : 
                       (N7418)? lru_i[122] : 
                       (N7420)? lru_i[123] : 
                       (N7422)? lru_i[124] : 
                       (N7424)? lru_i[125] : 
                       (N7426)? lru_i[126] : 1'b0;
  assign mask[1] = 1'b1 & N8825;
  assign N8825 = ~lru_i[0];
  assign mask[2] = 1'b1 & lru_i[0];
  assign mask[3] = mask[1] & N8826;
  assign N8826 = ~lru_i[1];
  assign mask[4] = mask[1] & lru_i[1];
  assign mask[5] = mask[2] & N8827;
  assign N8827 = ~lru_i[2];
  assign mask[6] = mask[2] & lru_i[2];
  assign mask[7] = mask[3] & N8828;
  assign N8828 = ~lru_i[3];
  assign mask[8] = mask[3] & lru_i[3];
  assign mask[9] = mask[4] & N8829;
  assign N8829 = ~lru_i[4];
  assign mask[10] = mask[4] & lru_i[4];
  assign mask[11] = mask[5] & N8830;
  assign N8830 = ~lru_i[5];
  assign mask[12] = mask[5] & lru_i[5];
  assign mask[13] = mask[6] & N8831;
  assign N8831 = ~lru_i[6];
  assign mask[14] = mask[6] & lru_i[6];
  assign mask[15] = mask[7] & N8832;
  assign N8832 = ~lru_i[7];
  assign mask[16] = mask[7] & lru_i[7];
  assign mask[17] = mask[8] & N8833;
  assign N8833 = ~lru_i[8];
  assign mask[18] = mask[8] & lru_i[8];
  assign mask[19] = mask[9] & N8834;
  assign N8834 = ~lru_i[9];
  assign mask[20] = mask[9] & lru_i[9];
  assign mask[21] = mask[10] & N8835;
  assign N8835 = ~lru_i[10];
  assign mask[22] = mask[10] & lru_i[10];
  assign mask[23] = mask[11] & N8836;
  assign N8836 = ~lru_i[11];
  assign mask[24] = mask[11] & lru_i[11];
  assign mask[25] = mask[12] & N8837;
  assign N8837 = ~lru_i[12];
  assign mask[26] = mask[12] & lru_i[12];
  assign mask[27] = mask[13] & N8838;
  assign N8838 = ~lru_i[13];
  assign mask[28] = mask[13] & lru_i[13];
  assign mask[29] = mask[14] & N8839;
  assign N8839 = ~lru_i[14];
  assign mask[30] = mask[14] & lru_i[14];
  assign mask[31] = mask[15] & N8840;
  assign N8840 = ~lru_i[15];
  assign mask[32] = mask[15] & lru_i[15];
  assign mask[33] = mask[16] & N8841;
  assign N8841 = ~lru_i[16];
  assign mask[34] = mask[16] & lru_i[16];
  assign mask[35] = mask[17] & N8842;
  assign N8842 = ~lru_i[17];
  assign mask[36] = mask[17] & lru_i[17];
  assign mask[37] = mask[18] & N8843;
  assign N8843 = ~lru_i[18];
  assign mask[38] = mask[18] & lru_i[18];
  assign mask[39] = mask[19] & N8844;
  assign N8844 = ~lru_i[19];
  assign mask[40] = mask[19] & lru_i[19];
  assign mask[41] = mask[20] & N8845;
  assign N8845 = ~lru_i[20];
  assign mask[42] = mask[20] & lru_i[20];
  assign mask[43] = mask[21] & N8846;
  assign N8846 = ~lru_i[21];
  assign mask[44] = mask[21] & lru_i[21];
  assign mask[45] = mask[22] & N8847;
  assign N8847 = ~lru_i[22];
  assign mask[46] = mask[22] & lru_i[22];
  assign mask[47] = mask[23] & N8848;
  assign N8848 = ~lru_i[23];
  assign mask[48] = mask[23] & lru_i[23];
  assign mask[49] = mask[24] & N8849;
  assign N8849 = ~lru_i[24];
  assign mask[50] = mask[24] & lru_i[24];
  assign mask[51] = mask[25] & N8850;
  assign N8850 = ~lru_i[25];
  assign mask[52] = mask[25] & lru_i[25];
  assign mask[53] = mask[26] & N8851;
  assign N8851 = ~lru_i[26];
  assign mask[54] = mask[26] & lru_i[26];
  assign mask[55] = mask[27] & N8852;
  assign N8852 = ~lru_i[27];
  assign mask[56] = mask[27] & lru_i[27];
  assign mask[57] = mask[28] & N8853;
  assign N8853 = ~lru_i[28];
  assign mask[58] = mask[28] & lru_i[28];
  assign mask[59] = mask[29] & N8854;
  assign N8854 = ~lru_i[29];
  assign mask[60] = mask[29] & lru_i[29];
  assign mask[61] = mask[30] & N8855;
  assign N8855 = ~lru_i[30];
  assign mask[62] = mask[30] & lru_i[30];
  assign mask[63] = mask[31] & N8856;
  assign N8856 = ~lru_i[31];
  assign mask[64] = mask[31] & lru_i[31];
  assign mask[65] = mask[32] & N8857;
  assign N8857 = ~lru_i[32];
  assign mask[66] = mask[32] & lru_i[32];
  assign mask[67] = mask[33] & N8858;
  assign N8858 = ~lru_i[33];
  assign mask[68] = mask[33] & lru_i[33];
  assign mask[69] = mask[34] & N8859;
  assign N8859 = ~lru_i[34];
  assign mask[70] = mask[34] & lru_i[34];
  assign mask[71] = mask[35] & N8860;
  assign N8860 = ~lru_i[35];
  assign mask[72] = mask[35] & lru_i[35];
  assign mask[73] = mask[36] & N8861;
  assign N8861 = ~lru_i[36];
  assign mask[74] = mask[36] & lru_i[36];
  assign mask[75] = mask[37] & N8862;
  assign N8862 = ~lru_i[37];
  assign mask[76] = mask[37] & lru_i[37];
  assign mask[77] = mask[38] & N8863;
  assign N8863 = ~lru_i[38];
  assign mask[78] = mask[38] & lru_i[38];
  assign mask[79] = mask[39] & N8864;
  assign N8864 = ~lru_i[39];
  assign mask[80] = mask[39] & lru_i[39];
  assign mask[81] = mask[40] & N8865;
  assign N8865 = ~lru_i[40];
  assign mask[82] = mask[40] & lru_i[40];
  assign mask[83] = mask[41] & N8866;
  assign N8866 = ~lru_i[41];
  assign mask[84] = mask[41] & lru_i[41];
  assign mask[85] = mask[42] & N8867;
  assign N8867 = ~lru_i[42];
  assign mask[86] = mask[42] & lru_i[42];
  assign mask[87] = mask[43] & N8868;
  assign N8868 = ~lru_i[43];
  assign mask[88] = mask[43] & lru_i[43];
  assign mask[89] = mask[44] & N8869;
  assign N8869 = ~lru_i[44];
  assign mask[90] = mask[44] & lru_i[44];
  assign mask[91] = mask[45] & N8870;
  assign N8870 = ~lru_i[45];
  assign mask[92] = mask[45] & lru_i[45];
  assign mask[93] = mask[46] & N8871;
  assign N8871 = ~lru_i[46];
  assign mask[94] = mask[46] & lru_i[46];
  assign mask[95] = mask[47] & N8872;
  assign N8872 = ~lru_i[47];
  assign mask[96] = mask[47] & lru_i[47];
  assign mask[97] = mask[48] & N8873;
  assign N8873 = ~lru_i[48];
  assign mask[98] = mask[48] & lru_i[48];
  assign mask[99] = mask[49] & N8874;
  assign N8874 = ~lru_i[49];
  assign mask[100] = mask[49] & lru_i[49];
  assign mask[101] = mask[50] & N8875;
  assign N8875 = ~lru_i[50];
  assign mask[102] = mask[50] & lru_i[50];
  assign mask[103] = mask[51] & N8876;
  assign N8876 = ~lru_i[51];
  assign mask[104] = mask[51] & lru_i[51];
  assign mask[105] = mask[52] & N8877;
  assign N8877 = ~lru_i[52];
  assign mask[106] = mask[52] & lru_i[52];
  assign mask[107] = mask[53] & N8878;
  assign N8878 = ~lru_i[53];
  assign mask[108] = mask[53] & lru_i[53];
  assign mask[109] = mask[54] & N8879;
  assign N8879 = ~lru_i[54];
  assign mask[110] = mask[54] & lru_i[54];
  assign mask[111] = mask[55] & N8880;
  assign N8880 = ~lru_i[55];
  assign mask[112] = mask[55] & lru_i[55];
  assign mask[113] = mask[56] & N8881;
  assign N8881 = ~lru_i[56];
  assign mask[114] = mask[56] & lru_i[56];
  assign mask[115] = mask[57] & N8882;
  assign N8882 = ~lru_i[57];
  assign mask[116] = mask[57] & lru_i[57];
  assign mask[117] = mask[58] & N8883;
  assign N8883 = ~lru_i[58];
  assign mask[118] = mask[58] & lru_i[58];
  assign mask[119] = mask[59] & N8884;
  assign N8884 = ~lru_i[59];
  assign mask[120] = mask[59] & lru_i[59];
  assign mask[121] = mask[60] & N8885;
  assign N8885 = ~lru_i[60];
  assign mask[122] = mask[60] & lru_i[60];
  assign mask[123] = mask[61] & N8886;
  assign N8886 = ~lru_i[61];
  assign mask[124] = mask[61] & lru_i[61];
  assign mask[125] = mask[62] & N8887;
  assign N8887 = ~lru_i[62];
  assign mask[126] = mask[62] & lru_i[62];
  assign N7176 = N7236 & N7236;
  assign N7177 = N7236 & 1'b0;
  assign N7178 = 1'b0 & N7236;
  assign N7179 = 1'b0 & 1'b0;
  assign N7180 = N7176 & N7236;
  assign N7181 = N7176 & 1'b0;
  assign N7182 = N7178 & N7236;
  assign N7183 = N7178 & 1'b0;
  assign N7184 = N7177 & N7236;
  assign N7185 = N7177 & 1'b0;
  assign N7186 = N7179 & N7236;
  assign N7187 = N7179 & 1'b0;
  assign N7188 = N7180 & N7236;
  assign N7189 = N7180 & 1'b0;
  assign N7190 = N7182 & N7236;
  assign N7191 = N7182 & 1'b0;
  assign N7192 = N7184 & N7236;
  assign N7193 = N7184 & 1'b0;
  assign N7194 = N7186 & N7236;
  assign N7195 = N7186 & 1'b0;
  assign N7196 = N7181 & N7236;
  assign N7197 = N7181 & 1'b0;
  assign N7198 = N7183 & N7236;
  assign N7199 = N7183 & 1'b0;
  assign N7200 = N7185 & N7236;
  assign N7201 = N7185 & 1'b0;
  assign N7202 = N7187 & N7236;
  assign N7203 = N7187 & 1'b0;
  assign N7204 = N7188 & N7236;
  assign N7205 = N7188 & 1'b0;
  assign N7206 = N7190 & N7236;
  assign N7207 = N7190 & 1'b0;
  assign N7208 = N7192 & N7236;
  assign N7209 = N7192 & 1'b0;
  assign N7210 = N7194 & N7236;
  assign N7211 = N7194 & 1'b0;
  assign N7212 = N7196 & N7236;
  assign N7213 = N7196 & 1'b0;
  assign N7214 = N7198 & N7236;
  assign N7215 = N7198 & 1'b0;
  assign N7216 = N7200 & N7236;
  assign N7217 = N7200 & 1'b0;
  assign N7218 = N7202 & N7236;
  assign N7219 = N7202 & 1'b0;
  assign N7220 = N7189 & N7236;
  assign N7221 = N7189 & 1'b0;
  assign N7222 = N7191 & N7236;
  assign N7223 = N7191 & 1'b0;
  assign N7224 = N7193 & N7236;
  assign N7225 = N7193 & 1'b0;
  assign N7226 = N7195 & N7236;
  assign N7227 = N7195 & 1'b0;
  assign N7228 = N7197 & N7236;
  assign N7229 = N7197 & 1'b0;
  assign N7230 = N7199 & N7236;
  assign N7231 = N7199 & 1'b0;
  assign N7232 = N7201 & N7236;
  assign N7233 = N7201 & 1'b0;
  assign N7234 = N7203 & N7236;
  assign N7235 = N7203 & 1'b0;
  assign N7236 = ~1'b0;
  assign N7237 = N7204 & N7236;
  assign N7238 = N7204 & 1'b0;
  assign N7239 = N7206 & N7236;
  assign N7240 = N7206 & 1'b0;
  assign N7241 = N7208 & N7236;
  assign N7242 = N7208 & 1'b0;
  assign N7243 = N7210 & N7236;
  assign N7244 = N7210 & 1'b0;
  assign N7245 = N7212 & N7236;
  assign N7246 = N7212 & 1'b0;
  assign N7247 = N7214 & N7236;
  assign N7248 = N7214 & 1'b0;
  assign N7249 = N7216 & N7236;
  assign N7250 = N7216 & 1'b0;
  assign N7251 = N7218 & N7236;
  assign N7252 = N7218 & 1'b0;
  assign N7253 = N7220 & N7236;
  assign N7254 = N7220 & 1'b0;
  assign N7255 = N7222 & N7236;
  assign N7256 = N7222 & 1'b0;
  assign N7257 = N7224 & N7236;
  assign N7258 = N7224 & 1'b0;
  assign N7259 = N7226 & N7236;
  assign N7260 = N7226 & 1'b0;
  assign N7261 = N7228 & N7236;
  assign N7262 = N7228 & 1'b0;
  assign N7263 = N7230 & N7236;
  assign N7264 = N7230 & 1'b0;
  assign N7265 = N7232 & N7236;
  assign N7266 = N7232 & 1'b0;
  assign N7267 = N7234 & N7236;
  assign N7268 = N7234 & 1'b0;
  assign N7269 = N7205 & N7236;
  assign N7270 = N7205 & 1'b0;
  assign N7271 = N7207 & N7236;
  assign N7272 = N7207 & 1'b0;
  assign N7273 = N7209 & N7236;
  assign N7274 = N7209 & 1'b0;
  assign N7275 = N7211 & N7236;
  assign N7276 = N7211 & 1'b0;
  assign N7277 = N7213 & N7236;
  assign N7278 = N7213 & 1'b0;
  assign N7279 = N7215 & N7236;
  assign N7280 = N7215 & 1'b0;
  assign N7281 = N7217 & N7236;
  assign N7282 = N7217 & 1'b0;
  assign N7283 = N7219 & N7236;
  assign N7284 = N7219 & 1'b0;
  assign N7285 = N7221 & N7236;
  assign N7286 = N7221 & 1'b0;
  assign N7287 = N7223 & N7236;
  assign N7288 = N7223 & 1'b0;
  assign N7289 = N7225 & N7236;
  assign N7290 = N7225 & 1'b0;
  assign N7291 = N7227 & N7236;
  assign N7292 = N7227 & 1'b0;
  assign N7293 = N7229 & N7236;
  assign N7294 = N7229 & 1'b0;
  assign N7295 = N7231 & N7236;
  assign N7296 = N7231 & 1'b0;
  assign N7297 = N7233 & N7236;
  assign N7298 = N7233 & 1'b0;
  assign N7299 = N7235 & N7236;
  assign N7300 = N7235 & 1'b0;
  assign N7301 = N7237 & N7236;
  assign N7302 = N7237 & 1'b0;
  assign N7303 = N7239 & N7236;
  assign N7304 = N7239 & 1'b0;
  assign N7305 = N7241 & N7236;
  assign N7306 = N7241 & 1'b0;
  assign N7307 = N7243 & N7236;
  assign N7308 = N7243 & 1'b0;
  assign N7309 = N7245 & N7236;
  assign N7310 = N7245 & 1'b0;
  assign N7311 = N7247 & N7236;
  assign N7312 = N7247 & 1'b0;
  assign N7313 = N7249 & N7236;
  assign N7314 = N7249 & 1'b0;
  assign N7315 = N7251 & N7236;
  assign N7316 = N7251 & 1'b0;
  assign N7317 = N7253 & N7236;
  assign N7318 = N7253 & 1'b0;
  assign N7319 = N7255 & N7236;
  assign N7320 = N7255 & 1'b0;
  assign N7321 = N7257 & N7236;
  assign N7322 = N7257 & 1'b0;
  assign N7323 = N7259 & N7236;
  assign N7324 = N7259 & 1'b0;
  assign N7325 = N7261 & N7236;
  assign N7326 = N7261 & 1'b0;
  assign N7327 = N7263 & N7236;
  assign N7328 = N7263 & 1'b0;
  assign N7329 = N7265 & N7236;
  assign N7330 = N7265 & 1'b0;
  assign N7331 = N7267 & N7236;
  assign N7332 = N7267 & 1'b0;
  assign N7333 = N7269 & N7236;
  assign N7334 = N7269 & 1'b0;
  assign N7335 = N7271 & N7236;
  assign N7336 = N7271 & 1'b0;
  assign N7337 = N7273 & N7236;
  assign N7338 = N7273 & 1'b0;
  assign N7339 = N7275 & N7236;
  assign N7340 = N7275 & 1'b0;
  assign N7341 = N7277 & N7236;
  assign N7342 = N7277 & 1'b0;
  assign N7343 = N7279 & N7236;
  assign N7344 = N7279 & 1'b0;
  assign N7345 = N7281 & N7236;
  assign N7346 = N7281 & 1'b0;
  assign N7347 = N7283 & N7236;
  assign N7348 = N7283 & 1'b0;
  assign N7349 = N7285 & N7236;
  assign N7350 = N7285 & 1'b0;
  assign N7351 = N7287 & N7236;
  assign N7352 = N7287 & 1'b0;
  assign N7353 = N7289 & N7236;
  assign N7354 = N7289 & 1'b0;
  assign N7355 = N7291 & N7236;
  assign N7356 = N7291 & 1'b0;
  assign N7357 = N7293 & N7236;
  assign N7358 = N7293 & 1'b0;
  assign N7359 = N7295 & N7236;
  assign N7360 = N7295 & 1'b0;
  assign N7361 = N7297 & N7236;
  assign N7362 = N7297 & 1'b0;
  assign N7363 = N7299 & N7236;
  assign N7364 = N7299 & 1'b0;
  assign N7365 = N7238 & N7236;
  assign N7366 = N7238 & 1'b0;
  assign N7367 = N7240 & N7236;
  assign N7368 = N7240 & 1'b0;
  assign N7369 = N7242 & N7236;
  assign N7370 = N7242 & 1'b0;
  assign N7371 = N7244 & N7236;
  assign N7372 = N7244 & 1'b0;
  assign N7373 = N7246 & N7236;
  assign N7374 = N7246 & 1'b0;
  assign N7375 = N7248 & N7236;
  assign N7376 = N7248 & 1'b0;
  assign N7377 = N7250 & N7236;
  assign N7378 = N7250 & 1'b0;
  assign N7379 = N7252 & N7236;
  assign N7380 = N7252 & 1'b0;
  assign N7381 = N7254 & N7236;
  assign N7382 = N7254 & 1'b0;
  assign N7383 = N7256 & N7236;
  assign N7384 = N7256 & 1'b0;
  assign N7385 = N7258 & N7236;
  assign N7386 = N7258 & 1'b0;
  assign N7387 = N7260 & N7236;
  assign N7388 = N7260 & 1'b0;
  assign N7389 = N7262 & N7236;
  assign N7390 = N7262 & 1'b0;
  assign N7391 = N7264 & N7236;
  assign N7392 = N7264 & 1'b0;
  assign N7393 = N7266 & N7236;
  assign N7394 = N7266 & 1'b0;
  assign N7395 = N7268 & N7236;
  assign N7396 = N7268 & 1'b0;
  assign N7397 = N7270 & N7236;
  assign N7398 = N7270 & 1'b0;
  assign N7399 = N7272 & N7236;
  assign N7400 = N7272 & 1'b0;
  assign N7401 = N7274 & N7236;
  assign N7402 = N7274 & 1'b0;
  assign N7403 = N7276 & N7236;
  assign N7404 = N7276 & 1'b0;
  assign N7405 = N7278 & N7236;
  assign N7406 = N7278 & 1'b0;
  assign N7407 = N7280 & N7236;
  assign N7408 = N7280 & 1'b0;
  assign N7409 = N7282 & N7236;
  assign N7410 = N7282 & 1'b0;
  assign N7411 = N7284 & N7236;
  assign N7412 = N7284 & 1'b0;
  assign N7413 = N7286 & N7236;
  assign N7414 = N7286 & 1'b0;
  assign N7415 = N7288 & N7236;
  assign N7416 = N7288 & 1'b0;
  assign N7417 = N7290 & N7236;
  assign N7418 = N7290 & 1'b0;
  assign N7419 = N7292 & N7236;
  assign N7420 = N7292 & 1'b0;
  assign N7421 = N7294 & N7236;
  assign N7422 = N7294 & 1'b0;
  assign N7423 = N7296 & N7236;
  assign N7424 = N7296 & 1'b0;
  assign N7425 = N7298 & N7236;
  assign N7426 = N7298 & 1'b0;
  assign N7427 = N7300 & N7236;
  assign pe_i_1__126_ = mask[126] ^ 1'b0;
  assign pe_i_1__125_ = mask[125] ^ 1'b0;
  assign pe_i_1__124_ = mask[124] ^ 1'b0;
  assign pe_i_1__123_ = mask[123] ^ 1'b0;
  assign pe_i_1__122_ = mask[122] ^ 1'b0;
  assign pe_i_1__121_ = mask[121] ^ 1'b0;
  assign pe_i_1__120_ = mask[120] ^ 1'b0;
  assign pe_i_1__119_ = mask[119] ^ 1'b0;
  assign pe_i_1__118_ = mask[118] ^ 1'b0;
  assign pe_i_1__117_ = mask[117] ^ 1'b0;
  assign pe_i_1__116_ = mask[116] ^ 1'b0;
  assign pe_i_1__115_ = mask[115] ^ 1'b0;
  assign pe_i_1__114_ = mask[114] ^ 1'b0;
  assign pe_i_1__113_ = mask[113] ^ 1'b0;
  assign pe_i_1__112_ = mask[112] ^ 1'b0;
  assign pe_i_1__111_ = mask[111] ^ 1'b0;
  assign pe_i_1__110_ = mask[110] ^ 1'b0;
  assign pe_i_1__109_ = mask[109] ^ 1'b0;
  assign pe_i_1__108_ = mask[108] ^ 1'b0;
  assign pe_i_1__107_ = mask[107] ^ 1'b0;
  assign pe_i_1__106_ = mask[106] ^ 1'b0;
  assign pe_i_1__105_ = mask[105] ^ 1'b0;
  assign pe_i_1__104_ = mask[104] ^ 1'b0;
  assign pe_i_1__103_ = mask[103] ^ 1'b0;
  assign pe_i_1__102_ = mask[102] ^ 1'b0;
  assign pe_i_1__101_ = mask[101] ^ 1'b0;
  assign pe_i_1__100_ = mask[100] ^ 1'b0;
  assign pe_i_1__99_ = mask[99] ^ 1'b0;
  assign pe_i_1__98_ = mask[98] ^ 1'b0;
  assign pe_i_1__97_ = mask[97] ^ 1'b0;
  assign pe_i_1__96_ = mask[96] ^ 1'b0;
  assign pe_i_1__95_ = mask[95] ^ 1'b0;
  assign pe_i_1__94_ = mask[94] ^ 1'b0;
  assign pe_i_1__93_ = mask[93] ^ 1'b0;
  assign pe_i_1__92_ = mask[92] ^ 1'b0;
  assign pe_i_1__91_ = mask[91] ^ 1'b0;
  assign pe_i_1__90_ = mask[90] ^ 1'b0;
  assign pe_i_1__89_ = mask[89] ^ 1'b0;
  assign pe_i_1__88_ = mask[88] ^ 1'b0;
  assign pe_i_1__87_ = mask[87] ^ 1'b0;
  assign pe_i_1__86_ = mask[86] ^ 1'b0;
  assign pe_i_1__85_ = mask[85] ^ 1'b0;
  assign pe_i_1__84_ = mask[84] ^ 1'b0;
  assign pe_i_1__83_ = mask[83] ^ 1'b0;
  assign pe_i_1__82_ = mask[82] ^ 1'b0;
  assign pe_i_1__81_ = mask[81] ^ 1'b0;
  assign pe_i_1__80_ = mask[80] ^ 1'b0;
  assign pe_i_1__79_ = mask[79] ^ 1'b0;
  assign pe_i_1__78_ = mask[78] ^ 1'b0;
  assign pe_i_1__77_ = mask[77] ^ 1'b0;
  assign pe_i_1__76_ = mask[76] ^ 1'b0;
  assign pe_i_1__75_ = mask[75] ^ 1'b0;
  assign pe_i_1__74_ = mask[74] ^ 1'b0;
  assign pe_i_1__73_ = mask[73] ^ 1'b0;
  assign pe_i_1__72_ = mask[72] ^ 1'b0;
  assign pe_i_1__71_ = mask[71] ^ 1'b0;
  assign pe_i_1__70_ = mask[70] ^ 1'b0;
  assign pe_i_1__69_ = mask[69] ^ 1'b0;
  assign pe_i_1__68_ = mask[68] ^ 1'b0;
  assign pe_i_1__67_ = mask[67] ^ 1'b0;
  assign pe_i_1__66_ = mask[66] ^ 1'b0;
  assign pe_i_1__65_ = mask[65] ^ 1'b0;
  assign pe_i_1__64_ = mask[64] ^ 1'b0;
  assign pe_i_1__63_ = mask[63] ^ 1'b0;
  assign pe_i_1__62_ = mask[62] ^ 1'b0;
  assign pe_i_1__61_ = mask[61] ^ 1'b0;
  assign pe_i_1__60_ = mask[60] ^ 1'b0;
  assign pe_i_1__59_ = mask[59] ^ 1'b0;
  assign pe_i_1__58_ = mask[58] ^ 1'b0;
  assign pe_i_1__57_ = mask[57] ^ 1'b0;
  assign pe_i_1__56_ = mask[56] ^ 1'b0;
  assign pe_i_1__55_ = mask[55] ^ 1'b0;
  assign pe_i_1__54_ = mask[54] ^ 1'b0;
  assign pe_i_1__53_ = mask[53] ^ 1'b0;
  assign pe_i_1__52_ = mask[52] ^ 1'b0;
  assign pe_i_1__51_ = mask[51] ^ 1'b0;
  assign pe_i_1__50_ = mask[50] ^ 1'b0;
  assign pe_i_1__49_ = mask[49] ^ 1'b0;
  assign pe_i_1__48_ = mask[48] ^ 1'b0;
  assign pe_i_1__47_ = mask[47] ^ 1'b0;
  assign pe_i_1__46_ = mask[46] ^ 1'b0;
  assign pe_i_1__45_ = mask[45] ^ 1'b0;
  assign pe_i_1__44_ = mask[44] ^ 1'b0;
  assign pe_i_1__43_ = mask[43] ^ 1'b0;
  assign pe_i_1__42_ = mask[42] ^ 1'b0;
  assign pe_i_1__41_ = mask[41] ^ 1'b0;
  assign pe_i_1__40_ = mask[40] ^ 1'b0;
  assign pe_i_1__39_ = mask[39] ^ 1'b0;
  assign pe_i_1__38_ = mask[38] ^ 1'b0;
  assign pe_i_1__37_ = mask[37] ^ 1'b0;
  assign pe_i_1__36_ = mask[36] ^ 1'b0;
  assign pe_i_1__35_ = mask[35] ^ 1'b0;
  assign pe_i_1__34_ = mask[34] ^ 1'b0;
  assign pe_i_1__33_ = mask[33] ^ 1'b0;
  assign pe_i_1__32_ = mask[32] ^ 1'b0;
  assign pe_i_1__31_ = mask[31] ^ 1'b0;
  assign pe_i_1__30_ = mask[30] ^ 1'b0;
  assign pe_i_1__29_ = mask[29] ^ 1'b0;
  assign pe_i_1__28_ = mask[28] ^ 1'b0;
  assign pe_i_1__27_ = mask[27] ^ 1'b0;
  assign pe_i_1__26_ = mask[26] ^ 1'b0;
  assign pe_i_1__25_ = mask[25] ^ 1'b0;
  assign pe_i_1__24_ = mask[24] ^ 1'b0;
  assign pe_i_1__23_ = mask[23] ^ 1'b0;
  assign pe_i_1__22_ = mask[22] ^ 1'b0;
  assign pe_i_1__21_ = mask[21] ^ 1'b0;
  assign pe_i_1__20_ = mask[20] ^ 1'b0;
  assign pe_i_1__19_ = mask[19] ^ 1'b0;
  assign pe_i_1__18_ = mask[18] ^ 1'b0;
  assign pe_i_1__17_ = mask[17] ^ 1'b0;
  assign pe_i_1__16_ = mask[16] ^ 1'b0;
  assign pe_i_1__15_ = mask[15] ^ 1'b0;
  assign pe_i_1__14_ = mask[14] ^ 1'b0;
  assign pe_i_1__13_ = mask[13] ^ 1'b0;
  assign pe_i_1__12_ = mask[12] ^ 1'b0;
  assign pe_i_1__11_ = mask[11] ^ 1'b0;
  assign pe_i_1__10_ = mask[10] ^ 1'b0;
  assign pe_i_1__9_ = mask[9] ^ 1'b0;
  assign pe_i_1__8_ = mask[8] ^ 1'b0;
  assign pe_i_1__7_ = mask[7] ^ 1'b0;
  assign pe_i_1__6_ = mask[6] ^ 1'b0;
  assign pe_i_1__5_ = mask[5] ^ 1'b0;
  assign pe_i_1__4_ = mask[4] ^ 1'b0;
  assign pe_i_1__3_ = mask[3] ^ 1'b0;
  assign pe_i_1__2_ = mask[2] ^ 1'b0;
  assign pe_i_1__1_ = mask[1] ^ 1'b0;
  assign pe_i_1__0_ = 1'b1 ^ 1'b1;
  assign pe_i_2__126_ = pe_i_1__126_ ^ N7808;
  assign pe_i_2__125_ = pe_i_1__125_ ^ N7807;
  assign pe_i_2__124_ = pe_i_1__124_ ^ N7806;
  assign pe_i_2__123_ = pe_i_1__123_ ^ N7805;
  assign pe_i_2__122_ = pe_i_1__122_ ^ N7804;
  assign pe_i_2__121_ = pe_i_1__121_ ^ N7803;
  assign pe_i_2__120_ = pe_i_1__120_ ^ N7802;
  assign pe_i_2__119_ = pe_i_1__119_ ^ N7801;
  assign pe_i_2__118_ = pe_i_1__118_ ^ N7800;
  assign pe_i_2__117_ = pe_i_1__117_ ^ N7799;
  assign pe_i_2__116_ = pe_i_1__116_ ^ N7798;
  assign pe_i_2__115_ = pe_i_1__115_ ^ N7797;
  assign pe_i_2__114_ = pe_i_1__114_ ^ N7796;
  assign pe_i_2__113_ = pe_i_1__113_ ^ N7795;
  assign pe_i_2__112_ = pe_i_1__112_ ^ N7794;
  assign pe_i_2__111_ = pe_i_1__111_ ^ N7793;
  assign pe_i_2__110_ = pe_i_1__110_ ^ N7792;
  assign pe_i_2__109_ = pe_i_1__109_ ^ N7791;
  assign pe_i_2__108_ = pe_i_1__108_ ^ N7790;
  assign pe_i_2__107_ = pe_i_1__107_ ^ N7789;
  assign pe_i_2__106_ = pe_i_1__106_ ^ N7788;
  assign pe_i_2__105_ = pe_i_1__105_ ^ N7787;
  assign pe_i_2__104_ = pe_i_1__104_ ^ N7786;
  assign pe_i_2__103_ = pe_i_1__103_ ^ N7785;
  assign pe_i_2__102_ = pe_i_1__102_ ^ N7784;
  assign pe_i_2__101_ = pe_i_1__101_ ^ N7783;
  assign pe_i_2__100_ = pe_i_1__100_ ^ N7782;
  assign pe_i_2__99_ = pe_i_1__99_ ^ N7781;
  assign pe_i_2__98_ = pe_i_1__98_ ^ N7780;
  assign pe_i_2__97_ = pe_i_1__97_ ^ N7779;
  assign pe_i_2__96_ = pe_i_1__96_ ^ N7778;
  assign pe_i_2__95_ = pe_i_1__95_ ^ N7777;
  assign pe_i_2__94_ = pe_i_1__94_ ^ N7776;
  assign pe_i_2__93_ = pe_i_1__93_ ^ N7775;
  assign pe_i_2__92_ = pe_i_1__92_ ^ N7774;
  assign pe_i_2__91_ = pe_i_1__91_ ^ N7773;
  assign pe_i_2__90_ = pe_i_1__90_ ^ N7772;
  assign pe_i_2__89_ = pe_i_1__89_ ^ N7771;
  assign pe_i_2__88_ = pe_i_1__88_ ^ N7770;
  assign pe_i_2__87_ = pe_i_1__87_ ^ N7769;
  assign pe_i_2__86_ = pe_i_1__86_ ^ N7768;
  assign pe_i_2__85_ = pe_i_1__85_ ^ N7767;
  assign pe_i_2__84_ = pe_i_1__84_ ^ N7766;
  assign pe_i_2__83_ = pe_i_1__83_ ^ N7765;
  assign pe_i_2__82_ = pe_i_1__82_ ^ N7764;
  assign pe_i_2__81_ = pe_i_1__81_ ^ N7763;
  assign pe_i_2__80_ = pe_i_1__80_ ^ N7762;
  assign pe_i_2__79_ = pe_i_1__79_ ^ N7761;
  assign pe_i_2__78_ = pe_i_1__78_ ^ N7760;
  assign pe_i_2__77_ = pe_i_1__77_ ^ N7759;
  assign pe_i_2__76_ = pe_i_1__76_ ^ N7758;
  assign pe_i_2__75_ = pe_i_1__75_ ^ N7757;
  assign pe_i_2__74_ = pe_i_1__74_ ^ N7756;
  assign pe_i_2__73_ = pe_i_1__73_ ^ N7755;
  assign pe_i_2__72_ = pe_i_1__72_ ^ N7754;
  assign pe_i_2__71_ = pe_i_1__71_ ^ N7753;
  assign pe_i_2__70_ = pe_i_1__70_ ^ N7752;
  assign pe_i_2__69_ = pe_i_1__69_ ^ N7751;
  assign pe_i_2__68_ = pe_i_1__68_ ^ N7750;
  assign pe_i_2__67_ = pe_i_1__67_ ^ N7749;
  assign pe_i_2__66_ = pe_i_1__66_ ^ N7748;
  assign pe_i_2__65_ = pe_i_1__65_ ^ N7747;
  assign pe_i_2__64_ = pe_i_1__64_ ^ N7746;
  assign pe_i_2__63_ = pe_i_1__63_ ^ N7745;
  assign pe_i_2__62_ = pe_i_1__62_ ^ N7744;
  assign pe_i_2__61_ = pe_i_1__61_ ^ N7743;
  assign pe_i_2__60_ = pe_i_1__60_ ^ N7742;
  assign pe_i_2__59_ = pe_i_1__59_ ^ N7741;
  assign pe_i_2__58_ = pe_i_1__58_ ^ N7740;
  assign pe_i_2__57_ = pe_i_1__57_ ^ N7739;
  assign pe_i_2__56_ = pe_i_1__56_ ^ N7738;
  assign pe_i_2__55_ = pe_i_1__55_ ^ N7737;
  assign pe_i_2__54_ = pe_i_1__54_ ^ N7736;
  assign pe_i_2__53_ = pe_i_1__53_ ^ N7735;
  assign pe_i_2__52_ = pe_i_1__52_ ^ N7734;
  assign pe_i_2__51_ = pe_i_1__51_ ^ N7733;
  assign pe_i_2__50_ = pe_i_1__50_ ^ N7732;
  assign pe_i_2__49_ = pe_i_1__49_ ^ N7731;
  assign pe_i_2__48_ = pe_i_1__48_ ^ N7730;
  assign pe_i_2__47_ = pe_i_1__47_ ^ N7729;
  assign pe_i_2__46_ = pe_i_1__46_ ^ N7728;
  assign pe_i_2__45_ = pe_i_1__45_ ^ N7727;
  assign pe_i_2__44_ = pe_i_1__44_ ^ N7726;
  assign pe_i_2__43_ = pe_i_1__43_ ^ N7725;
  assign pe_i_2__42_ = pe_i_1__42_ ^ N7724;
  assign pe_i_2__41_ = pe_i_1__41_ ^ N7723;
  assign pe_i_2__40_ = pe_i_1__40_ ^ N7722;
  assign pe_i_2__39_ = pe_i_1__39_ ^ N7721;
  assign pe_i_2__38_ = pe_i_1__38_ ^ N7720;
  assign pe_i_2__37_ = pe_i_1__37_ ^ N7719;
  assign pe_i_2__36_ = pe_i_1__36_ ^ N7718;
  assign pe_i_2__35_ = pe_i_1__35_ ^ N7717;
  assign pe_i_2__34_ = pe_i_1__34_ ^ N7716;
  assign pe_i_2__33_ = pe_i_1__33_ ^ N7715;
  assign pe_i_2__32_ = pe_i_1__32_ ^ N7714;
  assign pe_i_2__31_ = pe_i_1__31_ ^ N7713;
  assign pe_i_2__30_ = pe_i_1__30_ ^ N7712;
  assign pe_i_2__29_ = pe_i_1__29_ ^ N7711;
  assign pe_i_2__28_ = pe_i_1__28_ ^ N7710;
  assign pe_i_2__27_ = pe_i_1__27_ ^ N7709;
  assign pe_i_2__26_ = pe_i_1__26_ ^ N7708;
  assign pe_i_2__25_ = pe_i_1__25_ ^ N7707;
  assign pe_i_2__24_ = pe_i_1__24_ ^ N7706;
  assign pe_i_2__23_ = pe_i_1__23_ ^ N7705;
  assign pe_i_2__22_ = pe_i_1__22_ ^ N7704;
  assign pe_i_2__21_ = pe_i_1__21_ ^ N7703;
  assign pe_i_2__20_ = pe_i_1__20_ ^ N7702;
  assign pe_i_2__19_ = pe_i_1__19_ ^ N7701;
  assign pe_i_2__18_ = pe_i_1__18_ ^ N7700;
  assign pe_i_2__17_ = pe_i_1__17_ ^ N7699;
  assign pe_i_2__16_ = pe_i_1__16_ ^ N7698;
  assign pe_i_2__15_ = pe_i_1__15_ ^ N7697;
  assign pe_i_2__14_ = pe_i_1__14_ ^ N7696;
  assign pe_i_2__13_ = pe_i_1__13_ ^ N7695;
  assign pe_i_2__12_ = pe_i_1__12_ ^ N7694;
  assign pe_i_2__11_ = pe_i_1__11_ ^ N7693;
  assign pe_i_2__10_ = pe_i_1__10_ ^ N7692;
  assign pe_i_2__9_ = pe_i_1__9_ ^ N7691;
  assign pe_i_2__8_ = pe_i_1__8_ ^ N7690;
  assign pe_i_2__7_ = pe_i_1__7_ ^ N7689;
  assign pe_i_2__6_ = pe_i_1__6_ ^ N7688;
  assign pe_i_2__5_ = pe_i_1__5_ ^ N7687;
  assign pe_i_2__4_ = pe_i_1__4_ ^ N7686;
  assign pe_i_2__3_ = pe_i_1__3_ ^ N7685;
  assign pe_i_2__2_ = pe_i_1__2_ ^ N7684;
  assign pe_i_2__1_ = pe_i_1__1_ ^ N7683;
  assign pe_i_2__0_ = pe_i_1__0_ ^ N7682;
  assign pe_i_3__126_ = pe_i_2__126_ ^ N8062;
  assign pe_i_3__125_ = pe_i_2__125_ ^ N8061;
  assign pe_i_3__124_ = pe_i_2__124_ ^ N8060;
  assign pe_i_3__123_ = pe_i_2__123_ ^ N8059;
  assign pe_i_3__122_ = pe_i_2__122_ ^ N8058;
  assign pe_i_3__121_ = pe_i_2__121_ ^ N8057;
  assign pe_i_3__120_ = pe_i_2__120_ ^ N8056;
  assign pe_i_3__119_ = pe_i_2__119_ ^ N8055;
  assign pe_i_3__118_ = pe_i_2__118_ ^ N8054;
  assign pe_i_3__117_ = pe_i_2__117_ ^ N8053;
  assign pe_i_3__116_ = pe_i_2__116_ ^ N8052;
  assign pe_i_3__115_ = pe_i_2__115_ ^ N8051;
  assign pe_i_3__114_ = pe_i_2__114_ ^ N8050;
  assign pe_i_3__113_ = pe_i_2__113_ ^ N8049;
  assign pe_i_3__112_ = pe_i_2__112_ ^ N8048;
  assign pe_i_3__111_ = pe_i_2__111_ ^ N8047;
  assign pe_i_3__110_ = pe_i_2__110_ ^ N8046;
  assign pe_i_3__109_ = pe_i_2__109_ ^ N8045;
  assign pe_i_3__108_ = pe_i_2__108_ ^ N8044;
  assign pe_i_3__107_ = pe_i_2__107_ ^ N8043;
  assign pe_i_3__106_ = pe_i_2__106_ ^ N8042;
  assign pe_i_3__105_ = pe_i_2__105_ ^ N8041;
  assign pe_i_3__104_ = pe_i_2__104_ ^ N8040;
  assign pe_i_3__103_ = pe_i_2__103_ ^ N8039;
  assign pe_i_3__102_ = pe_i_2__102_ ^ N8038;
  assign pe_i_3__101_ = pe_i_2__101_ ^ N8037;
  assign pe_i_3__100_ = pe_i_2__100_ ^ N8036;
  assign pe_i_3__99_ = pe_i_2__99_ ^ N8035;
  assign pe_i_3__98_ = pe_i_2__98_ ^ N8034;
  assign pe_i_3__97_ = pe_i_2__97_ ^ N8033;
  assign pe_i_3__96_ = pe_i_2__96_ ^ N8032;
  assign pe_i_3__95_ = pe_i_2__95_ ^ N8031;
  assign pe_i_3__94_ = pe_i_2__94_ ^ N8030;
  assign pe_i_3__93_ = pe_i_2__93_ ^ N8029;
  assign pe_i_3__92_ = pe_i_2__92_ ^ N8028;
  assign pe_i_3__91_ = pe_i_2__91_ ^ N8027;
  assign pe_i_3__90_ = pe_i_2__90_ ^ N8026;
  assign pe_i_3__89_ = pe_i_2__89_ ^ N8025;
  assign pe_i_3__88_ = pe_i_2__88_ ^ N8024;
  assign pe_i_3__87_ = pe_i_2__87_ ^ N8023;
  assign pe_i_3__86_ = pe_i_2__86_ ^ N8022;
  assign pe_i_3__85_ = pe_i_2__85_ ^ N8021;
  assign pe_i_3__84_ = pe_i_2__84_ ^ N8020;
  assign pe_i_3__83_ = pe_i_2__83_ ^ N8019;
  assign pe_i_3__82_ = pe_i_2__82_ ^ N8018;
  assign pe_i_3__81_ = pe_i_2__81_ ^ N8017;
  assign pe_i_3__80_ = pe_i_2__80_ ^ N8016;
  assign pe_i_3__79_ = pe_i_2__79_ ^ N8015;
  assign pe_i_3__78_ = pe_i_2__78_ ^ N8014;
  assign pe_i_3__77_ = pe_i_2__77_ ^ N8013;
  assign pe_i_3__76_ = pe_i_2__76_ ^ N8012;
  assign pe_i_3__75_ = pe_i_2__75_ ^ N8011;
  assign pe_i_3__74_ = pe_i_2__74_ ^ N8010;
  assign pe_i_3__73_ = pe_i_2__73_ ^ N8009;
  assign pe_i_3__72_ = pe_i_2__72_ ^ N8008;
  assign pe_i_3__71_ = pe_i_2__71_ ^ N8007;
  assign pe_i_3__70_ = pe_i_2__70_ ^ N8006;
  assign pe_i_3__69_ = pe_i_2__69_ ^ N8005;
  assign pe_i_3__68_ = pe_i_2__68_ ^ N8004;
  assign pe_i_3__67_ = pe_i_2__67_ ^ N8003;
  assign pe_i_3__66_ = pe_i_2__66_ ^ N8002;
  assign pe_i_3__65_ = pe_i_2__65_ ^ N8001;
  assign pe_i_3__64_ = pe_i_2__64_ ^ N8000;
  assign pe_i_3__63_ = pe_i_2__63_ ^ N7999;
  assign pe_i_3__62_ = pe_i_2__62_ ^ N7998;
  assign pe_i_3__61_ = pe_i_2__61_ ^ N7997;
  assign pe_i_3__60_ = pe_i_2__60_ ^ N7996;
  assign pe_i_3__59_ = pe_i_2__59_ ^ N7995;
  assign pe_i_3__58_ = pe_i_2__58_ ^ N7994;
  assign pe_i_3__57_ = pe_i_2__57_ ^ N7993;
  assign pe_i_3__56_ = pe_i_2__56_ ^ N7992;
  assign pe_i_3__55_ = pe_i_2__55_ ^ N7991;
  assign pe_i_3__54_ = pe_i_2__54_ ^ N7990;
  assign pe_i_3__53_ = pe_i_2__53_ ^ N7989;
  assign pe_i_3__52_ = pe_i_2__52_ ^ N7988;
  assign pe_i_3__51_ = pe_i_2__51_ ^ N7987;
  assign pe_i_3__50_ = pe_i_2__50_ ^ N7986;
  assign pe_i_3__49_ = pe_i_2__49_ ^ N7985;
  assign pe_i_3__48_ = pe_i_2__48_ ^ N7984;
  assign pe_i_3__47_ = pe_i_2__47_ ^ N7983;
  assign pe_i_3__46_ = pe_i_2__46_ ^ N7982;
  assign pe_i_3__45_ = pe_i_2__45_ ^ N7981;
  assign pe_i_3__44_ = pe_i_2__44_ ^ N7980;
  assign pe_i_3__43_ = pe_i_2__43_ ^ N7979;
  assign pe_i_3__42_ = pe_i_2__42_ ^ N7978;
  assign pe_i_3__41_ = pe_i_2__41_ ^ N7977;
  assign pe_i_3__40_ = pe_i_2__40_ ^ N7976;
  assign pe_i_3__39_ = pe_i_2__39_ ^ N7975;
  assign pe_i_3__38_ = pe_i_2__38_ ^ N7974;
  assign pe_i_3__37_ = pe_i_2__37_ ^ N7973;
  assign pe_i_3__36_ = pe_i_2__36_ ^ N7972;
  assign pe_i_3__35_ = pe_i_2__35_ ^ N7971;
  assign pe_i_3__34_ = pe_i_2__34_ ^ N7970;
  assign pe_i_3__33_ = pe_i_2__33_ ^ N7969;
  assign pe_i_3__32_ = pe_i_2__32_ ^ N7968;
  assign pe_i_3__31_ = pe_i_2__31_ ^ N7967;
  assign pe_i_3__30_ = pe_i_2__30_ ^ N7966;
  assign pe_i_3__29_ = pe_i_2__29_ ^ N7965;
  assign pe_i_3__28_ = pe_i_2__28_ ^ N7964;
  assign pe_i_3__27_ = pe_i_2__27_ ^ N7963;
  assign pe_i_3__26_ = pe_i_2__26_ ^ N7962;
  assign pe_i_3__25_ = pe_i_2__25_ ^ N7961;
  assign pe_i_3__24_ = pe_i_2__24_ ^ N7960;
  assign pe_i_3__23_ = pe_i_2__23_ ^ N7959;
  assign pe_i_3__22_ = pe_i_2__22_ ^ N7958;
  assign pe_i_3__21_ = pe_i_2__21_ ^ N7957;
  assign pe_i_3__20_ = pe_i_2__20_ ^ N7956;
  assign pe_i_3__19_ = pe_i_2__19_ ^ N7955;
  assign pe_i_3__18_ = pe_i_2__18_ ^ N7954;
  assign pe_i_3__17_ = pe_i_2__17_ ^ N7953;
  assign pe_i_3__16_ = pe_i_2__16_ ^ N7952;
  assign pe_i_3__15_ = pe_i_2__15_ ^ N7951;
  assign pe_i_3__14_ = pe_i_2__14_ ^ N7950;
  assign pe_i_3__13_ = pe_i_2__13_ ^ N7949;
  assign pe_i_3__12_ = pe_i_2__12_ ^ N7948;
  assign pe_i_3__11_ = pe_i_2__11_ ^ N7947;
  assign pe_i_3__10_ = pe_i_2__10_ ^ N7946;
  assign pe_i_3__9_ = pe_i_2__9_ ^ N7945;
  assign pe_i_3__8_ = pe_i_2__8_ ^ N7944;
  assign pe_i_3__7_ = pe_i_2__7_ ^ N7943;
  assign pe_i_3__6_ = pe_i_2__6_ ^ N7942;
  assign pe_i_3__5_ = pe_i_2__5_ ^ N7941;
  assign pe_i_3__4_ = pe_i_2__4_ ^ N7940;
  assign pe_i_3__3_ = pe_i_2__3_ ^ N7939;
  assign pe_i_3__2_ = pe_i_2__2_ ^ N7938;
  assign pe_i_3__1_ = pe_i_2__1_ ^ N7937;
  assign pe_i_3__0_ = pe_i_2__0_ ^ N7936;
  assign pe_i_4__126_ = pe_i_3__126_ ^ N8316;
  assign pe_i_4__125_ = pe_i_3__125_ ^ N8315;
  assign pe_i_4__124_ = pe_i_3__124_ ^ N8314;
  assign pe_i_4__123_ = pe_i_3__123_ ^ N8313;
  assign pe_i_4__122_ = pe_i_3__122_ ^ N8312;
  assign pe_i_4__121_ = pe_i_3__121_ ^ N8311;
  assign pe_i_4__120_ = pe_i_3__120_ ^ N8310;
  assign pe_i_4__119_ = pe_i_3__119_ ^ N8309;
  assign pe_i_4__118_ = pe_i_3__118_ ^ N8308;
  assign pe_i_4__117_ = pe_i_3__117_ ^ N8307;
  assign pe_i_4__116_ = pe_i_3__116_ ^ N8306;
  assign pe_i_4__115_ = pe_i_3__115_ ^ N8305;
  assign pe_i_4__114_ = pe_i_3__114_ ^ N8304;
  assign pe_i_4__113_ = pe_i_3__113_ ^ N8303;
  assign pe_i_4__112_ = pe_i_3__112_ ^ N8302;
  assign pe_i_4__111_ = pe_i_3__111_ ^ N8301;
  assign pe_i_4__110_ = pe_i_3__110_ ^ N8300;
  assign pe_i_4__109_ = pe_i_3__109_ ^ N8299;
  assign pe_i_4__108_ = pe_i_3__108_ ^ N8298;
  assign pe_i_4__107_ = pe_i_3__107_ ^ N8297;
  assign pe_i_4__106_ = pe_i_3__106_ ^ N8296;
  assign pe_i_4__105_ = pe_i_3__105_ ^ N8295;
  assign pe_i_4__104_ = pe_i_3__104_ ^ N8294;
  assign pe_i_4__103_ = pe_i_3__103_ ^ N8293;
  assign pe_i_4__102_ = pe_i_3__102_ ^ N8292;
  assign pe_i_4__101_ = pe_i_3__101_ ^ N8291;
  assign pe_i_4__100_ = pe_i_3__100_ ^ N8290;
  assign pe_i_4__99_ = pe_i_3__99_ ^ N8289;
  assign pe_i_4__98_ = pe_i_3__98_ ^ N8288;
  assign pe_i_4__97_ = pe_i_3__97_ ^ N8287;
  assign pe_i_4__96_ = pe_i_3__96_ ^ N8286;
  assign pe_i_4__95_ = pe_i_3__95_ ^ N8285;
  assign pe_i_4__94_ = pe_i_3__94_ ^ N8284;
  assign pe_i_4__93_ = pe_i_3__93_ ^ N8283;
  assign pe_i_4__92_ = pe_i_3__92_ ^ N8282;
  assign pe_i_4__91_ = pe_i_3__91_ ^ N8281;
  assign pe_i_4__90_ = pe_i_3__90_ ^ N8280;
  assign pe_i_4__89_ = pe_i_3__89_ ^ N8279;
  assign pe_i_4__88_ = pe_i_3__88_ ^ N8278;
  assign pe_i_4__87_ = pe_i_3__87_ ^ N8277;
  assign pe_i_4__86_ = pe_i_3__86_ ^ N8276;
  assign pe_i_4__85_ = pe_i_3__85_ ^ N8275;
  assign pe_i_4__84_ = pe_i_3__84_ ^ N8274;
  assign pe_i_4__83_ = pe_i_3__83_ ^ N8273;
  assign pe_i_4__82_ = pe_i_3__82_ ^ N8272;
  assign pe_i_4__81_ = pe_i_3__81_ ^ N8271;
  assign pe_i_4__80_ = pe_i_3__80_ ^ N8270;
  assign pe_i_4__79_ = pe_i_3__79_ ^ N8269;
  assign pe_i_4__78_ = pe_i_3__78_ ^ N8268;
  assign pe_i_4__77_ = pe_i_3__77_ ^ N8267;
  assign pe_i_4__76_ = pe_i_3__76_ ^ N8266;
  assign pe_i_4__75_ = pe_i_3__75_ ^ N8265;
  assign pe_i_4__74_ = pe_i_3__74_ ^ N8264;
  assign pe_i_4__73_ = pe_i_3__73_ ^ N8263;
  assign pe_i_4__72_ = pe_i_3__72_ ^ N8262;
  assign pe_i_4__71_ = pe_i_3__71_ ^ N8261;
  assign pe_i_4__70_ = pe_i_3__70_ ^ N8260;
  assign pe_i_4__69_ = pe_i_3__69_ ^ N8259;
  assign pe_i_4__68_ = pe_i_3__68_ ^ N8258;
  assign pe_i_4__67_ = pe_i_3__67_ ^ N8257;
  assign pe_i_4__66_ = pe_i_3__66_ ^ N8256;
  assign pe_i_4__65_ = pe_i_3__65_ ^ N8255;
  assign pe_i_4__64_ = pe_i_3__64_ ^ N8254;
  assign pe_i_4__63_ = pe_i_3__63_ ^ N8253;
  assign pe_i_4__62_ = pe_i_3__62_ ^ N8252;
  assign pe_i_4__61_ = pe_i_3__61_ ^ N8251;
  assign pe_i_4__60_ = pe_i_3__60_ ^ N8250;
  assign pe_i_4__59_ = pe_i_3__59_ ^ N8249;
  assign pe_i_4__58_ = pe_i_3__58_ ^ N8248;
  assign pe_i_4__57_ = pe_i_3__57_ ^ N8247;
  assign pe_i_4__56_ = pe_i_3__56_ ^ N8246;
  assign pe_i_4__55_ = pe_i_3__55_ ^ N8245;
  assign pe_i_4__54_ = pe_i_3__54_ ^ N8244;
  assign pe_i_4__53_ = pe_i_3__53_ ^ N8243;
  assign pe_i_4__52_ = pe_i_3__52_ ^ N8242;
  assign pe_i_4__51_ = pe_i_3__51_ ^ N8241;
  assign pe_i_4__50_ = pe_i_3__50_ ^ N8240;
  assign pe_i_4__49_ = pe_i_3__49_ ^ N8239;
  assign pe_i_4__48_ = pe_i_3__48_ ^ N8238;
  assign pe_i_4__47_ = pe_i_3__47_ ^ N8237;
  assign pe_i_4__46_ = pe_i_3__46_ ^ N8236;
  assign pe_i_4__45_ = pe_i_3__45_ ^ N8235;
  assign pe_i_4__44_ = pe_i_3__44_ ^ N8234;
  assign pe_i_4__43_ = pe_i_3__43_ ^ N8233;
  assign pe_i_4__42_ = pe_i_3__42_ ^ N8232;
  assign pe_i_4__41_ = pe_i_3__41_ ^ N8231;
  assign pe_i_4__40_ = pe_i_3__40_ ^ N8230;
  assign pe_i_4__39_ = pe_i_3__39_ ^ N8229;
  assign pe_i_4__38_ = pe_i_3__38_ ^ N8228;
  assign pe_i_4__37_ = pe_i_3__37_ ^ N8227;
  assign pe_i_4__36_ = pe_i_3__36_ ^ N8226;
  assign pe_i_4__35_ = pe_i_3__35_ ^ N8225;
  assign pe_i_4__34_ = pe_i_3__34_ ^ N8224;
  assign pe_i_4__33_ = pe_i_3__33_ ^ N8223;
  assign pe_i_4__32_ = pe_i_3__32_ ^ N8222;
  assign pe_i_4__31_ = pe_i_3__31_ ^ N8221;
  assign pe_i_4__30_ = pe_i_3__30_ ^ N8220;
  assign pe_i_4__29_ = pe_i_3__29_ ^ N8219;
  assign pe_i_4__28_ = pe_i_3__28_ ^ N8218;
  assign pe_i_4__27_ = pe_i_3__27_ ^ N8217;
  assign pe_i_4__26_ = pe_i_3__26_ ^ N8216;
  assign pe_i_4__25_ = pe_i_3__25_ ^ N8215;
  assign pe_i_4__24_ = pe_i_3__24_ ^ N8214;
  assign pe_i_4__23_ = pe_i_3__23_ ^ N8213;
  assign pe_i_4__22_ = pe_i_3__22_ ^ N8212;
  assign pe_i_4__21_ = pe_i_3__21_ ^ N8211;
  assign pe_i_4__20_ = pe_i_3__20_ ^ N8210;
  assign pe_i_4__19_ = pe_i_3__19_ ^ N8209;
  assign pe_i_4__18_ = pe_i_3__18_ ^ N8208;
  assign pe_i_4__17_ = pe_i_3__17_ ^ N8207;
  assign pe_i_4__16_ = pe_i_3__16_ ^ N8206;
  assign pe_i_4__15_ = pe_i_3__15_ ^ N8205;
  assign pe_i_4__14_ = pe_i_3__14_ ^ N8204;
  assign pe_i_4__13_ = pe_i_3__13_ ^ N8203;
  assign pe_i_4__12_ = pe_i_3__12_ ^ N8202;
  assign pe_i_4__11_ = pe_i_3__11_ ^ N8201;
  assign pe_i_4__10_ = pe_i_3__10_ ^ N8200;
  assign pe_i_4__9_ = pe_i_3__9_ ^ N8199;
  assign pe_i_4__8_ = pe_i_3__8_ ^ N8198;
  assign pe_i_4__7_ = pe_i_3__7_ ^ N8197;
  assign pe_i_4__6_ = pe_i_3__6_ ^ N8196;
  assign pe_i_4__5_ = pe_i_3__5_ ^ N8195;
  assign pe_i_4__4_ = pe_i_3__4_ ^ N8194;
  assign pe_i_4__3_ = pe_i_3__3_ ^ N8193;
  assign pe_i_4__2_ = pe_i_3__2_ ^ N8192;
  assign pe_i_4__1_ = pe_i_3__1_ ^ N8191;
  assign pe_i_4__0_ = pe_i_3__0_ ^ N8190;
  assign pe_i_5__126_ = pe_i_4__126_ ^ N8570;
  assign pe_i_5__125_ = pe_i_4__125_ ^ N8569;
  assign pe_i_5__124_ = pe_i_4__124_ ^ N8568;
  assign pe_i_5__123_ = pe_i_4__123_ ^ N8567;
  assign pe_i_5__122_ = pe_i_4__122_ ^ N8566;
  assign pe_i_5__121_ = pe_i_4__121_ ^ N8565;
  assign pe_i_5__120_ = pe_i_4__120_ ^ N8564;
  assign pe_i_5__119_ = pe_i_4__119_ ^ N8563;
  assign pe_i_5__118_ = pe_i_4__118_ ^ N8562;
  assign pe_i_5__117_ = pe_i_4__117_ ^ N8561;
  assign pe_i_5__116_ = pe_i_4__116_ ^ N8560;
  assign pe_i_5__115_ = pe_i_4__115_ ^ N8559;
  assign pe_i_5__114_ = pe_i_4__114_ ^ N8558;
  assign pe_i_5__113_ = pe_i_4__113_ ^ N8557;
  assign pe_i_5__112_ = pe_i_4__112_ ^ N8556;
  assign pe_i_5__111_ = pe_i_4__111_ ^ N8555;
  assign pe_i_5__110_ = pe_i_4__110_ ^ N8554;
  assign pe_i_5__109_ = pe_i_4__109_ ^ N8553;
  assign pe_i_5__108_ = pe_i_4__108_ ^ N8552;
  assign pe_i_5__107_ = pe_i_4__107_ ^ N8551;
  assign pe_i_5__106_ = pe_i_4__106_ ^ N8550;
  assign pe_i_5__105_ = pe_i_4__105_ ^ N8549;
  assign pe_i_5__104_ = pe_i_4__104_ ^ N8548;
  assign pe_i_5__103_ = pe_i_4__103_ ^ N8547;
  assign pe_i_5__102_ = pe_i_4__102_ ^ N8546;
  assign pe_i_5__101_ = pe_i_4__101_ ^ N8545;
  assign pe_i_5__100_ = pe_i_4__100_ ^ N8544;
  assign pe_i_5__99_ = pe_i_4__99_ ^ N8543;
  assign pe_i_5__98_ = pe_i_4__98_ ^ N8542;
  assign pe_i_5__97_ = pe_i_4__97_ ^ N8541;
  assign pe_i_5__96_ = pe_i_4__96_ ^ N8540;
  assign pe_i_5__95_ = pe_i_4__95_ ^ N8539;
  assign pe_i_5__94_ = pe_i_4__94_ ^ N8538;
  assign pe_i_5__93_ = pe_i_4__93_ ^ N8537;
  assign pe_i_5__92_ = pe_i_4__92_ ^ N8536;
  assign pe_i_5__91_ = pe_i_4__91_ ^ N8535;
  assign pe_i_5__90_ = pe_i_4__90_ ^ N8534;
  assign pe_i_5__89_ = pe_i_4__89_ ^ N8533;
  assign pe_i_5__88_ = pe_i_4__88_ ^ N8532;
  assign pe_i_5__87_ = pe_i_4__87_ ^ N8531;
  assign pe_i_5__86_ = pe_i_4__86_ ^ N8530;
  assign pe_i_5__85_ = pe_i_4__85_ ^ N8529;
  assign pe_i_5__84_ = pe_i_4__84_ ^ N8528;
  assign pe_i_5__83_ = pe_i_4__83_ ^ N8527;
  assign pe_i_5__82_ = pe_i_4__82_ ^ N8526;
  assign pe_i_5__81_ = pe_i_4__81_ ^ N8525;
  assign pe_i_5__80_ = pe_i_4__80_ ^ N8524;
  assign pe_i_5__79_ = pe_i_4__79_ ^ N8523;
  assign pe_i_5__78_ = pe_i_4__78_ ^ N8522;
  assign pe_i_5__77_ = pe_i_4__77_ ^ N8521;
  assign pe_i_5__76_ = pe_i_4__76_ ^ N8520;
  assign pe_i_5__75_ = pe_i_4__75_ ^ N8519;
  assign pe_i_5__74_ = pe_i_4__74_ ^ N8518;
  assign pe_i_5__73_ = pe_i_4__73_ ^ N8517;
  assign pe_i_5__72_ = pe_i_4__72_ ^ N8516;
  assign pe_i_5__71_ = pe_i_4__71_ ^ N8515;
  assign pe_i_5__70_ = pe_i_4__70_ ^ N8514;
  assign pe_i_5__69_ = pe_i_4__69_ ^ N8513;
  assign pe_i_5__68_ = pe_i_4__68_ ^ N8512;
  assign pe_i_5__67_ = pe_i_4__67_ ^ N8511;
  assign pe_i_5__66_ = pe_i_4__66_ ^ N8510;
  assign pe_i_5__65_ = pe_i_4__65_ ^ N8509;
  assign pe_i_5__64_ = pe_i_4__64_ ^ N8508;
  assign pe_i_5__63_ = pe_i_4__63_ ^ N8507;
  assign pe_i_5__62_ = pe_i_4__62_ ^ N8506;
  assign pe_i_5__61_ = pe_i_4__61_ ^ N8505;
  assign pe_i_5__60_ = pe_i_4__60_ ^ N8504;
  assign pe_i_5__59_ = pe_i_4__59_ ^ N8503;
  assign pe_i_5__58_ = pe_i_4__58_ ^ N8502;
  assign pe_i_5__57_ = pe_i_4__57_ ^ N8501;
  assign pe_i_5__56_ = pe_i_4__56_ ^ N8500;
  assign pe_i_5__55_ = pe_i_4__55_ ^ N8499;
  assign pe_i_5__54_ = pe_i_4__54_ ^ N8498;
  assign pe_i_5__53_ = pe_i_4__53_ ^ N8497;
  assign pe_i_5__52_ = pe_i_4__52_ ^ N8496;
  assign pe_i_5__51_ = pe_i_4__51_ ^ N8495;
  assign pe_i_5__50_ = pe_i_4__50_ ^ N8494;
  assign pe_i_5__49_ = pe_i_4__49_ ^ N8493;
  assign pe_i_5__48_ = pe_i_4__48_ ^ N8492;
  assign pe_i_5__47_ = pe_i_4__47_ ^ N8491;
  assign pe_i_5__46_ = pe_i_4__46_ ^ N8490;
  assign pe_i_5__45_ = pe_i_4__45_ ^ N8489;
  assign pe_i_5__44_ = pe_i_4__44_ ^ N8488;
  assign pe_i_5__43_ = pe_i_4__43_ ^ N8487;
  assign pe_i_5__42_ = pe_i_4__42_ ^ N8486;
  assign pe_i_5__41_ = pe_i_4__41_ ^ N8485;
  assign pe_i_5__40_ = pe_i_4__40_ ^ N8484;
  assign pe_i_5__39_ = pe_i_4__39_ ^ N8483;
  assign pe_i_5__38_ = pe_i_4__38_ ^ N8482;
  assign pe_i_5__37_ = pe_i_4__37_ ^ N8481;
  assign pe_i_5__36_ = pe_i_4__36_ ^ N8480;
  assign pe_i_5__35_ = pe_i_4__35_ ^ N8479;
  assign pe_i_5__34_ = pe_i_4__34_ ^ N8478;
  assign pe_i_5__33_ = pe_i_4__33_ ^ N8477;
  assign pe_i_5__32_ = pe_i_4__32_ ^ N8476;
  assign pe_i_5__31_ = pe_i_4__31_ ^ N8475;
  assign pe_i_5__30_ = pe_i_4__30_ ^ N8474;
  assign pe_i_5__29_ = pe_i_4__29_ ^ N8473;
  assign pe_i_5__28_ = pe_i_4__28_ ^ N8472;
  assign pe_i_5__27_ = pe_i_4__27_ ^ N8471;
  assign pe_i_5__26_ = pe_i_4__26_ ^ N8470;
  assign pe_i_5__25_ = pe_i_4__25_ ^ N8469;
  assign pe_i_5__24_ = pe_i_4__24_ ^ N8468;
  assign pe_i_5__23_ = pe_i_4__23_ ^ N8467;
  assign pe_i_5__22_ = pe_i_4__22_ ^ N8466;
  assign pe_i_5__21_ = pe_i_4__21_ ^ N8465;
  assign pe_i_5__20_ = pe_i_4__20_ ^ N8464;
  assign pe_i_5__19_ = pe_i_4__19_ ^ N8463;
  assign pe_i_5__18_ = pe_i_4__18_ ^ N8462;
  assign pe_i_5__17_ = pe_i_4__17_ ^ N8461;
  assign pe_i_5__16_ = pe_i_4__16_ ^ N8460;
  assign pe_i_5__15_ = pe_i_4__15_ ^ N8459;
  assign pe_i_5__14_ = pe_i_4__14_ ^ N8458;
  assign pe_i_5__13_ = pe_i_4__13_ ^ N8457;
  assign pe_i_5__12_ = pe_i_4__12_ ^ N8456;
  assign pe_i_5__11_ = pe_i_4__11_ ^ N8455;
  assign pe_i_5__10_ = pe_i_4__10_ ^ N8454;
  assign pe_i_5__9_ = pe_i_4__9_ ^ N8453;
  assign pe_i_5__8_ = pe_i_4__8_ ^ N8452;
  assign pe_i_5__7_ = pe_i_4__7_ ^ N8451;
  assign pe_i_5__6_ = pe_i_4__6_ ^ N8450;
  assign pe_i_5__5_ = pe_i_4__5_ ^ N8449;
  assign pe_i_5__4_ = pe_i_4__4_ ^ N8448;
  assign pe_i_5__3_ = pe_i_4__3_ ^ N8447;
  assign pe_i_5__2_ = pe_i_4__2_ ^ N8446;
  assign pe_i_5__1_ = pe_i_4__1_ ^ N8445;
  assign pe_i_5__0_ = pe_i_4__0_ ^ N8444;
  assign pe_i_6__126_ = pe_i_5__126_ ^ N8824;
  assign pe_i_6__125_ = pe_i_5__125_ ^ N8823;
  assign pe_i_6__124_ = pe_i_5__124_ ^ N8822;
  assign pe_i_6__123_ = pe_i_5__123_ ^ N8821;
  assign pe_i_6__122_ = pe_i_5__122_ ^ N8820;
  assign pe_i_6__121_ = pe_i_5__121_ ^ N8819;
  assign pe_i_6__120_ = pe_i_5__120_ ^ N8818;
  assign pe_i_6__119_ = pe_i_5__119_ ^ N8817;
  assign pe_i_6__118_ = pe_i_5__118_ ^ N8816;
  assign pe_i_6__117_ = pe_i_5__117_ ^ N8815;
  assign pe_i_6__116_ = pe_i_5__116_ ^ N8814;
  assign pe_i_6__115_ = pe_i_5__115_ ^ N8813;
  assign pe_i_6__114_ = pe_i_5__114_ ^ N8812;
  assign pe_i_6__113_ = pe_i_5__113_ ^ N8811;
  assign pe_i_6__112_ = pe_i_5__112_ ^ N8810;
  assign pe_i_6__111_ = pe_i_5__111_ ^ N8809;
  assign pe_i_6__110_ = pe_i_5__110_ ^ N8808;
  assign pe_i_6__109_ = pe_i_5__109_ ^ N8807;
  assign pe_i_6__108_ = pe_i_5__108_ ^ N8806;
  assign pe_i_6__107_ = pe_i_5__107_ ^ N8805;
  assign pe_i_6__106_ = pe_i_5__106_ ^ N8804;
  assign pe_i_6__105_ = pe_i_5__105_ ^ N8803;
  assign pe_i_6__104_ = pe_i_5__104_ ^ N8802;
  assign pe_i_6__103_ = pe_i_5__103_ ^ N8801;
  assign pe_i_6__102_ = pe_i_5__102_ ^ N8800;
  assign pe_i_6__101_ = pe_i_5__101_ ^ N8799;
  assign pe_i_6__100_ = pe_i_5__100_ ^ N8798;
  assign pe_i_6__99_ = pe_i_5__99_ ^ N8797;
  assign pe_i_6__98_ = pe_i_5__98_ ^ N8796;
  assign pe_i_6__97_ = pe_i_5__97_ ^ N8795;
  assign pe_i_6__96_ = pe_i_5__96_ ^ N8794;
  assign pe_i_6__95_ = pe_i_5__95_ ^ N8793;
  assign pe_i_6__94_ = pe_i_5__94_ ^ N8792;
  assign pe_i_6__93_ = pe_i_5__93_ ^ N8791;
  assign pe_i_6__92_ = pe_i_5__92_ ^ N8790;
  assign pe_i_6__91_ = pe_i_5__91_ ^ N8789;
  assign pe_i_6__90_ = pe_i_5__90_ ^ N8788;
  assign pe_i_6__89_ = pe_i_5__89_ ^ N8787;
  assign pe_i_6__88_ = pe_i_5__88_ ^ N8786;
  assign pe_i_6__87_ = pe_i_5__87_ ^ N8785;
  assign pe_i_6__86_ = pe_i_5__86_ ^ N8784;
  assign pe_i_6__85_ = pe_i_5__85_ ^ N8783;
  assign pe_i_6__84_ = pe_i_5__84_ ^ N8782;
  assign pe_i_6__83_ = pe_i_5__83_ ^ N8781;
  assign pe_i_6__82_ = pe_i_5__82_ ^ N8780;
  assign pe_i_6__81_ = pe_i_5__81_ ^ N8779;
  assign pe_i_6__80_ = pe_i_5__80_ ^ N8778;
  assign pe_i_6__79_ = pe_i_5__79_ ^ N8777;
  assign pe_i_6__78_ = pe_i_5__78_ ^ N8776;
  assign pe_i_6__77_ = pe_i_5__77_ ^ N8775;
  assign pe_i_6__76_ = pe_i_5__76_ ^ N8774;
  assign pe_i_6__75_ = pe_i_5__75_ ^ N8773;
  assign pe_i_6__74_ = pe_i_5__74_ ^ N8772;
  assign pe_i_6__73_ = pe_i_5__73_ ^ N8771;
  assign pe_i_6__72_ = pe_i_5__72_ ^ N8770;
  assign pe_i_6__71_ = pe_i_5__71_ ^ N8769;
  assign pe_i_6__70_ = pe_i_5__70_ ^ N8768;
  assign pe_i_6__69_ = pe_i_5__69_ ^ N8767;
  assign pe_i_6__68_ = pe_i_5__68_ ^ N8766;
  assign pe_i_6__67_ = pe_i_5__67_ ^ N8765;
  assign pe_i_6__66_ = pe_i_5__66_ ^ N8764;
  assign pe_i_6__65_ = pe_i_5__65_ ^ N8763;
  assign pe_i_6__64_ = pe_i_5__64_ ^ N8762;
  assign pe_i_6__63_ = pe_i_5__63_ ^ N8761;
  assign pe_i_6__62_ = pe_i_5__62_ ^ N8760;
  assign pe_i_6__61_ = pe_i_5__61_ ^ N8759;
  assign pe_i_6__60_ = pe_i_5__60_ ^ N8758;
  assign pe_i_6__59_ = pe_i_5__59_ ^ N8757;
  assign pe_i_6__58_ = pe_i_5__58_ ^ N8756;
  assign pe_i_6__57_ = pe_i_5__57_ ^ N8755;
  assign pe_i_6__56_ = pe_i_5__56_ ^ N8754;
  assign pe_i_6__55_ = pe_i_5__55_ ^ N8753;
  assign pe_i_6__54_ = pe_i_5__54_ ^ N8752;
  assign pe_i_6__53_ = pe_i_5__53_ ^ N8751;
  assign pe_i_6__52_ = pe_i_5__52_ ^ N8750;
  assign pe_i_6__51_ = pe_i_5__51_ ^ N8749;
  assign pe_i_6__50_ = pe_i_5__50_ ^ N8748;
  assign pe_i_6__49_ = pe_i_5__49_ ^ N8747;
  assign pe_i_6__48_ = pe_i_5__48_ ^ N8746;
  assign pe_i_6__47_ = pe_i_5__47_ ^ N8745;
  assign pe_i_6__46_ = pe_i_5__46_ ^ N8744;
  assign pe_i_6__45_ = pe_i_5__45_ ^ N8743;
  assign pe_i_6__44_ = pe_i_5__44_ ^ N8742;
  assign pe_i_6__43_ = pe_i_5__43_ ^ N8741;
  assign pe_i_6__42_ = pe_i_5__42_ ^ N8740;
  assign pe_i_6__41_ = pe_i_5__41_ ^ N8739;
  assign pe_i_6__40_ = pe_i_5__40_ ^ N8738;
  assign pe_i_6__39_ = pe_i_5__39_ ^ N8737;
  assign pe_i_6__38_ = pe_i_5__38_ ^ N8736;
  assign pe_i_6__37_ = pe_i_5__37_ ^ N8735;
  assign pe_i_6__36_ = pe_i_5__36_ ^ N8734;
  assign pe_i_6__35_ = pe_i_5__35_ ^ N8733;
  assign pe_i_6__34_ = pe_i_5__34_ ^ N8732;
  assign pe_i_6__33_ = pe_i_5__33_ ^ N8731;
  assign pe_i_6__32_ = pe_i_5__32_ ^ N8730;
  assign pe_i_6__31_ = pe_i_5__31_ ^ N8729;
  assign pe_i_6__30_ = pe_i_5__30_ ^ N8728;
  assign pe_i_6__29_ = pe_i_5__29_ ^ N8727;
  assign pe_i_6__28_ = pe_i_5__28_ ^ N8726;
  assign pe_i_6__27_ = pe_i_5__27_ ^ N8725;
  assign pe_i_6__26_ = pe_i_5__26_ ^ N8724;
  assign pe_i_6__25_ = pe_i_5__25_ ^ N8723;
  assign pe_i_6__24_ = pe_i_5__24_ ^ N8722;
  assign pe_i_6__23_ = pe_i_5__23_ ^ N8721;
  assign pe_i_6__22_ = pe_i_5__22_ ^ N8720;
  assign pe_i_6__21_ = pe_i_5__21_ ^ N8719;
  assign pe_i_6__20_ = pe_i_5__20_ ^ N8718;
  assign pe_i_6__19_ = pe_i_5__19_ ^ N8717;
  assign pe_i_6__18_ = pe_i_5__18_ ^ N8716;
  assign pe_i_6__17_ = pe_i_5__17_ ^ N8715;
  assign pe_i_6__16_ = pe_i_5__16_ ^ N8714;
  assign pe_i_6__15_ = pe_i_5__15_ ^ N8713;
  assign pe_i_6__14_ = pe_i_5__14_ ^ N8712;
  assign pe_i_6__13_ = pe_i_5__13_ ^ N8711;
  assign pe_i_6__12_ = pe_i_5__12_ ^ N8710;
  assign pe_i_6__11_ = pe_i_5__11_ ^ N8709;
  assign pe_i_6__10_ = pe_i_5__10_ ^ N8708;
  assign pe_i_6__9_ = pe_i_5__9_ ^ N8707;
  assign pe_i_6__8_ = pe_i_5__8_ ^ N8706;
  assign pe_i_6__7_ = pe_i_5__7_ ^ N8705;
  assign pe_i_6__6_ = pe_i_5__6_ ^ N8704;
  assign pe_i_6__5_ = pe_i_5__5_ ^ N8703;
  assign pe_i_6__4_ = pe_i_5__4_ ^ N8702;
  assign pe_i_6__3_ = pe_i_5__3_ ^ N8701;
  assign pe_i_6__2_ = pe_i_5__2_ ^ N8700;
  assign pe_i_6__1_ = pe_i_5__1_ ^ N8699;
  assign pe_i_6__0_ = pe_i_5__0_ ^ N8698;

endmodule

